-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 12 2019 13:57:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : inout std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__37526\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal \c0.tx.n4414\ : std_logic;
signal \c0.tx.n4415\ : std_logic;
signal \c0.tx.n4416\ : std_logic;
signal \c0.tx.n4417\ : std_logic;
signal \c0.tx.n4418\ : std_logic;
signal \c0.tx.n4419\ : std_logic;
signal \c0.tx.n4420\ : std_logic;
signal \c0.tx.n4421\ : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal \n5037_cascade_\ : std_logic;
signal n3611 : std_logic;
signal \n4_adj_2008_cascade_\ : std_logic;
signal \c0.tx2.n5312_cascade_\ : std_logic;
signal \c0.n5815_cascade_\ : std_logic;
signal \c0.n5818\ : std_logic;
signal \c0.tx2.n5932_cascade_\ : std_logic;
signal \c0.n5917_cascade_\ : std_logic;
signal \c0.n5920_cascade_\ : std_logic;
signal \c0.n5662\ : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal \c0.tx2.n5929\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal \c0.n5399_cascade_\ : std_logic;
signal \c0.n5857_cascade_\ : std_logic;
signal \c0.n5860\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_1798\ : std_logic;
signal \n3_cascade_\ : std_logic;
signal \c0.data_in_frame_19_0\ : std_logic;
signal tx2_o : std_logic;
signal tx2_enable : std_logic;
signal \c0.n5402\ : std_logic;
signal \c0.data_in_frame_19_3\ : std_logic;
signal \c0.n5863\ : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal \c0.rx.n4422\ : std_logic;
signal \c0.rx.n4423\ : std_logic;
signal \c0.rx.n4424\ : std_logic;
signal \c0.rx.n4425\ : std_logic;
signal \c0.rx.n4426\ : std_logic;
signal \c0.rx.n4427\ : std_logic;
signal \c0.rx.n4428\ : std_logic;
signal \n2156_cascade_\ : std_logic;
signal n8 : std_logic;
signal \c0.rx.n5298_cascade_\ : std_logic;
signal \c0.rx.n5536\ : std_logic;
signal \c0.rx.n5049\ : std_logic;
signal n5050 : std_logic;
signal \c0.rx.n5923_cascade_\ : std_logic;
signal \c0.rx.n5926_cascade_\ : std_logic;
signal \c0.rx.n5537\ : std_logic;
signal n5490 : std_logic;
signal \c0.rx.n3980_cascade_\ : std_logic;
signal \c0.rx.n5532\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \c0.n4378\ : std_logic;
signal \c0.tx_transmit_N_568_2\ : std_logic;
signal \c0.n4379\ : std_logic;
signal \c0.tx_transmit_N_568_3\ : std_logic;
signal \c0.n4380\ : std_logic;
signal \c0.n4381\ : std_logic;
signal \c0.byte_transmit_counter_5\ : std_logic;
signal \c0.n4382\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.n4383\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.n4384\ : std_logic;
signal \c0.n50\ : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \c0.n5540_cascade_\ : std_logic;
signal \c0.n5977_cascade_\ : std_logic;
signal \n1760_cascade_\ : std_logic;
signal n1760 : std_logic;
signal \c0.n1529_cascade_\ : std_logic;
signal \c0.n1801\ : std_logic;
signal \c0.tx.n315\ : std_logic;
signal n319 : std_logic;
signal \c0.tx.n320\ : std_logic;
signal \c0.tx.n321\ : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal \c0.tx.n313\ : std_logic;
signal n316 : std_logic;
signal n314 : std_logic;
signal n317 : std_logic;
signal \r_Clock_Count_2\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \r_Clock_Count_5\ : std_logic;
signal \r_Clock_Count_4\ : std_logic;
signal \c0.tx.n5_cascade_\ : std_logic;
signal \r_Clock_Count_7\ : std_logic;
signal \n3595_cascade_\ : std_logic;
signal \c0.tx.n5520\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx2.n5_cascade_\ : std_logic;
signal \c0.tx2.n3591\ : std_logic;
signal \c0.tx2.n3591_cascade_\ : std_logic;
signal \r_SM_Main_2_N_1767_1_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_0\ : std_logic;
signal n2460 : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal \c0.tx2.r_Clock_Count_1\ : std_logic;
signal n2399 : std_logic;
signal \c0.tx2.n4429\ : std_logic;
signal \c0.tx2.n4430\ : std_logic;
signal \c0.tx2.n4431\ : std_logic;
signal \c0.tx2.r_Clock_Count_4\ : std_logic;
signal n2382 : std_logic;
signal \c0.tx2.n4432\ : std_logic;
signal \c0.tx2.r_Clock_Count_5\ : std_logic;
signal n2379 : std_logic;
signal \c0.tx2.n4433\ : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal n2376 : std_logic;
signal \c0.tx2.n4434\ : std_logic;
signal \c0.tx2.n4435\ : std_logic;
signal \c0.tx2.n4436\ : std_logic;
signal \r_Clock_Count_8_adj_2012\ : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal n2369 : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal \c0.tx2.n5947\ : std_logic;
signal \c0.tx2.n5950\ : std_logic;
signal n1345 : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal \c0.n5665_cascade_\ : std_logic;
signal \c0.n5372_cascade_\ : std_logic;
signal \c0.n5659\ : std_logic;
signal \c0.n5938\ : std_logic;
signal \c0.n5971_cascade_\ : std_logic;
signal \c0.n5725_cascade_\ : std_logic;
signal \c0.n1058\ : std_logic;
signal \c0.n5728_cascade_\ : std_logic;
signal \c0.n5974\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.tx2.n1592\ : std_logic;
signal \c0.n5803_cascade_\ : std_logic;
signal \c0.data_in_frame_18_1\ : std_logic;
signal \c0.n5369\ : std_logic;
signal \c0.n5869\ : std_logic;
signal \c0.n5959\ : std_logic;
signal \c0.n5962\ : std_logic;
signal \c0.data_in_frame_18_3\ : std_logic;
signal n5051 : std_logic;
signal n5491 : std_logic;
signal \c0.rx.n5535\ : std_logic;
signal \c0.rx.n2157\ : std_logic;
signal \c0.rx.n5538\ : std_logic;
signal \c0.rx.n5539\ : std_logic;
signal \c0.rx.n40\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_1824_2_cascade_\ : std_logic;
signal n4474 : std_logic;
signal n2156 : std_logic;
signal \n4474_cascade_\ : std_logic;
signal \c0.rx.n4_adj_1866_cascade_\ : std_logic;
signal \c0.rx.n4011\ : std_logic;
signal data_in_5_1 : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal \c0.rx.n37\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.n37_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \r_SM_Main_2_N_1830_0\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \n12_adj_1995_cascade_\ : std_logic;
signal n5316 : std_logic;
signal n16_adj_1993 : std_logic;
signal \c0.rx.n3573\ : std_logic;
signal \c0.rx.n3573_cascade_\ : std_logic;
signal \c0.n20_adj_1918_cascade_\ : std_logic;
signal \c0.n87\ : std_logic;
signal \c0.n87_cascade_\ : std_logic;
signal \c0.n16_adj_1909\ : std_logic;
signal \c0.tx_transmit_N_568_5\ : std_logic;
signal \c0.tx_transmit_N_568_6\ : std_logic;
signal \c0.tx_transmit_N_568_7\ : std_logic;
signal \c0.tx_transmit_N_568_4\ : std_logic;
signal \c0.n103\ : std_logic;
signal \c0.n109\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.n109_cascade_\ : std_logic;
signal \n4315_cascade_\ : std_logic;
signal \n4316_cascade_\ : std_logic;
signal n7_adj_2002 : std_logic;
signal n5066 : std_logic;
signal tx_active : std_logic;
signal data_out_19_4 : std_logic;
signal data_out_18_4 : std_logic;
signal \c0.n17_cascade_\ : std_logic;
signal \tx_data_4_N_keep_cascade_\ : std_logic;
signal n8_adj_2001 : std_logic;
signal \c0.tx.r_SM_Main_2_N_1767_1_cascade_\ : std_logic;
signal n5041 : std_logic;
signal \c0.tx_transmit\ : std_logic;
signal \c0.tx.n12_cascade_\ : std_logic;
signal \r_Clock_Count_8\ : std_logic;
signal \n1307_cascade_\ : std_logic;
signal n3595 : std_logic;
signal n4221 : std_logic;
signal n2 : std_logic;
signal n1307 : std_logic;
signal \n4_adj_2003_cascade_\ : std_logic;
signal n4155 : std_logic;
signal n2372 : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal n2395 : std_logic;
signal \c0.tx2.r_Clock_Count_2\ : std_logic;
signal \r_SM_Main_0_adj_2011\ : std_logic;
signal \r_SM_Main_2_N_1767_1\ : std_logic;
signal \r_SM_Main_1_adj_2010\ : std_logic;
signal \c0.tx2.n2218_cascade_\ : std_logic;
signal \c0.tx2.n3577\ : std_logic;
signal \c0.n5953\ : std_logic;
signal \c0.n5956\ : std_logic;
signal n2392 : std_logic;
signal \r_SM_Main_2_adj_2009\ : std_logic;
signal n5037 : std_logic;
signal \c0.tx2.r_Clock_Count_3\ : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal \c0.n4400\ : std_logic;
signal \c0.n4401\ : std_logic;
signal \c0.n4402\ : std_logic;
signal \c0.n4403\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.n5785_cascade_\ : std_logic;
signal \c0.n5426\ : std_logic;
signal \c0.n5788\ : std_logic;
signal \c0.n5968\ : std_logic;
signal \c0.n5363\ : std_logic;
signal \c0.data_in_frame_19_7\ : std_logic;
signal \c0.n5935\ : std_logic;
signal \c0.n5944\ : std_logic;
signal \c0.data_in_frame_19_6\ : std_logic;
signal \c0.n5456\ : std_logic;
signal data_in_18_3 : std_logic;
signal \c0.n1893_cascade_\ : std_logic;
signal \c0.n20_adj_1921\ : std_logic;
signal \c0.n5459\ : std_logic;
signal \c0.n5737\ : std_logic;
signal \c0.data_in_frame_19_1\ : std_logic;
signal \c0.data_in_field_131\ : std_logic;
signal \c0.n2036_cascade_\ : std_logic;
signal \c0.n5273_cascade_\ : std_logic;
signal \c0.data_in_frame_18_7\ : std_logic;
signal \c0.n5671\ : std_logic;
signal rx_data_3 : std_logic;
signal rx_data_5 : std_logic;
signal \r_Clock_Count_7_adj_2004\ : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal \c0.rx.n6\ : std_logic;
signal \c0.rx.n2213\ : std_logic;
signal \c0.rx.n2317\ : std_logic;
signal \c0.rx.r_Bit_Index_1\ : std_logic;
signal \c0.rx.r_Bit_Index_2\ : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal \r_Clock_Count_6\ : std_logic;
signal n8_adj_1996 : std_logic;
signal tx_enable : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.n4404\ : std_logic;
signal \c0.n4405\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.n4406\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.n4407\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.n4408\ : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.n4409\ : std_logic;
signal \c0.n4410\ : std_logic;
signal \c0.n4411\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal \c0.n4412\ : std_logic;
signal \c0.n4413\ : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal n5077 : std_logic;
signal n4_adj_1988 : std_logic;
signal data_out_19_0 : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.n18_adj_1908\ : std_logic;
signal n4_adj_2000 : std_logic;
signal \n5086_cascade_\ : std_logic;
signal n1525 : std_logic;
signal \n5156_cascade_\ : std_logic;
signal data_out_18_0 : std_logic;
signal n5156 : std_logic;
signal n5063 : std_logic;
signal data_out_18_3 : std_logic;
signal data_out_19_7 : std_logic;
signal n7_adj_1998 : std_logic;
signal n8_adj_1997 : std_logic;
signal data_out_18_7 : std_logic;
signal data_out_19_3 : std_logic;
signal data_out_18_1 : std_logic;
signal n4_adj_2007 : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \c0.n9\ : std_logic;
signal \c0.n5501\ : std_logic;
signal \c0.n1173_cascade_\ : std_logic;
signal \tx_data_0_N_keep_cascade_\ : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \c0.n5531\ : std_logic;
signal \c0.n15_cascade_\ : std_logic;
signal \tx_data_1_N_keep\ : std_logic;
signal \c0.tx.r_SM_Main_2_N_1767_1\ : std_logic;
signal \c0.tx.n3507\ : std_logic;
signal \c0.tx.n3507_cascade_\ : std_logic;
signal n2307 : std_logic;
signal n2200 : std_logic;
signal \n2307_cascade_\ : std_logic;
signal n805 : std_logic;
signal \c0.tx2.r_Bit_Index_0\ : std_logic;
signal \c0.tx2.r_Bit_Index_1\ : std_logic;
signal \c0.tx2.r_Bit_Index_2\ : std_logic;
signal \c0.tx2.n2218\ : std_logic;
signal \c0.tx2.n2319\ : std_logic;
signal n5153 : std_logic;
signal \c0.n3414_cascade_\ : std_logic;
signal \c0.n3414\ : std_logic;
signal \c0.FRAME_MATCHER_wait_for_transmission_N_909\ : std_logic;
signal \c0.r_SM_Main_2_N_1770_0\ : std_logic;
signal tx2_active : std_logic;
signal \c0.n195\ : std_logic;
signal \c0.n5845_cascade_\ : std_logic;
signal \c0.n2275\ : std_logic;
signal \c0.data_in_field_81\ : std_logic;
signal \c0.n1918_cascade_\ : std_logic;
signal \c0.n5192_cascade_\ : std_logic;
signal \c0.n30_adj_1897_cascade_\ : std_logic;
signal \c0.n36_cascade_\ : std_logic;
signal \c0.n5080_cascade_\ : std_logic;
signal \c0.n1990\ : std_logic;
signal \c0.n5192\ : std_logic;
signal \c0.n5080\ : std_logic;
signal \c0.n23_adj_1931\ : std_logic;
signal \c0.n21_adj_1928\ : std_logic;
signal \c0.n22_adj_1927_cascade_\ : std_logic;
signal \c0.n24_adj_1907\ : std_logic;
signal data_in_19_3 : std_logic;
signal \c0.data_in_frame_18_0\ : std_logic;
signal \c0.data_in_frame_18_4\ : std_logic;
signal \c0.n22_adj_1881\ : std_logic;
signal \c0.n5266\ : std_logic;
signal \c0.data_in_field_101\ : std_logic;
signal \c0.n18_adj_1882_cascade_\ : std_logic;
signal \c0.n26_adj_1883\ : std_logic;
signal \c0.n5462\ : std_logic;
signal data_in_12_5 : std_logic;
signal \c0.n5222_cascade_\ : std_logic;
signal \c0.n42\ : std_logic;
signal \c0.n33_cascade_\ : std_logic;
signal \c0.n2008_cascade_\ : std_logic;
signal \c0.n38_cascade_\ : std_logic;
signal \c0.data_in_frame_18_6\ : std_logic;
signal data_in_2_5 : std_logic;
signal rx_data_6 : std_logic;
signal \c0.rx.n2151_cascade_\ : std_logic;
signal \n1709_cascade_\ : std_logic;
signal n4_adj_1990 : std_logic;
signal rx_data_4 : std_logic;
signal n4_adj_1992 : std_logic;
signal data_out_11_0 : std_logic;
signal data_out_18_2 : std_logic;
signal data_out_19_2 : std_logic;
signal \c0.n2249\ : std_logic;
signal \c0.n5522_cascade_\ : std_logic;
signal n4_adj_1991 : std_logic;
signal data_out_18_5 : std_logic;
signal n4_adj_1994 : std_logic;
signal n5135 : std_logic;
signal n5117 : std_logic;
signal \n5117_cascade_\ : std_logic;
signal n4316 : std_logic;
signal data_out_19_5 : std_logic;
signal \tx_data_2_N_keep\ : std_logic;
signal data_out_11_3 : std_logic;
signal data_out_11_2 : std_logic;
signal \c0.n1805_cascade_\ : std_logic;
signal n135 : std_logic;
signal \c0.n1805\ : std_logic;
signal n5173 : std_logic;
signal data_out_11_7 : std_logic;
signal data_out_10_7 : std_logic;
signal n5079 : std_logic;
signal data_out_19_1 : std_logic;
signal \c0.n5519\ : std_logic;
signal \c0.n5980\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.tx.n5713_cascade_\ : std_logic;
signal data_out_11_1 : std_logic;
signal \c0.n9_adj_1880\ : std_logic;
signal \c0.n9_adj_1890\ : std_logic;
signal \c0.n5489\ : std_logic;
signal \c0.n991_cascade_\ : std_logic;
signal \tx_data_5_N_keep_cascade_\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \tx_data_3_N_keep\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \c0.tx.n5719\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \c0.tx.n5716\ : std_logic;
signal \c0.tx.n5722\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \c0.tx.o_Tx_Serial_N_1798_cascade_\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \c0.tx.n3_cascade_\ : std_logic;
signal tx_o : std_logic;
signal \c0.n2018\ : std_logic;
signal \c0.data_in_frame_18_2\ : std_logic;
signal \c0.n5965\ : std_logic;
signal data_in_19_6 : std_logic;
signal \c0.n22_adj_1901_cascade_\ : std_logic;
signal \c0.n23_adj_1932\ : std_logic;
signal \c0.n30_adj_1940_cascade_\ : std_logic;
signal \c0.n3563\ : std_logic;
signal \c0.n5280\ : std_logic;
signal \c0.n5277\ : std_logic;
signal \c0.n25_adj_1941\ : std_logic;
signal \c0.n5072\ : std_logic;
signal \c0.n26_adj_1915_cascade_\ : std_logic;
signal data_in_17_3 : std_logic;
signal \c0.data_in_field_71\ : std_logic;
signal \c0.n26_cascade_\ : std_logic;
signal \c0.n27_adj_1919\ : std_logic;
signal \c0.n5250\ : std_logic;
signal \c0.n28_adj_1917_cascade_\ : std_logic;
signal \c0.n26_adj_1939\ : std_logic;
signal \c0.data_in_field_41\ : std_logic;
signal \c0.n14_cascade_\ : std_logic;
signal \c0.n15_adj_1894\ : std_logic;
signal \c0.n16_adj_1893_cascade_\ : std_logic;
signal \c0.n22_adj_1930\ : std_logic;
signal \c0.n2058\ : std_logic;
signal \c0.n5096_cascade_\ : std_logic;
signal \c0.n1785_cascade_\ : std_logic;
signal \c0.n22\ : std_logic;
signal data_in_13_5 : std_logic;
signal \c0.n5150\ : std_logic;
signal \c0.data_in_field_109\ : std_logic;
signal \c0.n39\ : std_logic;
signal \c0.n45_adj_1885\ : std_logic;
signal \c0.n43\ : std_logic;
signal \c0.n30\ : std_logic;
signal \c0.n5275_cascade_\ : std_logic;
signal \c0.n24_adj_1929\ : std_logic;
signal \c0.n5182\ : std_logic;
signal \c0.n5147\ : std_logic;
signal \c0.n5182_cascade_\ : std_logic;
signal \c0.n40\ : std_logic;
signal \c0.data_in_field_119\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n20_adj_1906\ : std_logic;
signal data_in_4_3 : std_logic;
signal data_in_16_6 : std_logic;
signal \c0.n5731\ : std_logic;
signal \c0.n5264\ : std_logic;
signal \c0.n5264_cascade_\ : std_logic;
signal data_in_19_1 : std_logic;
signal data_in_2_3 : std_logic;
signal \r_SM_Main_2_adj_2005\ : std_logic;
signal \c0.rx.r_SM_Main_1\ : std_logic;
signal \c0.rx.n5058\ : std_logic;
signal \c0.rx.r_Bit_Index_0\ : std_logic;
signal \r_SM_Main_0_adj_2006\ : std_logic;
signal \c0.rx.n5058_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_1824_2\ : std_logic;
signal n4 : std_logic;
signal \n1714_cascade_\ : std_logic;
signal rx_data_1 : std_logic;
signal data_in_0_7 : std_logic;
signal n4_adj_1986 : std_logic;
signal n1709 : std_logic;
signal data_0 : std_logic;
signal \bfn_6_17_0_\ : std_logic;
signal data_1 : std_logic;
signal \c0.n4385\ : std_logic;
signal data_2 : std_logic;
signal \c0.n4386\ : std_logic;
signal data_3 : std_logic;
signal \c0.n4387\ : std_logic;
signal \c0.n4388\ : std_logic;
signal data_5 : std_logic;
signal \c0.n4389\ : std_logic;
signal data_6 : std_logic;
signal \c0.n4390\ : std_logic;
signal data_7 : std_logic;
signal \c0.n4391\ : std_logic;
signal \c0.n4392\ : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal data_9 : std_logic;
signal \c0.n4393\ : std_logic;
signal \c0.n4394\ : std_logic;
signal data_11 : std_logic;
signal \c0.n4395\ : std_logic;
signal data_12 : std_logic;
signal \c0.n4396\ : std_logic;
signal data_13 : std_logic;
signal \c0.n4397\ : std_logic;
signal \c0.n4398\ : std_logic;
signal \c0.n4399\ : std_logic;
signal data_15 : std_logic;
signal data_4 : std_logic;
signal data_14 : std_logic;
signal data_out_11_4 : std_logic;
signal data_out_10_4 : std_logic;
signal \c0.n9_adj_1887_cascade_\ : std_logic;
signal \c0.n15_adj_1889\ : std_logic;
signal data_8 : std_logic;
signal \c0.n17_adj_1961\ : std_logic;
signal \c0.n1236_cascade_\ : std_logic;
signal \c0.n2247\ : std_logic;
signal \c0.n1227\ : std_logic;
signal \c0.n5511_cascade_\ : std_logic;
signal \tx_data_7_N_keep_cascade_\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal n1442 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal data_out_10_0 : std_logic;
signal n1748 : std_logic;
signal n21_adj_1999 : std_logic;
signal data_10 : std_logic;
signal n4315 : std_logic;
signal data_out_10_2 : std_logic;
signal \c0.n5411\ : std_logic;
signal \c0.n5830\ : std_logic;
signal \c0.n5941\ : std_logic;
signal \c0.data_in_frame_19_2\ : std_logic;
signal \c0.data_in_frame_18_5\ : std_logic;
signal \c0.data_in_frame_19_5\ : std_logic;
signal data_in_14_5 : std_logic;
signal \c0.n5809\ : std_logic;
signal \c0.n5241\ : std_logic;
signal \c0.tx2_transmit_N_1031_cascade_\ : std_logic;
signal \c0.n38_adj_1934\ : std_logic;
signal \c0.n14_adj_1900\ : std_logic;
signal data_in_15_0 : std_logic;
signal \c0.n5210\ : std_logic;
signal \c0.tx2_transmit_N_1031\ : std_logic;
signal \c0.n1785\ : std_logic;
signal \c0.n11\ : std_logic;
signal \c0.n24_adj_1924\ : std_logic;
signal \c0.n5259_cascade_\ : std_logic;
signal \c0.n21_adj_1933\ : std_logic;
signal \c0.n16\ : std_logic;
signal \c0.n1893\ : std_logic;
signal \c0.n2008\ : std_logic;
signal \c0.n5225\ : std_logic;
signal \c0.n5198_cascade_\ : std_logic;
signal \c0.n6103\ : std_logic;
signal \c0.n28\ : std_logic;
signal \c0.n5198\ : std_logic;
signal \c0.n1918\ : std_logic;
signal \c0.n18_adj_1910\ : std_logic;
signal \c0.n17_adj_1912_cascade_\ : std_logic;
signal \c0.n12_adj_1911\ : std_logic;
signal \c0.n19_adj_1920\ : std_logic;
signal \c0.n28_adj_1902\ : std_logic;
signal \c0.n32\ : std_logic;
signal \c0.n29_adj_1905_cascade_\ : std_logic;
signal \c0.n31_adj_1904\ : std_logic;
signal \c0.n5278\ : std_logic;
signal \c0.data_in_field_134\ : std_logic;
signal \c0.n12_cascade_\ : std_logic;
signal \c0.n1880\ : std_logic;
signal \c0.n2036\ : std_logic;
signal \c0.n20_adj_1892\ : std_logic;
signal \c0.n2033\ : std_logic;
signal \c0.n10_adj_1963_cascade_\ : std_logic;
signal \c0.n5114\ : std_logic;
signal \c0.n5114_cascade_\ : std_logic;
signal \c0.n30_adj_1903\ : std_logic;
signal \c0.n5743\ : std_logic;
signal \c0.data_in_field_87\ : std_logic;
signal \c0.data_in_field_57\ : std_logic;
signal \c0.data_in_field_7\ : std_logic;
signal \c0.n5162_cascade_\ : std_logic;
signal data_in_18_1 : std_logic;
signal \c0.n1825_cascade_\ : std_logic;
signal \c0.data_in_field_133\ : std_logic;
signal \c0.data_in_field_73\ : std_logic;
signal \c0.data_in_field_35\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.data_in_field_137\ : std_logic;
signal \c0.n6_adj_1877\ : std_logic;
signal \c0.data_in_field_31\ : std_logic;
signal \c0.n28_adj_1886\ : std_logic;
signal \c0.n5222\ : std_logic;
signal \c0.n34\ : std_logic;
signal data_in_15_5 : std_logic;
signal \c0.n1686_cascade_\ : std_logic;
signal \c0.data_in_field_25\ : std_logic;
signal data_in_19_7 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n1714 : std_logic;
signal n3342 : std_logic;
signal rx_data_7 : std_logic;
signal data_in_17_1 : std_logic;
signal data_out_19_6 : std_logic;
signal data_out_18_6 : std_logic;
signal data_out_11_5 : std_logic;
signal n5176 : std_logic;
signal \c0.n1590\ : std_logic;
signal data_out_11_6 : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal data_out_10_6 : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.n3567\ : std_logic;
signal \c0.byte_transmit_counter_3\ : std_logic;
signal \c0.n5523_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal \c0.n1236\ : std_logic;
signal \c0.n5515\ : std_logic;
signal \c0.n5513_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_4\ : std_logic;
signal \tx_data_6_N_keep\ : std_logic;
signal data_out_10_5 : std_logic;
signal data_out_10_1 : std_logic;
signal data_out_10_3 : std_logic;
signal n5132 : std_logic;
signal \c0.n5839_cascade_\ : std_logic;
signal \c0.n5833_cascade_\ : std_logic;
signal \c0.n5417_cascade_\ : std_logic;
signal \c0.n5414\ : std_logic;
signal \c0.n5827\ : std_logic;
signal \c0.n5683_cascade_\ : std_logic;
signal \c0.n5695\ : std_logic;
signal \c0.n5480_cascade_\ : std_logic;
signal \c0.n5483\ : std_logic;
signal \c0.n5677_cascade_\ : std_logic;
signal \c0.n5680\ : std_logic;
signal data_in_18_5 : std_logic;
signal \c0.n24_adj_1895\ : std_logic;
signal rx_data_0 : std_logic;
signal data_in_19_0 : std_logic;
signal \c0.n5429\ : std_logic;
signal \c0.n5791\ : std_logic;
signal \c0.n5432\ : std_logic;
signal \c0.data_in_field_30\ : std_logic;
signal \c0.data_in_field_13\ : std_logic;
signal \c0.n5393\ : std_logic;
signal data_in_14_7 : std_logic;
signal \c0.n10_adj_1898\ : std_logic;
signal \c0.data_in_field_69\ : std_logic;
signal \c0.n5159\ : std_logic;
signal \c0.data_in_field_99\ : std_logic;
signal \c0.n5159_cascade_\ : std_logic;
signal \c0.data_in_field_105\ : std_logic;
signal \c0.n2095_cascade_\ : std_logic;
signal \c0.n1821\ : std_logic;
signal \c0.n34_adj_1896\ : std_logic;
signal \c0.data_in_field_11\ : std_logic;
signal \c0.n5821_cascade_\ : std_logic;
signal \c0.n5423\ : std_logic;
signal \c0.data_in_field_27\ : std_logic;
signal \c0.n2080\ : std_logic;
signal \c0.n2080_cascade_\ : std_logic;
signal \c0.n5243\ : std_logic;
signal \c0.n16_adj_1922\ : std_logic;
signal \c0.n25_adj_1926\ : std_logic;
signal \c0.n1978\ : std_logic;
signal \c0.n5261\ : std_logic;
signal \c0.n5689_cascade_\ : std_logic;
signal \c0.n5366\ : std_logic;
signal \c0.n14_adj_1967\ : std_logic;
signal \c0.n5276\ : std_logic;
signal \c0.n5201\ : std_logic;
signal \c0.n5276_cascade_\ : std_logic;
signal \c0.n37\ : std_logic;
signal \c0.data_in_field_36\ : std_logic;
signal \c0.data_in_field_22\ : std_logic;
signal \c0.n2005_cascade_\ : std_logic;
signal \c0.n10_adj_1873_cascade_\ : std_logic;
signal \c0.n1825\ : std_logic;
signal \c0.data_in_field_55\ : std_logic;
signal \c0.n13_adj_1951\ : std_logic;
signal \c0.data_in_field_23\ : std_logic;
signal \c0.n6107\ : std_logic;
signal \c0.n18_adj_1891\ : std_logic;
signal \c0.n5249\ : std_logic;
signal rx_data_2 : std_logic;
signal \c0.n5255\ : std_logic;
signal data_in_1_3 : std_logic;
signal \c0.n28_adj_1954\ : std_logic;
signal \c0.n26_adj_1955\ : std_logic;
signal \c0.n25_adj_1957_cascade_\ : std_logic;
signal \c0.n4465\ : std_logic;
signal \c0.data_in_field_17\ : std_logic;
signal data_in_1_4 : std_logic;
signal data_in_11_7 : std_logic;
signal data_in_10_7 : std_logic;
signal data_in_2_7 : std_logic;
signal \c0.n27_adj_1956\ : std_logic;
signal \c0.n26_adj_1958\ : std_logic;
signal \c0.data_in_field_135\ : std_logic;
signal \c0.data_in_field_113\ : std_logic;
signal \c0.n1772\ : std_logic;
signal \c0.n5144\ : std_logic;
signal \c0.n5144_cascade_\ : std_logic;
signal \c0.n31\ : std_logic;
signal data_in_8_5 : std_logic;
signal data_in_8_7 : std_logic;
signal \c0.n5447_cascade_\ : std_logic;
signal \c0.n5755_cascade_\ : std_logic;
signal \c0.n5758\ : std_logic;
signal \c0.data_in_field_54\ : std_logic;
signal \c0.data_in_field_10\ : std_logic;
signal \c0.n5438\ : std_logic;
signal \c0.data_in_field_82\ : std_logic;
signal \c0.n5767_cascade_\ : std_logic;
signal \c0.n5444\ : std_logic;
signal \c0.n5761\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.data_in_field_117\ : std_logic;
signal \c0.n2074_cascade_\ : std_logic;
signal \c0.n10_adj_1888\ : std_logic;
signal \c0.data_in_field_95\ : std_logic;
signal \c0.n1851\ : std_logic;
signal \c0.data_in_field_96\ : std_logic;
signal \c0.n5099\ : std_logic;
signal \c0.n5162\ : std_logic;
signal \c0.n5213\ : std_logic;
signal \c0.n5099_cascade_\ : std_logic;
signal \c0.n19\ : std_logic;
signal \c0.data_in_field_104\ : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_12_0 : std_logic;
signal \c0.data_in_field_89\ : std_logic;
signal \c0.data_in_field_120\ : std_logic;
signal \c0.n23_adj_1925\ : std_logic;
signal \c0.data_in_field_83\ : std_logic;
signal \c0.n5797\ : std_logic;
signal \c0.data_in_field_19\ : std_logic;
signal \c0.n23\ : std_logic;
signal data_in_3_3 : std_logic;
signal \c0.n25_adj_1960\ : std_logic;
signal \c0.data_in_field_67\ : std_logic;
signal \c0.n5093\ : std_logic;
signal \c0.data_in_field_21\ : std_logic;
signal \c0.n5881\ : std_logic;
signal data_in_15_6 : std_logic;
signal \c0.data_in_field_29\ : std_logic;
signal \c0.n2046\ : std_logic;
signal \c0.data_in_field_85\ : std_logic;
signal \c0.n2046_cascade_\ : std_logic;
signal \c0.n5108\ : std_logic;
signal data_in_7_1 : std_logic;
signal data_in_6_1 : std_logic;
signal \c0.data_in_field_141\ : std_logic;
signal data_in_1_6 : std_logic;
signal data_in_9_7 : std_logic;
signal data_in_6_7 : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_7_5 : std_logic;
signal data_in_18_6 : std_logic;
signal data_in_17_6 : std_logic;
signal data_in_1_5 : std_logic;
signal data_in_7_7 : std_logic;
signal \c0.data_in_field_121\ : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_17_5 : std_logic;
signal data_in_16_5 : std_logic;
signal data_in_19_2 : std_logic;
signal \c0.n5779\ : std_logic;
signal data_in_13_0 : std_logic;
signal data_in_14_0 : std_logic;
signal \c0.n1929\ : std_logic;
signal \c0.data_in_field_112\ : std_logic;
signal \c0.n1929_cascade_\ : std_logic;
signal \c0.n10_adj_1870_cascade_\ : std_logic;
signal \c0.n5204\ : std_logic;
signal \c0.data_in_field_28\ : std_logic;
signal \c0.data_in_field_20\ : std_logic;
signal \c0.data_in_field_12\ : std_logic;
signal \c0.n5851_cascade_\ : std_logic;
signal \c0.n5408\ : std_logic;
signal \c0.n5267\ : std_logic;
signal \c0.n5905\ : std_logic;
signal \c0.n2074\ : std_logic;
signal data_in_19_5 : std_logic;
signal \c0.n22_adj_1914\ : std_logic;
signal \c0.data_in_field_139\ : std_logic;
signal \c0.n1947_cascade_\ : std_logic;
signal \c0.n10\ : std_logic;
signal \c0.data_in_field_51\ : std_logic;
signal \c0.n1922\ : std_logic;
signal \c0.data_in_field_75\ : std_logic;
signal \c0.n5474\ : std_logic;
signal \c0.n26_adj_1884\ : std_logic;
signal \c0.data_in_field_98\ : std_logic;
signal data_in_12_7 : std_logic;
signal \c0.data_in_field_103\ : std_logic;
signal \c0.data_in_field_61\ : std_logic;
signal \c0.n5875_cascade_\ : std_logic;
signal \c0.data_in_field_37\ : std_logic;
signal \c0.n5396\ : std_logic;
signal \c0.data_in_field_53\ : std_logic;
signal \c0.data_in_field_88\ : std_logic;
signal \c0.data_in_field_124\ : std_logic;
signal \c0.n1944\ : std_logic;
signal \c0.n1944_cascade_\ : std_logic;
signal \c0.n20_cascade_\ : std_logic;
signal \c0.data_in_field_43\ : std_logic;
signal \c0.n24\ : std_logic;
signal data_in_4_7 : std_logic;
signal \c0.data_in_field_39\ : std_logic;
signal \c0.data_in_field_5\ : std_logic;
signal \c0.data_in_field_79\ : std_logic;
signal \c0.data_in_field_77\ : std_logic;
signal \c0.n10_adj_1871_cascade_\ : std_logic;
signal \c0.n5234\ : std_logic;
signal \c0.n1975\ : std_logic;
signal \c0.data_in_field_38\ : std_logic;
signal data_in_12_1 : std_logic;
signal \c0.n2062\ : std_logic;
signal \c0.n1830\ : std_logic;
signal \c0.n5141\ : std_logic;
signal \c0.data_in_field_106\ : std_logic;
signal data_in_13_7 : std_logic;
signal \c0.data_in_field_111\ : std_logic;
signal \c0.data_in_field_143\ : std_logic;
signal data_in_16_7 : std_logic;
signal data_in_18_7 : std_logic;
signal data_in_17_7 : std_logic;
signal \c0.data_in_field_49\ : std_logic;
signal \c0.n2092_cascade_\ : std_logic;
signal \c0.n2043\ : std_logic;
signal \c0.n5246\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.data_in_field_9\ : std_logic;
signal \c0.n5749\ : std_logic;
signal \c0.data_in_field_1\ : std_logic;
signal \c0.n5453\ : std_logic;
signal \c0.data_in_field_59\ : std_logic;
signal data_in_6_6 : std_logic;
signal data_in_13_4 : std_logic;
signal data_in_2_4 : std_logic;
signal \c0.data_in_field_115\ : std_logic;
signal data_in_9_1 : std_logic;
signal data_in_7_6 : std_logic;
signal data_in_10_4 : std_logic;
signal data_in_10_3 : std_logic;
signal data_in_9_3 : std_logic;
signal \c0.n26_adj_1878\ : std_logic;
signal data_in_0_4 : std_logic;
signal \c0.data_in_field_68\ : std_logic;
signal \c0.n5105\ : std_logic;
signal \c0.n5111\ : std_logic;
signal \c0.n35\ : std_logic;
signal data_in_16_3 : std_logic;
signal data_in_18_4 : std_logic;
signal data_in_17_4 : std_logic;
signal \c0.data_in_field_63\ : std_logic;
signal \c0.data_in_field_62\ : std_logic;
signal \c0.n1795_cascade_\ : std_logic;
signal \c0.n6097\ : std_logic;
signal data_in_6_3 : std_logic;
signal data_in_5_3 : std_logic;
signal \c0.data_in_field_142\ : std_logic;
signal \c0.n1795\ : std_logic;
signal \c0.n11_adj_1913\ : std_logic;
signal data_in_11_4 : std_logic;
signal \c0.data_in_field_92\ : std_logic;
signal data_in_11_5 : std_logic;
signal \c0.data_in_field_93\ : std_logic;
signal \c0.n5707\ : std_logic;
signal \c0.n1838\ : std_logic;
signal data_in_5_0 : std_logic;
signal \c0.n6_adj_1876_cascade_\ : std_logic;
signal \c0.data_in_field_132\ : std_logic;
signal \c0.n5129\ : std_logic;
signal \c0.n6_adj_1874\ : std_logic;
signal data_in_0_0 : std_logic;
signal \c0.data_in_field_0\ : std_logic;
signal \c0.data_in_field_90\ : std_logic;
signal \c0.n22_adj_1935\ : std_logic;
signal data_in_5_6 : std_logic;
signal \c0.data_in_field_2\ : std_logic;
signal \c0.data_in_field_108\ : std_logic;
signal \c0.n5102\ : std_logic;
signal data_in_5_7 : std_logic;
signal \c0.data_in_field_47\ : std_logic;
signal data_in_15_7 : std_logic;
signal \c0.data_in_field_127\ : std_logic;
signal data_in_16_0 : std_logic;
signal data_in_1_7 : std_logic;
signal data_in_10_5 : std_logic;
signal data_in_9_5 : std_logic;
signal data_in_0_5 : std_logic;
signal data_in_1_2 : std_logic;
signal data_in_6_5 : std_logic;
signal data_in_4_6 : std_logic;
signal data_in_6_0 : std_logic;
signal \c0.data_in_field_60\ : std_logic;
signal \c0.n6_adj_1875\ : std_logic;
signal data_in_3_5 : std_logic;
signal data_in_3_4 : std_logic;
signal data_in_2_6 : std_logic;
signal data_in_3_6 : std_logic;
signal \c0.n28_adj_1953_cascade_\ : std_logic;
signal \c0.n22_adj_1952\ : std_logic;
signal \c0.n30_adj_1959\ : std_logic;
signal data_in_4_5 : std_logic;
signal data_in_8_0 : std_logic;
signal \c0.data_in_field_58\ : std_logic;
signal \c0.n5773_cascade_\ : std_logic;
signal \c0.data_in_field_34\ : std_logic;
signal \c0.n5441\ : std_logic;
signal \c0.n5477\ : std_logic;
signal data_in_16_4 : std_logic;
signal data_in_15_4 : std_logic;
signal data_in_8_6 : std_logic;
signal data_in_11_1 : std_logic;
signal data_in_10_1 : std_logic;
signal data_in_11_0 : std_logic;
signal \c0.data_in_field_14\ : std_logic;
signal \c0.n5911\ : std_logic;
signal \c0.data_in_field_6\ : std_logic;
signal \c0.data_in_field_138\ : std_logic;
signal \c0.data_in_field_130\ : std_logic;
signal \c0.n5123\ : std_logic;
signal \c0.n5123_cascade_\ : std_logic;
signal \c0.n5231\ : std_logic;
signal data_in_13_2 : std_logic;
signal data_in_12_2 : std_logic;
signal \c0.data_in_field_64\ : std_logic;
signal \c0.n5179\ : std_logic;
signal \c0.data_in_field_46\ : std_logic;
signal \c0.data_in_field_4\ : std_logic;
signal \c0.n1767_cascade_\ : std_logic;
signal \c0.n1899\ : std_logic;
signal \c0.n5126\ : std_logic;
signal \c0.data_in_field_140\ : std_logic;
signal \c0.n5126_cascade_\ : std_logic;
signal \c0.data_in_field_125\ : std_logic;
signal \c0.n20_adj_1899\ : std_logic;
signal data_in_14_6 : std_logic;
signal \c0.n10_adj_1872\ : std_logic;
signal data_in_12_4 : std_logic;
signal \c0.data_in_field_100\ : std_logic;
signal \c0.data_in_field_40\ : std_logic;
signal \c0.data_in_field_128\ : std_logic;
signal \c0.data_in_field_16\ : std_logic;
signal \c0.data_in_field_72\ : std_logic;
signal \c0.n5188\ : std_logic;
signal \c0.n5138_cascade_\ : std_logic;
signal \c0.n15_adj_1968\ : std_logic;
signal data_in_3_2 : std_logic;
signal \c0.data_in_field_26\ : std_logic;
signal data_in_4_1 : std_logic;
signal \c0.data_in_field_33\ : std_logic;
signal data_in_2_2 : std_logic;
signal \c0.data_in_field_18\ : std_logic;
signal \c0.n6\ : std_logic;
signal data_in_4_0 : std_logic;
signal \c0.data_in_field_32\ : std_logic;
signal data_in_13_6 : std_logic;
signal n5332 : std_logic;
signal \n5331_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal \c0.data_in_field_97\ : std_logic;
signal \c0.n1972\ : std_logic;
signal data_in_9_4 : std_logic;
signal \c0.data_in_field_76\ : std_logic;
signal data_in_0_1 : std_logic;
signal data_in_5_5 : std_logic;
signal \c0.data_in_field_45\ : std_logic;
signal data_in_9_0 : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_1_1 : std_logic;
signal \c0.data_in_field_48\ : std_logic;
signal \c0.n5701\ : std_logic;
signal data_in_4_4 : std_logic;
signal data_in_6_4 : std_logic;
signal data_in_7_2 : std_logic;
signal data_in_10_6 : std_logic;
signal data_in_9_6 : std_logic;
signal data_in_10_0 : std_logic;
signal \c0.data_in_field_80\ : std_logic;
signal data_in_8_2 : std_logic;
signal data_in_14_2 : std_logic;
signal \c0.data_in_field_114\ : std_logic;
signal data_in_4_2 : std_logic;
signal \c0.data_in_field_66\ : std_logic;
signal \c0.data_in_field_84\ : std_logic;
signal \c0.n1969\ : std_logic;
signal \c0.n25\ : std_logic;
signal data_in_5_2 : std_logic;
signal \c0.data_in_field_42\ : std_logic;
signal \c0.data_in_field_107\ : std_logic;
signal \c0.data_in_field_15\ : std_logic;
signal \c0.n20_adj_1916\ : std_logic;
signal data_in_8_1 : std_logic;
signal \c0.data_in_field_65\ : std_logic;
signal data_in_16_1 : std_logic;
signal data_in_15_1 : std_logic;
signal data_in_14_4 : std_logic;
signal \c0.data_in_field_116\ : std_logic;
signal \c0.n1815\ : std_logic;
signal \c0.n1815_cascade_\ : std_logic;
signal \c0.data_in_field_52\ : std_logic;
signal \c0.n27\ : std_logic;
signal data_in_14_1 : std_logic;
signal data_in_13_1 : std_logic;
signal data_in_7_0 : std_logic;
signal \c0.data_in_field_56\ : std_logic;
signal \c0.data_in_field_129\ : std_logic;
signal \c0.n15_adj_1923\ : std_logic;
signal data_in_6_2 : std_logic;
signal \c0.data_in_field_50\ : std_logic;
signal \c0.data_in_field_8\ : std_logic;
signal data_in_5_4 : std_logic;
signal \c0.data_in_field_44\ : std_logic;
signal \c0.n1962\ : std_logic;
signal data_in_3_0 : std_logic;
signal \c0.data_in_field_24\ : std_logic;
signal data_in_2_0 : std_logic;
signal data_in_1_0 : std_logic;
signal data_in_15_3 : std_logic;
signal \c0.data_in_field_123\ : std_logic;
signal data_in_12_6 : std_logic;
signal data_in_11_6 : std_logic;
signal data_in_18_2 : std_logic;
signal \c0.data_in_field_74\ : std_logic;
signal \c0.data_in_field_136\ : std_logic;
signal data_in_15_2 : std_logic;
signal \c0.data_in_field_122\ : std_logic;
signal data_in_14_3 : std_logic;
signal data_in_13_3 : std_logic;
signal data_in_12_3 : std_logic;
signal data_in_11_3 : std_logic;
signal \c0.data_in_field_91\ : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.data_in_field_3\ : std_logic;
signal data_in_11_2 : std_logic;
signal data_in_10_2 : std_logic;
signal data_in_9_2 : std_logic;
signal data_in_8_3 : std_logic;
signal data_in_7_3 : std_logic;
signal data_in_18_0 : std_logic;
signal data_in_17_0 : std_logic;
signal \c0.data_in_field_118\ : std_logic;
signal \c0.data_in_field_126\ : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal \c0.data_in_field_86\ : std_logic;
signal \c0.data_in_field_94\ : std_logic;
signal \c0.data_in_field_70\ : std_logic;
signal \c0.n5899_cascade_\ : std_logic;
signal \c0.data_in_field_78\ : std_logic;
signal \c0.n5893\ : std_logic;
signal \c0.data_in_field_102\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.data_in_field_110\ : std_logic;
signal \c0.n5384\ : std_logic;
signal \c0.n5387_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.n5378\ : std_logic;
signal \c0.n5381\ : std_logic;
signal \c0.n5887_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.n5890\ : std_logic;
signal \c0.n5219\ : std_logic;
signal \c0.n5138\ : std_logic;
signal \c0.n1896\ : std_logic;
signal data_in_8_4 : std_logic;
signal data_in_7_4 : std_logic;
signal rx_data_ready : std_logic;
signal data_in_17_2 : std_logic;
signal data_in_16_2 : std_logic;
signal n26 : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal n25 : std_logic;
signal n4437 : std_logic;
signal n24 : std_logic;
signal n4438 : std_logic;
signal n23 : std_logic;
signal n4439 : std_logic;
signal n22 : std_logic;
signal n4440 : std_logic;
signal n21 : std_logic;
signal n4441 : std_logic;
signal n20 : std_logic;
signal n4442 : std_logic;
signal n19 : std_logic;
signal n4443 : std_logic;
signal n4444 : std_logic;
signal n18 : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal n17 : std_logic;
signal n4445 : std_logic;
signal n16 : std_logic;
signal n4446 : std_logic;
signal n15 : std_logic;
signal n4447 : std_logic;
signal n14 : std_logic;
signal n4448 : std_logic;
signal n13 : std_logic;
signal n4449 : std_logic;
signal n12 : std_logic;
signal n4450 : std_logic;
signal n11 : std_logic;
signal n4451 : std_logic;
signal n4452 : std_logic;
signal n10 : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal n9 : std_logic;
signal n4453 : std_logic;
signal n8_adj_1989 : std_logic;
signal n4454 : std_logic;
signal n7 : std_logic;
signal n4455 : std_logic;
signal n6 : std_logic;
signal n4456 : std_logic;
signal blink_counter_21 : std_logic;
signal n4457 : std_logic;
signal blink_counter_22 : std_logic;
signal n4458 : std_logic;
signal blink_counter_23 : std_logic;
signal n4459 : std_logic;
signal n4460 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal n4461 : std_logic;
signal blink_counter_25 : std_logic;
signal data_in_19_4 : std_logic;
signal \c0.FRAME_MATCHER_wait_for_transmission\ : std_logic;
signal \c0.n1686\ : std_logic;
signal \c0.data_in_frame_19_4\ : std_logic;
signal \CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37526\,
            DIN => \N__37525\,
            DOUT => \N__37524\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37526\,
            PADOUT => \N__37525\,
            PADIN => \N__37524\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29815\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37517\,
            DIN => \N__37516\,
            DOUT => \N__37515\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37517\,
            PADOUT => \N__37516\,
            PADIN => \N__37515\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__37508\,
            DIN => \N__37507\,
            DOUT => \N__37506\,
            PACKAGEPIN => PIN_2
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37508\,
            PADOUT => \N__37507\,
            PADIN => \N__37506\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__35351\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__37499\,
            DIN => \N__37498\,
            DOUT => \N__37497\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37499\,
            PADOUT => \N__37498\,
            PADIN => \N__37497\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12276\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__12256\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__37490\,
            DIN => \N__37489\,
            DOUT => \N__37488\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37490\,
            PADOUT => \N__37489\,
            PADIN => \N__37488\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__16890\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__14842\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37481\,
            DIN => \N__37480\,
            DOUT => \N__37479\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37481\,
            PADOUT => \N__37480\,
            PADIN => \N__37479\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__9468\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37456\
        );

    \I__9467\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37456\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37453\
        );

    \I__9465\ : Span4Mux_v
    port map (
            O => \N__37453\,
            I => \N__37449\
        );

    \I__9464\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37446\
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__37449\,
            I => blink_counter_21
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__37446\,
            I => blink_counter_21
        );

    \I__9461\ : InMux
    port map (
            O => \N__37441\,
            I => n4457
        );

    \I__9460\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37432\
        );

    \I__9459\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37432\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__37432\,
            I => \N__37429\
        );

    \I__9457\ : Span4Mux_v
    port map (
            O => \N__37429\,
            I => \N__37425\
        );

    \I__9456\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37422\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__37425\,
            I => blink_counter_22
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__37422\,
            I => blink_counter_22
        );

    \I__9453\ : InMux
    port map (
            O => \N__37417\,
            I => n4458
        );

    \I__9452\ : CascadeMux
    port map (
            O => \N__37414\,
            I => \N__37410\
        );

    \I__9451\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37405\
        );

    \I__9450\ : InMux
    port map (
            O => \N__37410\,
            I => \N__37405\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__37405\,
            I => \N__37402\
        );

    \I__9448\ : Span4Mux_h
    port map (
            O => \N__37402\,
            I => \N__37398\
        );

    \I__9447\ : InMux
    port map (
            O => \N__37401\,
            I => \N__37395\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__37398\,
            I => blink_counter_23
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__37395\,
            I => blink_counter_23
        );

    \I__9444\ : InMux
    port map (
            O => \N__37390\,
            I => n4459
        );

    \I__9443\ : CascadeMux
    port map (
            O => \N__37387\,
            I => \N__37384\
        );

    \I__9442\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37378\
        );

    \I__9441\ : InMux
    port map (
            O => \N__37383\,
            I => \N__37378\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__37378\,
            I => \N__37375\
        );

    \I__9439\ : Span4Mux_v
    port map (
            O => \N__37375\,
            I => \N__37371\
        );

    \I__9438\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37368\
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__37371\,
            I => blink_counter_24
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__37368\,
            I => blink_counter_24
        );

    \I__9435\ : InMux
    port map (
            O => \N__37363\,
            I => \bfn_15_28_0_\
        );

    \I__9434\ : InMux
    port map (
            O => \N__37360\,
            I => n4461
        );

    \I__9433\ : InMux
    port map (
            O => \N__37357\,
            I => \N__37354\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__37354\,
            I => \N__37351\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__37351\,
            I => \N__37347\
        );

    \I__9430\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37344\
        );

    \I__9429\ : Odrv4
    port map (
            O => \N__37347\,
            I => blink_counter_25
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__37344\,
            I => blink_counter_25
        );

    \I__9427\ : InMux
    port map (
            O => \N__37339\,
            I => \N__37335\
        );

    \I__9426\ : CascadeMux
    port map (
            O => \N__37338\,
            I => \N__37331\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__37335\,
            I => \N__37328\
        );

    \I__9424\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37325\
        );

    \I__9423\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37322\
        );

    \I__9422\ : Span12Mux_s7_v
    port map (
            O => \N__37328\,
            I => \N__37319\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__37325\,
            I => \N__37316\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__37322\,
            I => \N__37312\
        );

    \I__9419\ : Span12Mux_h
    port map (
            O => \N__37319\,
            I => \N__37309\
        );

    \I__9418\ : Span4Mux_h
    port map (
            O => \N__37316\,
            I => \N__37306\
        );

    \I__9417\ : InMux
    port map (
            O => \N__37315\,
            I => \N__37303\
        );

    \I__9416\ : Span12Mux_v
    port map (
            O => \N__37312\,
            I => \N__37300\
        );

    \I__9415\ : Odrv12
    port map (
            O => \N__37309\,
            I => data_in_19_4
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__37306\,
            I => data_in_19_4
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__37303\,
            I => data_in_19_4
        );

    \I__9412\ : Odrv12
    port map (
            O => \N__37300\,
            I => data_in_19_4
        );

    \I__9411\ : CascadeMux
    port map (
            O => \N__37291\,
            I => \N__37286\
        );

    \I__9410\ : CascadeMux
    port map (
            O => \N__37290\,
            I => \N__37282\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__37289\,
            I => \N__37262\
        );

    \I__9408\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37258\
        );

    \I__9407\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37251\
        );

    \I__9406\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37251\
        );

    \I__9405\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37251\
        );

    \I__9404\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37243\
        );

    \I__9403\ : InMux
    port map (
            O => \N__37279\,
            I => \N__37243\
        );

    \I__9402\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37243\
        );

    \I__9401\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37232\
        );

    \I__9400\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37232\
        );

    \I__9399\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37232\
        );

    \I__9398\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37232\
        );

    \I__9397\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37232\
        );

    \I__9396\ : CascadeMux
    port map (
            O => \N__37272\,
            I => \N__37223\
        );

    \I__9395\ : CascadeMux
    port map (
            O => \N__37271\,
            I => \N__37219\
        );

    \I__9394\ : CascadeMux
    port map (
            O => \N__37270\,
            I => \N__37215\
        );

    \I__9393\ : CascadeMux
    port map (
            O => \N__37269\,
            I => \N__37209\
        );

    \I__9392\ : CascadeMux
    port map (
            O => \N__37268\,
            I => \N__37204\
        );

    \I__9391\ : CascadeMux
    port map (
            O => \N__37267\,
            I => \N__37196\
        );

    \I__9390\ : CascadeMux
    port map (
            O => \N__37266\,
            I => \N__37191\
        );

    \I__9389\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37181\
        );

    \I__9388\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37176\
        );

    \I__9387\ : InMux
    port map (
            O => \N__37261\,
            I => \N__37176\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__37258\,
            I => \N__37171\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37171\
        );

    \I__9384\ : CascadeMux
    port map (
            O => \N__37250\,
            I => \N__37168\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37158\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__37232\,
            I => \N__37155\
        );

    \I__9381\ : CascadeMux
    port map (
            O => \N__37231\,
            I => \N__37139\
        );

    \I__9380\ : CascadeMux
    port map (
            O => \N__37230\,
            I => \N__37136\
        );

    \I__9379\ : CascadeMux
    port map (
            O => \N__37229\,
            I => \N__37133\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__37228\,
            I => \N__37129\
        );

    \I__9377\ : CascadeMux
    port map (
            O => \N__37227\,
            I => \N__37120\
        );

    \I__9376\ : CascadeMux
    port map (
            O => \N__37226\,
            I => \N__37117\
        );

    \I__9375\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37111\
        );

    \I__9374\ : InMux
    port map (
            O => \N__37222\,
            I => \N__37111\
        );

    \I__9373\ : InMux
    port map (
            O => \N__37219\,
            I => \N__37106\
        );

    \I__9372\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37106\
        );

    \I__9371\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37099\
        );

    \I__9370\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37099\
        );

    \I__9369\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37099\
        );

    \I__9368\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37090\
        );

    \I__9367\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37090\
        );

    \I__9366\ : InMux
    port map (
            O => \N__37208\,
            I => \N__37090\
        );

    \I__9365\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37090\
        );

    \I__9364\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37083\
        );

    \I__9363\ : CascadeMux
    port map (
            O => \N__37203\,
            I => \N__37080\
        );

    \I__9362\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37074\
        );

    \I__9361\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37074\
        );

    \I__9360\ : CascadeMux
    port map (
            O => \N__37200\,
            I => \N__37071\
        );

    \I__9359\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37061\
        );

    \I__9358\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37061\
        );

    \I__9357\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37061\
        );

    \I__9356\ : CascadeMux
    port map (
            O => \N__37194\,
            I => \N__37055\
        );

    \I__9355\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37050\
        );

    \I__9354\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37045\
        );

    \I__9353\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37045\
        );

    \I__9352\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37042\
        );

    \I__9351\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37033\
        );

    \I__9350\ : InMux
    port map (
            O => \N__37186\,
            I => \N__37033\
        );

    \I__9349\ : InMux
    port map (
            O => \N__37185\,
            I => \N__37033\
        );

    \I__9348\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37033\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37026\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__37176\,
            I => \N__37026\
        );

    \I__9345\ : Span4Mux_h
    port map (
            O => \N__37171\,
            I => \N__37026\
        );

    \I__9344\ : InMux
    port map (
            O => \N__37168\,
            I => \N__37021\
        );

    \I__9343\ : InMux
    port map (
            O => \N__37167\,
            I => \N__37021\
        );

    \I__9342\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37010\
        );

    \I__9341\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37010\
        );

    \I__9340\ : InMux
    port map (
            O => \N__37164\,
            I => \N__37010\
        );

    \I__9339\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37010\
        );

    \I__9338\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37010\
        );

    \I__9337\ : CascadeMux
    port map (
            O => \N__37161\,
            I => \N__36993\
        );

    \I__9336\ : Span4Mux_v
    port map (
            O => \N__37158\,
            I => \N__36984\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__37155\,
            I => \N__36984\
        );

    \I__9334\ : InMux
    port map (
            O => \N__37154\,
            I => \N__36977\
        );

    \I__9333\ : InMux
    port map (
            O => \N__37153\,
            I => \N__36977\
        );

    \I__9332\ : InMux
    port map (
            O => \N__37152\,
            I => \N__36977\
        );

    \I__9331\ : InMux
    port map (
            O => \N__37151\,
            I => \N__36966\
        );

    \I__9330\ : InMux
    port map (
            O => \N__37150\,
            I => \N__36966\
        );

    \I__9329\ : InMux
    port map (
            O => \N__37149\,
            I => \N__36966\
        );

    \I__9328\ : InMux
    port map (
            O => \N__37148\,
            I => \N__36966\
        );

    \I__9327\ : InMux
    port map (
            O => \N__37147\,
            I => \N__36966\
        );

    \I__9326\ : InMux
    port map (
            O => \N__37146\,
            I => \N__36957\
        );

    \I__9325\ : InMux
    port map (
            O => \N__37145\,
            I => \N__36957\
        );

    \I__9324\ : InMux
    port map (
            O => \N__37144\,
            I => \N__36957\
        );

    \I__9323\ : InMux
    port map (
            O => \N__37143\,
            I => \N__36957\
        );

    \I__9322\ : InMux
    port map (
            O => \N__37142\,
            I => \N__36945\
        );

    \I__9321\ : InMux
    port map (
            O => \N__37139\,
            I => \N__36945\
        );

    \I__9320\ : InMux
    port map (
            O => \N__37136\,
            I => \N__36938\
        );

    \I__9319\ : InMux
    port map (
            O => \N__37133\,
            I => \N__36938\
        );

    \I__9318\ : InMux
    port map (
            O => \N__37132\,
            I => \N__36938\
        );

    \I__9317\ : InMux
    port map (
            O => \N__37129\,
            I => \N__36934\
        );

    \I__9316\ : InMux
    port map (
            O => \N__37128\,
            I => \N__36927\
        );

    \I__9315\ : InMux
    port map (
            O => \N__37127\,
            I => \N__36927\
        );

    \I__9314\ : InMux
    port map (
            O => \N__37126\,
            I => \N__36927\
        );

    \I__9313\ : InMux
    port map (
            O => \N__37125\,
            I => \N__36922\
        );

    \I__9312\ : InMux
    port map (
            O => \N__37124\,
            I => \N__36922\
        );

    \I__9311\ : InMux
    port map (
            O => \N__37123\,
            I => \N__36913\
        );

    \I__9310\ : InMux
    port map (
            O => \N__37120\,
            I => \N__36913\
        );

    \I__9309\ : InMux
    port map (
            O => \N__37117\,
            I => \N__36913\
        );

    \I__9308\ : InMux
    port map (
            O => \N__37116\,
            I => \N__36913\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__37111\,
            I => \N__36910\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__36907\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__37099\,
            I => \N__36902\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__37090\,
            I => \N__36902\
        );

    \I__9303\ : InMux
    port map (
            O => \N__37089\,
            I => \N__36895\
        );

    \I__9302\ : InMux
    port map (
            O => \N__37088\,
            I => \N__36895\
        );

    \I__9301\ : InMux
    port map (
            O => \N__37087\,
            I => \N__36895\
        );

    \I__9300\ : CascadeMux
    port map (
            O => \N__37086\,
            I => \N__36890\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__37083\,
            I => \N__36885\
        );

    \I__9298\ : InMux
    port map (
            O => \N__37080\,
            I => \N__36882\
        );

    \I__9297\ : CascadeMux
    port map (
            O => \N__37079\,
            I => \N__36877\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__37074\,
            I => \N__36874\
        );

    \I__9295\ : InMux
    port map (
            O => \N__37071\,
            I => \N__36865\
        );

    \I__9294\ : InMux
    port map (
            O => \N__37070\,
            I => \N__36865\
        );

    \I__9293\ : InMux
    port map (
            O => \N__37069\,
            I => \N__36865\
        );

    \I__9292\ : InMux
    port map (
            O => \N__37068\,
            I => \N__36865\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__37061\,
            I => \N__36862\
        );

    \I__9290\ : InMux
    port map (
            O => \N__37060\,
            I => \N__36857\
        );

    \I__9289\ : InMux
    port map (
            O => \N__37059\,
            I => \N__36857\
        );

    \I__9288\ : InMux
    port map (
            O => \N__37058\,
            I => \N__36854\
        );

    \I__9287\ : InMux
    port map (
            O => \N__37055\,
            I => \N__36849\
        );

    \I__9286\ : InMux
    port map (
            O => \N__37054\,
            I => \N__36849\
        );

    \I__9285\ : InMux
    port map (
            O => \N__37053\,
            I => \N__36842\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__37050\,
            I => \N__36837\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__37045\,
            I => \N__36837\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__37042\,
            I => \N__36826\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__36826\
        );

    \I__9280\ : Span4Mux_h
    port map (
            O => \N__37026\,
            I => \N__36826\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__37021\,
            I => \N__36826\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__37010\,
            I => \N__36826\
        );

    \I__9277\ : InMux
    port map (
            O => \N__37009\,
            I => \N__36823\
        );

    \I__9276\ : InMux
    port map (
            O => \N__37008\,
            I => \N__36816\
        );

    \I__9275\ : InMux
    port map (
            O => \N__37007\,
            I => \N__36816\
        );

    \I__9274\ : InMux
    port map (
            O => \N__37006\,
            I => \N__36816\
        );

    \I__9273\ : CascadeMux
    port map (
            O => \N__37005\,
            I => \N__36811\
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__37004\,
            I => \N__36808\
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__37003\,
            I => \N__36799\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__37002\,
            I => \N__36795\
        );

    \I__9269\ : CascadeMux
    port map (
            O => \N__37001\,
            I => \N__36792\
        );

    \I__9268\ : CascadeMux
    port map (
            O => \N__37000\,
            I => \N__36788\
        );

    \I__9267\ : CascadeMux
    port map (
            O => \N__36999\,
            I => \N__36782\
        );

    \I__9266\ : InMux
    port map (
            O => \N__36998\,
            I => \N__36775\
        );

    \I__9265\ : InMux
    port map (
            O => \N__36997\,
            I => \N__36775\
        );

    \I__9264\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36775\
        );

    \I__9263\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36766\
        );

    \I__9262\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36766\
        );

    \I__9261\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36766\
        );

    \I__9260\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36766\
        );

    \I__9259\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36763\
        );

    \I__9258\ : Span4Mux_v
    port map (
            O => \N__36984\,
            I => \N__36760\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36757\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__36966\,
            I => \N__36752\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__36957\,
            I => \N__36752\
        );

    \I__9254\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36745\
        );

    \I__9253\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36745\
        );

    \I__9252\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36745\
        );

    \I__9251\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36742\
        );

    \I__9250\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36739\
        );

    \I__9249\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36734\
        );

    \I__9248\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36734\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__36945\,
            I => \N__36729\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__36938\,
            I => \N__36729\
        );

    \I__9245\ : InMux
    port map (
            O => \N__36937\,
            I => \N__36726\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__36934\,
            I => \N__36723\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__36927\,
            I => \N__36716\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__36922\,
            I => \N__36716\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__36913\,
            I => \N__36716\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__36910\,
            I => \N__36711\
        );

    \I__9239\ : Span4Mux_h
    port map (
            O => \N__36907\,
            I => \N__36711\
        );

    \I__9238\ : Span4Mux_h
    port map (
            O => \N__36902\,
            I => \N__36706\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__36895\,
            I => \N__36706\
        );

    \I__9236\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36699\
        );

    \I__9235\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36699\
        );

    \I__9234\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36692\
        );

    \I__9233\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36692\
        );

    \I__9232\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36692\
        );

    \I__9231\ : Span4Mux_s3_h
    port map (
            O => \N__36885\,
            I => \N__36686\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__36882\,
            I => \N__36686\
        );

    \I__9229\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36681\
        );

    \I__9228\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36681\
        );

    \I__9227\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36678\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__36874\,
            I => \N__36673\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36673\
        );

    \I__9224\ : Span4Mux_h
    port map (
            O => \N__36862\,
            I => \N__36666\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__36857\,
            I => \N__36666\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__36854\,
            I => \N__36666\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__36849\,
            I => \N__36663\
        );

    \I__9220\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36654\
        );

    \I__9219\ : InMux
    port map (
            O => \N__36847\,
            I => \N__36654\
        );

    \I__9218\ : InMux
    port map (
            O => \N__36846\,
            I => \N__36654\
        );

    \I__9217\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36654\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__36842\,
            I => \N__36651\
        );

    \I__9215\ : Span4Mux_h
    port map (
            O => \N__36837\,
            I => \N__36640\
        );

    \I__9214\ : Span4Mux_v
    port map (
            O => \N__36826\,
            I => \N__36640\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__36823\,
            I => \N__36640\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__36816\,
            I => \N__36640\
        );

    \I__9211\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36630\
        );

    \I__9210\ : InMux
    port map (
            O => \N__36814\,
            I => \N__36630\
        );

    \I__9209\ : InMux
    port map (
            O => \N__36811\,
            I => \N__36627\
        );

    \I__9208\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36622\
        );

    \I__9207\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36622\
        );

    \I__9206\ : InMux
    port map (
            O => \N__36806\,
            I => \N__36615\
        );

    \I__9205\ : InMux
    port map (
            O => \N__36805\,
            I => \N__36615\
        );

    \I__9204\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36615\
        );

    \I__9203\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36612\
        );

    \I__9202\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36609\
        );

    \I__9201\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36599\
        );

    \I__9200\ : InMux
    port map (
            O => \N__36798\,
            I => \N__36599\
        );

    \I__9199\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36592\
        );

    \I__9198\ : InMux
    port map (
            O => \N__36792\,
            I => \N__36592\
        );

    \I__9197\ : InMux
    port map (
            O => \N__36791\,
            I => \N__36592\
        );

    \I__9196\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36587\
        );

    \I__9195\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36587\
        );

    \I__9194\ : InMux
    port map (
            O => \N__36786\,
            I => \N__36584\
        );

    \I__9193\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36579\
        );

    \I__9192\ : InMux
    port map (
            O => \N__36782\,
            I => \N__36579\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__36775\,
            I => \N__36574\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__36766\,
            I => \N__36574\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__36763\,
            I => \N__36567\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__36760\,
            I => \N__36567\
        );

    \I__9187\ : Span4Mux_v
    port map (
            O => \N__36757\,
            I => \N__36567\
        );

    \I__9186\ : Span4Mux_s3_v
    port map (
            O => \N__36752\,
            I => \N__36562\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__36745\,
            I => \N__36562\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__36742\,
            I => \N__36557\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__36739\,
            I => \N__36557\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__36734\,
            I => \N__36542\
        );

    \I__9181\ : Span4Mux_s3_v
    port map (
            O => \N__36729\,
            I => \N__36542\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__36726\,
            I => \N__36542\
        );

    \I__9179\ : Span4Mux_h
    port map (
            O => \N__36723\,
            I => \N__36542\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__36716\,
            I => \N__36542\
        );

    \I__9177\ : Span4Mux_h
    port map (
            O => \N__36711\,
            I => \N__36542\
        );

    \I__9176\ : Span4Mux_h
    port map (
            O => \N__36706\,
            I => \N__36542\
        );

    \I__9175\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36537\
        );

    \I__9174\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36537\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__36699\,
            I => \N__36532\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__36692\,
            I => \N__36532\
        );

    \I__9171\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36529\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__36686\,
            I => \N__36524\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36524\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36513\
        );

    \I__9167\ : Span4Mux_v
    port map (
            O => \N__36673\,
            I => \N__36513\
        );

    \I__9166\ : Span4Mux_v
    port map (
            O => \N__36666\,
            I => \N__36513\
        );

    \I__9165\ : Span4Mux_v
    port map (
            O => \N__36663\,
            I => \N__36513\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__36654\,
            I => \N__36513\
        );

    \I__9163\ : Span4Mux_h
    port map (
            O => \N__36651\,
            I => \N__36510\
        );

    \I__9162\ : CascadeMux
    port map (
            O => \N__36650\,
            I => \N__36505\
        );

    \I__9161\ : CascadeMux
    port map (
            O => \N__36649\,
            I => \N__36502\
        );

    \I__9160\ : Span4Mux_v
    port map (
            O => \N__36640\,
            I => \N__36497\
        );

    \I__9159\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36491\
        );

    \I__9158\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36486\
        );

    \I__9157\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36486\
        );

    \I__9156\ : CascadeMux
    port map (
            O => \N__36636\,
            I => \N__36483\
        );

    \I__9155\ : CascadeMux
    port map (
            O => \N__36635\,
            I => \N__36479\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__36630\,
            I => \N__36466\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__36627\,
            I => \N__36466\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__36622\,
            I => \N__36466\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__36615\,
            I => \N__36466\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__36612\,
            I => \N__36466\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36466\
        );

    \I__9148\ : InMux
    port map (
            O => \N__36608\,
            I => \N__36455\
        );

    \I__9147\ : InMux
    port map (
            O => \N__36607\,
            I => \N__36455\
        );

    \I__9146\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36455\
        );

    \I__9145\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36455\
        );

    \I__9144\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36455\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__36599\,
            I => \N__36446\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__36592\,
            I => \N__36446\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__36587\,
            I => \N__36446\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__36584\,
            I => \N__36446\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__36579\,
            I => \N__36441\
        );

    \I__9138\ : Span4Mux_v
    port map (
            O => \N__36574\,
            I => \N__36441\
        );

    \I__9137\ : Span4Mux_h
    port map (
            O => \N__36567\,
            I => \N__36438\
        );

    \I__9136\ : Span4Mux_v
    port map (
            O => \N__36562\,
            I => \N__36430\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__36557\,
            I => \N__36430\
        );

    \I__9134\ : Span4Mux_v
    port map (
            O => \N__36542\,
            I => \N__36430\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__36537\,
            I => \N__36425\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__36532\,
            I => \N__36425\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__36529\,
            I => \N__36416\
        );

    \I__9130\ : Span4Mux_h
    port map (
            O => \N__36524\,
            I => \N__36416\
        );

    \I__9129\ : Span4Mux_h
    port map (
            O => \N__36513\,
            I => \N__36416\
        );

    \I__9128\ : Span4Mux_v
    port map (
            O => \N__36510\,
            I => \N__36416\
        );

    \I__9127\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36413\
        );

    \I__9126\ : InMux
    port map (
            O => \N__36508\,
            I => \N__36402\
        );

    \I__9125\ : InMux
    port map (
            O => \N__36505\,
            I => \N__36402\
        );

    \I__9124\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36402\
        );

    \I__9123\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36402\
        );

    \I__9122\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36402\
        );

    \I__9121\ : Span4Mux_h
    port map (
            O => \N__36497\,
            I => \N__36399\
        );

    \I__9120\ : InMux
    port map (
            O => \N__36496\,
            I => \N__36392\
        );

    \I__9119\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36392\
        );

    \I__9118\ : InMux
    port map (
            O => \N__36494\,
            I => \N__36392\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__36491\,
            I => \N__36387\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36387\
        );

    \I__9115\ : InMux
    port map (
            O => \N__36483\,
            I => \N__36380\
        );

    \I__9114\ : InMux
    port map (
            O => \N__36482\,
            I => \N__36380\
        );

    \I__9113\ : InMux
    port map (
            O => \N__36479\,
            I => \N__36380\
        );

    \I__9112\ : Span12Mux_h
    port map (
            O => \N__36466\,
            I => \N__36377\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__36455\,
            I => \N__36368\
        );

    \I__9110\ : Span4Mux_v
    port map (
            O => \N__36446\,
            I => \N__36368\
        );

    \I__9109\ : Span4Mux_v
    port map (
            O => \N__36441\,
            I => \N__36368\
        );

    \I__9108\ : Span4Mux_v
    port map (
            O => \N__36438\,
            I => \N__36368\
        );

    \I__9107\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36365\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__36430\,
            I => \N__36362\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__36425\,
            I => \N__36357\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__36416\,
            I => \N__36357\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__36413\,
            I => \N__36350\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__36402\,
            I => \N__36350\
        );

    \I__9101\ : Span4Mux_h
    port map (
            O => \N__36399\,
            I => \N__36350\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__36392\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9099\ : Odrv12
    port map (
            O => \N__36387\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__36380\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9097\ : Odrv12
    port map (
            O => \N__36377\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__36368\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__36365\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__36362\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__36357\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__36350\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__9091\ : CascadeMux
    port map (
            O => \N__36331\,
            I => \N__36324\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__36330\,
            I => \N__36316\
        );

    \I__9089\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36302\
        );

    \I__9088\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36302\
        );

    \I__9087\ : InMux
    port map (
            O => \N__36327\,
            I => \N__36302\
        );

    \I__9086\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36299\
        );

    \I__9085\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36294\
        );

    \I__9084\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36294\
        );

    \I__9083\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36282\
        );

    \I__9082\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36282\
        );

    \I__9081\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36282\
        );

    \I__9080\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36277\
        );

    \I__9079\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36277\
        );

    \I__9078\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36274\
        );

    \I__9077\ : CascadeMux
    port map (
            O => \N__36313\,
            I => \N__36267\
        );

    \I__9076\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36258\
        );

    \I__9075\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36244\
        );

    \I__9074\ : InMux
    port map (
            O => \N__36310\,
            I => \N__36244\
        );

    \I__9073\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36244\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__36302\,
            I => \N__36241\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__36299\,
            I => \N__36236\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36236\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__36293\,
            I => \N__36232\
        );

    \I__9068\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36219\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__36291\,
            I => \N__36212\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__36290\,
            I => \N__36209\
        );

    \I__9065\ : InMux
    port map (
            O => \N__36289\,
            I => \N__36190\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__36282\,
            I => \N__36183\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__36277\,
            I => \N__36183\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__36274\,
            I => \N__36183\
        );

    \I__9061\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36176\
        );

    \I__9060\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36176\
        );

    \I__9059\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36176\
        );

    \I__9058\ : CascadeMux
    port map (
            O => \N__36270\,
            I => \N__36164\
        );

    \I__9057\ : InMux
    port map (
            O => \N__36267\,
            I => \N__36154\
        );

    \I__9056\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36154\
        );

    \I__9055\ : InMux
    port map (
            O => \N__36265\,
            I => \N__36147\
        );

    \I__9054\ : InMux
    port map (
            O => \N__36264\,
            I => \N__36147\
        );

    \I__9053\ : InMux
    port map (
            O => \N__36263\,
            I => \N__36147\
        );

    \I__9052\ : CascadeMux
    port map (
            O => \N__36262\,
            I => \N__36143\
        );

    \I__9051\ : CascadeMux
    port map (
            O => \N__36261\,
            I => \N__36140\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__36258\,
            I => \N__36137\
        );

    \I__9049\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36130\
        );

    \I__9048\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36130\
        );

    \I__9047\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36130\
        );

    \I__9046\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36123\
        );

    \I__9045\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36123\
        );

    \I__9044\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36123\
        );

    \I__9043\ : InMux
    port map (
            O => \N__36251\,
            I => \N__36120\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__36244\,
            I => \N__36113\
        );

    \I__9041\ : Span4Mux_v
    port map (
            O => \N__36241\,
            I => \N__36113\
        );

    \I__9040\ : Span4Mux_v
    port map (
            O => \N__36236\,
            I => \N__36113\
        );

    \I__9039\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36102\
        );

    \I__9038\ : InMux
    port map (
            O => \N__36232\,
            I => \N__36102\
        );

    \I__9037\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36102\
        );

    \I__9036\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36102\
        );

    \I__9035\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36102\
        );

    \I__9034\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36096\
        );

    \I__9033\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36096\
        );

    \I__9032\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36091\
        );

    \I__9031\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36091\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__36224\,
            I => \N__36088\
        );

    \I__9029\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36076\
        );

    \I__9028\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36076\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36073\
        );

    \I__9026\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36064\
        );

    \I__9025\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36064\
        );

    \I__9024\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36064\
        );

    \I__9023\ : InMux
    port map (
            O => \N__36215\,
            I => \N__36064\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36050\
        );

    \I__9021\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36050\
        );

    \I__9020\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36050\
        );

    \I__9019\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36045\
        );

    \I__9018\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36045\
        );

    \I__9017\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36042\
        );

    \I__9016\ : CascadeMux
    port map (
            O => \N__36204\,
            I => \N__36027\
        );

    \I__9015\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36019\
        );

    \I__9014\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36019\
        );

    \I__9013\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36014\
        );

    \I__9012\ : CascadeMux
    port map (
            O => \N__36200\,
            I => \N__36007\
        );

    \I__9011\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36000\
        );

    \I__9010\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36000\
        );

    \I__9009\ : InMux
    port map (
            O => \N__36197\,
            I => \N__35997\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__35993\
        );

    \I__9007\ : InMux
    port map (
            O => \N__36195\,
            I => \N__35981\
        );

    \I__9006\ : InMux
    port map (
            O => \N__36194\,
            I => \N__35981\
        );

    \I__9005\ : CascadeMux
    port map (
            O => \N__36193\,
            I => \N__35978\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__36190\,
            I => \N__35975\
        );

    \I__9003\ : Span4Mux_v
    port map (
            O => \N__36183\,
            I => \N__35970\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__36176\,
            I => \N__35970\
        );

    \I__9001\ : InMux
    port map (
            O => \N__36175\,
            I => \N__35967\
        );

    \I__9000\ : InMux
    port map (
            O => \N__36174\,
            I => \N__35961\
        );

    \I__8999\ : InMux
    port map (
            O => \N__36173\,
            I => \N__35956\
        );

    \I__8998\ : InMux
    port map (
            O => \N__36172\,
            I => \N__35956\
        );

    \I__8997\ : InMux
    port map (
            O => \N__36171\,
            I => \N__35951\
        );

    \I__8996\ : InMux
    port map (
            O => \N__36170\,
            I => \N__35951\
        );

    \I__8995\ : InMux
    port map (
            O => \N__36169\,
            I => \N__35944\
        );

    \I__8994\ : InMux
    port map (
            O => \N__36168\,
            I => \N__35944\
        );

    \I__8993\ : InMux
    port map (
            O => \N__36167\,
            I => \N__35944\
        );

    \I__8992\ : InMux
    port map (
            O => \N__36164\,
            I => \N__35939\
        );

    \I__8991\ : InMux
    port map (
            O => \N__36163\,
            I => \N__35939\
        );

    \I__8990\ : InMux
    port map (
            O => \N__36162\,
            I => \N__35930\
        );

    \I__8989\ : InMux
    port map (
            O => \N__36161\,
            I => \N__35930\
        );

    \I__8988\ : InMux
    port map (
            O => \N__36160\,
            I => \N__35930\
        );

    \I__8987\ : InMux
    port map (
            O => \N__36159\,
            I => \N__35930\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__36154\,
            I => \N__35925\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__36147\,
            I => \N__35925\
        );

    \I__8984\ : InMux
    port map (
            O => \N__36146\,
            I => \N__35922\
        );

    \I__8983\ : InMux
    port map (
            O => \N__36143\,
            I => \N__35917\
        );

    \I__8982\ : InMux
    port map (
            O => \N__36140\,
            I => \N__35917\
        );

    \I__8981\ : Span4Mux_s1_v
    port map (
            O => \N__36137\,
            I => \N__35904\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__36130\,
            I => \N__35904\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__36123\,
            I => \N__35904\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__36120\,
            I => \N__35904\
        );

    \I__8977\ : Span4Mux_h
    port map (
            O => \N__36113\,
            I => \N__35904\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__36102\,
            I => \N__35904\
        );

    \I__8975\ : InMux
    port map (
            O => \N__36101\,
            I => \N__35901\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__35896\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__36091\,
            I => \N__35896\
        );

    \I__8972\ : InMux
    port map (
            O => \N__36088\,
            I => \N__35887\
        );

    \I__8971\ : InMux
    port map (
            O => \N__36087\,
            I => \N__35887\
        );

    \I__8970\ : InMux
    port map (
            O => \N__36086\,
            I => \N__35887\
        );

    \I__8969\ : InMux
    port map (
            O => \N__36085\,
            I => \N__35887\
        );

    \I__8968\ : InMux
    port map (
            O => \N__36084\,
            I => \N__35878\
        );

    \I__8967\ : InMux
    port map (
            O => \N__36083\,
            I => \N__35878\
        );

    \I__8966\ : InMux
    port map (
            O => \N__36082\,
            I => \N__35878\
        );

    \I__8965\ : InMux
    port map (
            O => \N__36081\,
            I => \N__35878\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__36076\,
            I => \N__35875\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__36073\,
            I => \N__35870\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__36064\,
            I => \N__35870\
        );

    \I__8961\ : InMux
    port map (
            O => \N__36063\,
            I => \N__35865\
        );

    \I__8960\ : InMux
    port map (
            O => \N__36062\,
            I => \N__35865\
        );

    \I__8959\ : InMux
    port map (
            O => \N__36061\,
            I => \N__35846\
        );

    \I__8958\ : InMux
    port map (
            O => \N__36060\,
            I => \N__35846\
        );

    \I__8957\ : InMux
    port map (
            O => \N__36059\,
            I => \N__35846\
        );

    \I__8956\ : InMux
    port map (
            O => \N__36058\,
            I => \N__35846\
        );

    \I__8955\ : InMux
    port map (
            O => \N__36057\,
            I => \N__35846\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__36050\,
            I => \N__35839\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__36045\,
            I => \N__35839\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__36042\,
            I => \N__35839\
        );

    \I__8951\ : InMux
    port map (
            O => \N__36041\,
            I => \N__35832\
        );

    \I__8950\ : InMux
    port map (
            O => \N__36040\,
            I => \N__35832\
        );

    \I__8949\ : InMux
    port map (
            O => \N__36039\,
            I => \N__35825\
        );

    \I__8948\ : InMux
    port map (
            O => \N__36038\,
            I => \N__35825\
        );

    \I__8947\ : InMux
    port map (
            O => \N__36037\,
            I => \N__35825\
        );

    \I__8946\ : InMux
    port map (
            O => \N__36036\,
            I => \N__35818\
        );

    \I__8945\ : InMux
    port map (
            O => \N__36035\,
            I => \N__35818\
        );

    \I__8944\ : InMux
    port map (
            O => \N__36034\,
            I => \N__35818\
        );

    \I__8943\ : InMux
    port map (
            O => \N__36033\,
            I => \N__35809\
        );

    \I__8942\ : InMux
    port map (
            O => \N__36032\,
            I => \N__35809\
        );

    \I__8941\ : InMux
    port map (
            O => \N__36031\,
            I => \N__35809\
        );

    \I__8940\ : InMux
    port map (
            O => \N__36030\,
            I => \N__35809\
        );

    \I__8939\ : InMux
    port map (
            O => \N__36027\,
            I => \N__35800\
        );

    \I__8938\ : InMux
    port map (
            O => \N__36026\,
            I => \N__35800\
        );

    \I__8937\ : InMux
    port map (
            O => \N__36025\,
            I => \N__35800\
        );

    \I__8936\ : InMux
    port map (
            O => \N__36024\,
            I => \N__35800\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__36019\,
            I => \N__35797\
        );

    \I__8934\ : InMux
    port map (
            O => \N__36018\,
            I => \N__35792\
        );

    \I__8933\ : InMux
    port map (
            O => \N__36017\,
            I => \N__35792\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__36014\,
            I => \N__35789\
        );

    \I__8931\ : InMux
    port map (
            O => \N__36013\,
            I => \N__35786\
        );

    \I__8930\ : InMux
    port map (
            O => \N__36012\,
            I => \N__35781\
        );

    \I__8929\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35781\
        );

    \I__8928\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35772\
        );

    \I__8927\ : InMux
    port map (
            O => \N__36007\,
            I => \N__35772\
        );

    \I__8926\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35772\
        );

    \I__8925\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35772\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__36000\,
            I => \N__35769\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__35997\,
            I => \N__35765\
        );

    \I__8922\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35762\
        );

    \I__8921\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35755\
        );

    \I__8920\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35755\
        );

    \I__8919\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35755\
        );

    \I__8918\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35744\
        );

    \I__8917\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35744\
        );

    \I__8916\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35744\
        );

    \I__8915\ : InMux
    port map (
            O => \N__35987\,
            I => \N__35744\
        );

    \I__8914\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35744\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__35981\,
            I => \N__35741\
        );

    \I__8912\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35738\
        );

    \I__8911\ : Span4Mux_v
    port map (
            O => \N__35975\,
            I => \N__35735\
        );

    \I__8910\ : Span4Mux_h
    port map (
            O => \N__35970\,
            I => \N__35730\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__35967\,
            I => \N__35730\
        );

    \I__8908\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35727\
        );

    \I__8907\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35722\
        );

    \I__8906\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35722\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__35961\,
            I => \N__35717\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__35956\,
            I => \N__35717\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__35951\,
            I => \N__35706\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__35944\,
            I => \N__35706\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__35939\,
            I => \N__35706\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__35930\,
            I => \N__35706\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__35925\,
            I => \N__35706\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__35922\,
            I => \N__35701\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__35917\,
            I => \N__35701\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__35904\,
            I => \N__35698\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__35901\,
            I => \N__35683\
        );

    \I__8894\ : Span4Mux_h
    port map (
            O => \N__35896\,
            I => \N__35683\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__35887\,
            I => \N__35683\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35683\
        );

    \I__8891\ : Span4Mux_v
    port map (
            O => \N__35875\,
            I => \N__35683\
        );

    \I__8890\ : Span4Mux_h
    port map (
            O => \N__35870\,
            I => \N__35683\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__35865\,
            I => \N__35683\
        );

    \I__8888\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35680\
        );

    \I__8887\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35677\
        );

    \I__8886\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35674\
        );

    \I__8885\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35663\
        );

    \I__8884\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35663\
        );

    \I__8883\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35663\
        );

    \I__8882\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35663\
        );

    \I__8881\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35663\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__35846\,
            I => \N__35660\
        );

    \I__8879\ : Span4Mux_v
    port map (
            O => \N__35839\,
            I => \N__35657\
        );

    \I__8878\ : InMux
    port map (
            O => \N__35838\,
            I => \N__35654\
        );

    \I__8877\ : CascadeMux
    port map (
            O => \N__35837\,
            I => \N__35636\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__35832\,
            I => \N__35633\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__35825\,
            I => \N__35628\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__35818\,
            I => \N__35628\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35625\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35620\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__35797\,
            I => \N__35620\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35615\
        );

    \I__8869\ : Span4Mux_v
    port map (
            O => \N__35789\,
            I => \N__35615\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__35786\,
            I => \N__35606\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__35781\,
            I => \N__35606\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__35772\,
            I => \N__35606\
        );

    \I__8865\ : Span4Mux_v
    port map (
            O => \N__35769\,
            I => \N__35606\
        );

    \I__8864\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35603\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__35765\,
            I => \N__35600\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__35762\,
            I => \N__35595\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35595\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__35744\,
            I => \N__35590\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__35741\,
            I => \N__35590\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35583\
        );

    \I__8857\ : Span4Mux_s0_h
    port map (
            O => \N__35735\,
            I => \N__35583\
        );

    \I__8856\ : Span4Mux_v
    port map (
            O => \N__35730\,
            I => \N__35583\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__35727\,
            I => \N__35574\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__35722\,
            I => \N__35574\
        );

    \I__8853\ : Span4Mux_v
    port map (
            O => \N__35717\,
            I => \N__35574\
        );

    \I__8852\ : Span4Mux_v
    port map (
            O => \N__35706\,
            I => \N__35574\
        );

    \I__8851\ : Span4Mux_v
    port map (
            O => \N__35701\,
            I => \N__35571\
        );

    \I__8850\ : Span4Mux_s1_v
    port map (
            O => \N__35698\,
            I => \N__35566\
        );

    \I__8849\ : Span4Mux_v
    port map (
            O => \N__35683\,
            I => \N__35566\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35559\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__35677\,
            I => \N__35559\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__35674\,
            I => \N__35559\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__35663\,
            I => \N__35556\
        );

    \I__8844\ : Span4Mux_h
    port map (
            O => \N__35660\,
            I => \N__35549\
        );

    \I__8843\ : Span4Mux_h
    port map (
            O => \N__35657\,
            I => \N__35549\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__35654\,
            I => \N__35549\
        );

    \I__8841\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35546\
        );

    \I__8840\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35543\
        );

    \I__8839\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35536\
        );

    \I__8838\ : InMux
    port map (
            O => \N__35650\,
            I => \N__35536\
        );

    \I__8837\ : InMux
    port map (
            O => \N__35649\,
            I => \N__35536\
        );

    \I__8836\ : InMux
    port map (
            O => \N__35648\,
            I => \N__35529\
        );

    \I__8835\ : InMux
    port map (
            O => \N__35647\,
            I => \N__35529\
        );

    \I__8834\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35529\
        );

    \I__8833\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35524\
        );

    \I__8832\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35524\
        );

    \I__8831\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35517\
        );

    \I__8830\ : InMux
    port map (
            O => \N__35642\,
            I => \N__35517\
        );

    \I__8829\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35517\
        );

    \I__8828\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35512\
        );

    \I__8827\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35512\
        );

    \I__8826\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35509\
        );

    \I__8825\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35506\
        );

    \I__8824\ : Span4Mux_h
    port map (
            O => \N__35628\,
            I => \N__35503\
        );

    \I__8823\ : Span4Mux_v
    port map (
            O => \N__35625\,
            I => \N__35494\
        );

    \I__8822\ : Span4Mux_h
    port map (
            O => \N__35620\,
            I => \N__35494\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__35615\,
            I => \N__35494\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__35606\,
            I => \N__35494\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__35603\,
            I => \N__35481\
        );

    \I__8818\ : Span4Mux_s1_v
    port map (
            O => \N__35600\,
            I => \N__35481\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__35595\,
            I => \N__35481\
        );

    \I__8816\ : Span4Mux_v
    port map (
            O => \N__35590\,
            I => \N__35481\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__35583\,
            I => \N__35481\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__35574\,
            I => \N__35481\
        );

    \I__8813\ : Span4Mux_s1_v
    port map (
            O => \N__35571\,
            I => \N__35476\
        );

    \I__8812\ : Span4Mux_h
    port map (
            O => \N__35566\,
            I => \N__35476\
        );

    \I__8811\ : Span12Mux_h
    port map (
            O => \N__35559\,
            I => \N__35469\
        );

    \I__8810\ : Span12Mux_v
    port map (
            O => \N__35556\,
            I => \N__35469\
        );

    \I__8809\ : Sp12to4
    port map (
            O => \N__35549\,
            I => \N__35469\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__35546\,
            I => \c0.n1686\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__35543\,
            I => \c0.n1686\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__35536\,
            I => \c0.n1686\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__35529\,
            I => \c0.n1686\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__35524\,
            I => \c0.n1686\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__35517\,
            I => \c0.n1686\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__35512\,
            I => \c0.n1686\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__35509\,
            I => \c0.n1686\
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__35506\,
            I => \c0.n1686\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__35503\,
            I => \c0.n1686\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__35494\,
            I => \c0.n1686\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__35481\,
            I => \c0.n1686\
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__35476\,
            I => \c0.n1686\
        );

    \I__8795\ : Odrv12
    port map (
            O => \N__35469\,
            I => \c0.n1686\
        );

    \I__8794\ : CascadeMux
    port map (
            O => \N__35440\,
            I => \N__35437\
        );

    \I__8793\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35434\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__35434\,
            I => \N__35431\
        );

    \I__8791\ : Span4Mux_s3_h
    port map (
            O => \N__35431\,
            I => \N__35428\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__35428\,
            I => \N__35425\
        );

    \I__8789\ : Span4Mux_h
    port map (
            O => \N__35425\,
            I => \N__35421\
        );

    \I__8788\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35418\
        );

    \I__8787\ : Span4Mux_h
    port map (
            O => \N__35421\,
            I => \N__35415\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__35418\,
            I => \c0.data_in_frame_19_4\
        );

    \I__8785\ : Odrv4
    port map (
            O => \N__35415\,
            I => \c0.data_in_frame_19_4\
        );

    \I__8784\ : ClkMux
    port map (
            O => \N__35410\,
            I => \N__34984\
        );

    \I__8783\ : ClkMux
    port map (
            O => \N__35409\,
            I => \N__34984\
        );

    \I__8782\ : ClkMux
    port map (
            O => \N__35408\,
            I => \N__34984\
        );

    \I__8781\ : ClkMux
    port map (
            O => \N__35407\,
            I => \N__34984\
        );

    \I__8780\ : ClkMux
    port map (
            O => \N__35406\,
            I => \N__34984\
        );

    \I__8779\ : ClkMux
    port map (
            O => \N__35405\,
            I => \N__34984\
        );

    \I__8778\ : ClkMux
    port map (
            O => \N__35404\,
            I => \N__34984\
        );

    \I__8777\ : ClkMux
    port map (
            O => \N__35403\,
            I => \N__34984\
        );

    \I__8776\ : ClkMux
    port map (
            O => \N__35402\,
            I => \N__34984\
        );

    \I__8775\ : ClkMux
    port map (
            O => \N__35401\,
            I => \N__34984\
        );

    \I__8774\ : ClkMux
    port map (
            O => \N__35400\,
            I => \N__34984\
        );

    \I__8773\ : ClkMux
    port map (
            O => \N__35399\,
            I => \N__34984\
        );

    \I__8772\ : ClkMux
    port map (
            O => \N__35398\,
            I => \N__34984\
        );

    \I__8771\ : ClkMux
    port map (
            O => \N__35397\,
            I => \N__34984\
        );

    \I__8770\ : ClkMux
    port map (
            O => \N__35396\,
            I => \N__34984\
        );

    \I__8769\ : ClkMux
    port map (
            O => \N__35395\,
            I => \N__34984\
        );

    \I__8768\ : ClkMux
    port map (
            O => \N__35394\,
            I => \N__34984\
        );

    \I__8767\ : ClkMux
    port map (
            O => \N__35393\,
            I => \N__34984\
        );

    \I__8766\ : ClkMux
    port map (
            O => \N__35392\,
            I => \N__34984\
        );

    \I__8765\ : ClkMux
    port map (
            O => \N__35391\,
            I => \N__34984\
        );

    \I__8764\ : ClkMux
    port map (
            O => \N__35390\,
            I => \N__34984\
        );

    \I__8763\ : ClkMux
    port map (
            O => \N__35389\,
            I => \N__34984\
        );

    \I__8762\ : ClkMux
    port map (
            O => \N__35388\,
            I => \N__34984\
        );

    \I__8761\ : ClkMux
    port map (
            O => \N__35387\,
            I => \N__34984\
        );

    \I__8760\ : ClkMux
    port map (
            O => \N__35386\,
            I => \N__34984\
        );

    \I__8759\ : ClkMux
    port map (
            O => \N__35385\,
            I => \N__34984\
        );

    \I__8758\ : ClkMux
    port map (
            O => \N__35384\,
            I => \N__34984\
        );

    \I__8757\ : ClkMux
    port map (
            O => \N__35383\,
            I => \N__34984\
        );

    \I__8756\ : ClkMux
    port map (
            O => \N__35382\,
            I => \N__34984\
        );

    \I__8755\ : ClkMux
    port map (
            O => \N__35381\,
            I => \N__34984\
        );

    \I__8754\ : ClkMux
    port map (
            O => \N__35380\,
            I => \N__34984\
        );

    \I__8753\ : ClkMux
    port map (
            O => \N__35379\,
            I => \N__34984\
        );

    \I__8752\ : ClkMux
    port map (
            O => \N__35378\,
            I => \N__34984\
        );

    \I__8751\ : ClkMux
    port map (
            O => \N__35377\,
            I => \N__34984\
        );

    \I__8750\ : ClkMux
    port map (
            O => \N__35376\,
            I => \N__34984\
        );

    \I__8749\ : ClkMux
    port map (
            O => \N__35375\,
            I => \N__34984\
        );

    \I__8748\ : ClkMux
    port map (
            O => \N__35374\,
            I => \N__34984\
        );

    \I__8747\ : ClkMux
    port map (
            O => \N__35373\,
            I => \N__34984\
        );

    \I__8746\ : ClkMux
    port map (
            O => \N__35372\,
            I => \N__34984\
        );

    \I__8745\ : ClkMux
    port map (
            O => \N__35371\,
            I => \N__34984\
        );

    \I__8744\ : ClkMux
    port map (
            O => \N__35370\,
            I => \N__34984\
        );

    \I__8743\ : ClkMux
    port map (
            O => \N__35369\,
            I => \N__34984\
        );

    \I__8742\ : ClkMux
    port map (
            O => \N__35368\,
            I => \N__34984\
        );

    \I__8741\ : ClkMux
    port map (
            O => \N__35367\,
            I => \N__34984\
        );

    \I__8740\ : ClkMux
    port map (
            O => \N__35366\,
            I => \N__34984\
        );

    \I__8739\ : ClkMux
    port map (
            O => \N__35365\,
            I => \N__34984\
        );

    \I__8738\ : ClkMux
    port map (
            O => \N__35364\,
            I => \N__34984\
        );

    \I__8737\ : ClkMux
    port map (
            O => \N__35363\,
            I => \N__34984\
        );

    \I__8736\ : ClkMux
    port map (
            O => \N__35362\,
            I => \N__34984\
        );

    \I__8735\ : ClkMux
    port map (
            O => \N__35361\,
            I => \N__34984\
        );

    \I__8734\ : ClkMux
    port map (
            O => \N__35360\,
            I => \N__34984\
        );

    \I__8733\ : ClkMux
    port map (
            O => \N__35359\,
            I => \N__34984\
        );

    \I__8732\ : ClkMux
    port map (
            O => \N__35358\,
            I => \N__34984\
        );

    \I__8731\ : ClkMux
    port map (
            O => \N__35357\,
            I => \N__34984\
        );

    \I__8730\ : ClkMux
    port map (
            O => \N__35356\,
            I => \N__34984\
        );

    \I__8729\ : ClkMux
    port map (
            O => \N__35355\,
            I => \N__34984\
        );

    \I__8728\ : ClkMux
    port map (
            O => \N__35354\,
            I => \N__34984\
        );

    \I__8727\ : ClkMux
    port map (
            O => \N__35353\,
            I => \N__34984\
        );

    \I__8726\ : ClkMux
    port map (
            O => \N__35352\,
            I => \N__34984\
        );

    \I__8725\ : ClkMux
    port map (
            O => \N__35351\,
            I => \N__34984\
        );

    \I__8724\ : ClkMux
    port map (
            O => \N__35350\,
            I => \N__34984\
        );

    \I__8723\ : ClkMux
    port map (
            O => \N__35349\,
            I => \N__34984\
        );

    \I__8722\ : ClkMux
    port map (
            O => \N__35348\,
            I => \N__34984\
        );

    \I__8721\ : ClkMux
    port map (
            O => \N__35347\,
            I => \N__34984\
        );

    \I__8720\ : ClkMux
    port map (
            O => \N__35346\,
            I => \N__34984\
        );

    \I__8719\ : ClkMux
    port map (
            O => \N__35345\,
            I => \N__34984\
        );

    \I__8718\ : ClkMux
    port map (
            O => \N__35344\,
            I => \N__34984\
        );

    \I__8717\ : ClkMux
    port map (
            O => \N__35343\,
            I => \N__34984\
        );

    \I__8716\ : ClkMux
    port map (
            O => \N__35342\,
            I => \N__34984\
        );

    \I__8715\ : ClkMux
    port map (
            O => \N__35341\,
            I => \N__34984\
        );

    \I__8714\ : ClkMux
    port map (
            O => \N__35340\,
            I => \N__34984\
        );

    \I__8713\ : ClkMux
    port map (
            O => \N__35339\,
            I => \N__34984\
        );

    \I__8712\ : ClkMux
    port map (
            O => \N__35338\,
            I => \N__34984\
        );

    \I__8711\ : ClkMux
    port map (
            O => \N__35337\,
            I => \N__34984\
        );

    \I__8710\ : ClkMux
    port map (
            O => \N__35336\,
            I => \N__34984\
        );

    \I__8709\ : ClkMux
    port map (
            O => \N__35335\,
            I => \N__34984\
        );

    \I__8708\ : ClkMux
    port map (
            O => \N__35334\,
            I => \N__34984\
        );

    \I__8707\ : ClkMux
    port map (
            O => \N__35333\,
            I => \N__34984\
        );

    \I__8706\ : ClkMux
    port map (
            O => \N__35332\,
            I => \N__34984\
        );

    \I__8705\ : ClkMux
    port map (
            O => \N__35331\,
            I => \N__34984\
        );

    \I__8704\ : ClkMux
    port map (
            O => \N__35330\,
            I => \N__34984\
        );

    \I__8703\ : ClkMux
    port map (
            O => \N__35329\,
            I => \N__34984\
        );

    \I__8702\ : ClkMux
    port map (
            O => \N__35328\,
            I => \N__34984\
        );

    \I__8701\ : ClkMux
    port map (
            O => \N__35327\,
            I => \N__34984\
        );

    \I__8700\ : ClkMux
    port map (
            O => \N__35326\,
            I => \N__34984\
        );

    \I__8699\ : ClkMux
    port map (
            O => \N__35325\,
            I => \N__34984\
        );

    \I__8698\ : ClkMux
    port map (
            O => \N__35324\,
            I => \N__34984\
        );

    \I__8697\ : ClkMux
    port map (
            O => \N__35323\,
            I => \N__34984\
        );

    \I__8696\ : ClkMux
    port map (
            O => \N__35322\,
            I => \N__34984\
        );

    \I__8695\ : ClkMux
    port map (
            O => \N__35321\,
            I => \N__34984\
        );

    \I__8694\ : ClkMux
    port map (
            O => \N__35320\,
            I => \N__34984\
        );

    \I__8693\ : ClkMux
    port map (
            O => \N__35319\,
            I => \N__34984\
        );

    \I__8692\ : ClkMux
    port map (
            O => \N__35318\,
            I => \N__34984\
        );

    \I__8691\ : ClkMux
    port map (
            O => \N__35317\,
            I => \N__34984\
        );

    \I__8690\ : ClkMux
    port map (
            O => \N__35316\,
            I => \N__34984\
        );

    \I__8689\ : ClkMux
    port map (
            O => \N__35315\,
            I => \N__34984\
        );

    \I__8688\ : ClkMux
    port map (
            O => \N__35314\,
            I => \N__34984\
        );

    \I__8687\ : ClkMux
    port map (
            O => \N__35313\,
            I => \N__34984\
        );

    \I__8686\ : ClkMux
    port map (
            O => \N__35312\,
            I => \N__34984\
        );

    \I__8685\ : ClkMux
    port map (
            O => \N__35311\,
            I => \N__34984\
        );

    \I__8684\ : ClkMux
    port map (
            O => \N__35310\,
            I => \N__34984\
        );

    \I__8683\ : ClkMux
    port map (
            O => \N__35309\,
            I => \N__34984\
        );

    \I__8682\ : ClkMux
    port map (
            O => \N__35308\,
            I => \N__34984\
        );

    \I__8681\ : ClkMux
    port map (
            O => \N__35307\,
            I => \N__34984\
        );

    \I__8680\ : ClkMux
    port map (
            O => \N__35306\,
            I => \N__34984\
        );

    \I__8679\ : ClkMux
    port map (
            O => \N__35305\,
            I => \N__34984\
        );

    \I__8678\ : ClkMux
    port map (
            O => \N__35304\,
            I => \N__34984\
        );

    \I__8677\ : ClkMux
    port map (
            O => \N__35303\,
            I => \N__34984\
        );

    \I__8676\ : ClkMux
    port map (
            O => \N__35302\,
            I => \N__34984\
        );

    \I__8675\ : ClkMux
    port map (
            O => \N__35301\,
            I => \N__34984\
        );

    \I__8674\ : ClkMux
    port map (
            O => \N__35300\,
            I => \N__34984\
        );

    \I__8673\ : ClkMux
    port map (
            O => \N__35299\,
            I => \N__34984\
        );

    \I__8672\ : ClkMux
    port map (
            O => \N__35298\,
            I => \N__34984\
        );

    \I__8671\ : ClkMux
    port map (
            O => \N__35297\,
            I => \N__34984\
        );

    \I__8670\ : ClkMux
    port map (
            O => \N__35296\,
            I => \N__34984\
        );

    \I__8669\ : ClkMux
    port map (
            O => \N__35295\,
            I => \N__34984\
        );

    \I__8668\ : ClkMux
    port map (
            O => \N__35294\,
            I => \N__34984\
        );

    \I__8667\ : ClkMux
    port map (
            O => \N__35293\,
            I => \N__34984\
        );

    \I__8666\ : ClkMux
    port map (
            O => \N__35292\,
            I => \N__34984\
        );

    \I__8665\ : ClkMux
    port map (
            O => \N__35291\,
            I => \N__34984\
        );

    \I__8664\ : ClkMux
    port map (
            O => \N__35290\,
            I => \N__34984\
        );

    \I__8663\ : ClkMux
    port map (
            O => \N__35289\,
            I => \N__34984\
        );

    \I__8662\ : ClkMux
    port map (
            O => \N__35288\,
            I => \N__34984\
        );

    \I__8661\ : ClkMux
    port map (
            O => \N__35287\,
            I => \N__34984\
        );

    \I__8660\ : ClkMux
    port map (
            O => \N__35286\,
            I => \N__34984\
        );

    \I__8659\ : ClkMux
    port map (
            O => \N__35285\,
            I => \N__34984\
        );

    \I__8658\ : ClkMux
    port map (
            O => \N__35284\,
            I => \N__34984\
        );

    \I__8657\ : ClkMux
    port map (
            O => \N__35283\,
            I => \N__34984\
        );

    \I__8656\ : ClkMux
    port map (
            O => \N__35282\,
            I => \N__34984\
        );

    \I__8655\ : ClkMux
    port map (
            O => \N__35281\,
            I => \N__34984\
        );

    \I__8654\ : ClkMux
    port map (
            O => \N__35280\,
            I => \N__34984\
        );

    \I__8653\ : ClkMux
    port map (
            O => \N__35279\,
            I => \N__34984\
        );

    \I__8652\ : ClkMux
    port map (
            O => \N__35278\,
            I => \N__34984\
        );

    \I__8651\ : ClkMux
    port map (
            O => \N__35277\,
            I => \N__34984\
        );

    \I__8650\ : ClkMux
    port map (
            O => \N__35276\,
            I => \N__34984\
        );

    \I__8649\ : ClkMux
    port map (
            O => \N__35275\,
            I => \N__34984\
        );

    \I__8648\ : ClkMux
    port map (
            O => \N__35274\,
            I => \N__34984\
        );

    \I__8647\ : ClkMux
    port map (
            O => \N__35273\,
            I => \N__34984\
        );

    \I__8646\ : ClkMux
    port map (
            O => \N__35272\,
            I => \N__34984\
        );

    \I__8645\ : ClkMux
    port map (
            O => \N__35271\,
            I => \N__34984\
        );

    \I__8644\ : ClkMux
    port map (
            O => \N__35270\,
            I => \N__34984\
        );

    \I__8643\ : ClkMux
    port map (
            O => \N__35269\,
            I => \N__34984\
        );

    \I__8642\ : GlobalMux
    port map (
            O => \N__34984\,
            I => \N__34981\
        );

    \I__8641\ : gio2CtrlBuf
    port map (
            O => \N__34981\,
            I => \CLK_c\
        );

    \I__8640\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34975\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__34975\,
            I => n13
        );

    \I__8638\ : InMux
    port map (
            O => \N__34972\,
            I => n4449
        );

    \I__8637\ : InMux
    port map (
            O => \N__34969\,
            I => \N__34966\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__34966\,
            I => n12
        );

    \I__8635\ : InMux
    port map (
            O => \N__34963\,
            I => n4450
        );

    \I__8634\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34957\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__34957\,
            I => n11
        );

    \I__8632\ : InMux
    port map (
            O => \N__34954\,
            I => n4451
        );

    \I__8631\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34948\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__34948\,
            I => n10
        );

    \I__8629\ : InMux
    port map (
            O => \N__34945\,
            I => \bfn_15_27_0_\
        );

    \I__8628\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34939\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__34939\,
            I => n9
        );

    \I__8626\ : InMux
    port map (
            O => \N__34936\,
            I => n4453
        );

    \I__8625\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34930\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__34930\,
            I => n8_adj_1989
        );

    \I__8623\ : InMux
    port map (
            O => \N__34927\,
            I => n4454
        );

    \I__8622\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34921\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__34921\,
            I => n7
        );

    \I__8620\ : InMux
    port map (
            O => \N__34918\,
            I => n4455
        );

    \I__8619\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34912\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__34912\,
            I => n6
        );

    \I__8617\ : InMux
    port map (
            O => \N__34909\,
            I => n4456
        );

    \I__8616\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34903\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__34903\,
            I => n21
        );

    \I__8614\ : InMux
    port map (
            O => \N__34900\,
            I => n4441
        );

    \I__8613\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34894\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__34894\,
            I => n20
        );

    \I__8611\ : InMux
    port map (
            O => \N__34891\,
            I => n4442
        );

    \I__8610\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34885\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__34885\,
            I => n19
        );

    \I__8608\ : InMux
    port map (
            O => \N__34882\,
            I => n4443
        );

    \I__8607\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34876\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__34876\,
            I => n18
        );

    \I__8605\ : InMux
    port map (
            O => \N__34873\,
            I => \bfn_15_26_0_\
        );

    \I__8604\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34867\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__34867\,
            I => n17
        );

    \I__8602\ : InMux
    port map (
            O => \N__34864\,
            I => n4445
        );

    \I__8601\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34858\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__34858\,
            I => n16
        );

    \I__8599\ : InMux
    port map (
            O => \N__34855\,
            I => n4446
        );

    \I__8598\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34849\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__34849\,
            I => n15
        );

    \I__8596\ : InMux
    port map (
            O => \N__34846\,
            I => n4447
        );

    \I__8595\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34840\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__34840\,
            I => n14
        );

    \I__8593\ : InMux
    port map (
            O => \N__34837\,
            I => n4448
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__34834\,
            I => \c0.n5887_cascade_\
        );

    \I__8591\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34822\
        );

    \I__8590\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34822\
        );

    \I__8589\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34817\
        );

    \I__8588\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34814\
        );

    \I__8587\ : CascadeMux
    port map (
            O => \N__34827\,
            I => \N__34808\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__34822\,
            I => \N__34801\
        );

    \I__8585\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34797\
        );

    \I__8584\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34794\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__34817\,
            I => \N__34789\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__34814\,
            I => \N__34789\
        );

    \I__8581\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34786\
        );

    \I__8580\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34783\
        );

    \I__8579\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34778\
        );

    \I__8578\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34778\
        );

    \I__8577\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34775\
        );

    \I__8576\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34772\
        );

    \I__8575\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34769\
        );

    \I__8574\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34766\
        );

    \I__8573\ : Span4Mux_v
    port map (
            O => \N__34801\,
            I => \N__34763\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__34800\,
            I => \N__34758\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__34797\,
            I => \N__34755\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__34794\,
            I => \N__34748\
        );

    \I__8569\ : Span4Mux_h
    port map (
            O => \N__34789\,
            I => \N__34748\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__34786\,
            I => \N__34748\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__34783\,
            I => \N__34744\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__34778\,
            I => \N__34735\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__34775\,
            I => \N__34735\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__34772\,
            I => \N__34735\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__34769\,
            I => \N__34735\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34730\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__34763\,
            I => \N__34730\
        );

    \I__8560\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34727\
        );

    \I__8559\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34722\
        );

    \I__8558\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34722\
        );

    \I__8557\ : Span4Mux_s3_h
    port map (
            O => \N__34755\,
            I => \N__34717\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__34748\,
            I => \N__34717\
        );

    \I__8555\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34714\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__34744\,
            I => \N__34707\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__34735\,
            I => \N__34707\
        );

    \I__8552\ : Span4Mux_h
    port map (
            O => \N__34730\,
            I => \N__34707\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__34727\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__34722\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__34717\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__34714\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__34707\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__8546\ : InMux
    port map (
            O => \N__34696\,
            I => \N__34693\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__34693\,
            I => \N__34690\
        );

    \I__8544\ : Span12Mux_h
    port map (
            O => \N__34690\,
            I => \N__34687\
        );

    \I__8543\ : Odrv12
    port map (
            O => \N__34687\,
            I => \c0.n5890\
        );

    \I__8542\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34681\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__34681\,
            I => \N__34677\
        );

    \I__8540\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34674\
        );

    \I__8539\ : Span4Mux_h
    port map (
            O => \N__34677\,
            I => \N__34671\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34668\
        );

    \I__8537\ : Span4Mux_h
    port map (
            O => \N__34671\,
            I => \N__34664\
        );

    \I__8536\ : Span4Mux_h
    port map (
            O => \N__34668\,
            I => \N__34661\
        );

    \I__8535\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34658\
        );

    \I__8534\ : Odrv4
    port map (
            O => \N__34664\,
            I => \c0.n5219\
        );

    \I__8533\ : Odrv4
    port map (
            O => \N__34661\,
            I => \c0.n5219\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__34658\,
            I => \c0.n5219\
        );

    \I__8531\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34648\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__34648\,
            I => \N__34644\
        );

    \I__8529\ : InMux
    port map (
            O => \N__34647\,
            I => \N__34641\
        );

    \I__8528\ : Odrv4
    port map (
            O => \N__34644\,
            I => \c0.n5138\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__34641\,
            I => \c0.n5138\
        );

    \I__8526\ : CascadeMux
    port map (
            O => \N__34636\,
            I => \N__34633\
        );

    \I__8525\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34627\
        );

    \I__8523\ : Span4Mux_h
    port map (
            O => \N__34627\,
            I => \N__34624\
        );

    \I__8522\ : Span4Mux_h
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__34621\,
            I => \c0.n1896\
        );

    \I__8520\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34614\
        );

    \I__8519\ : CascadeMux
    port map (
            O => \N__34617\,
            I => \N__34610\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__34614\,
            I => \N__34607\
        );

    \I__8517\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34604\
        );

    \I__8516\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34601\
        );

    \I__8515\ : Span4Mux_h
    port map (
            O => \N__34607\,
            I => \N__34598\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__34604\,
            I => data_in_8_4
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__34601\,
            I => data_in_8_4
        );

    \I__8512\ : Odrv4
    port map (
            O => \N__34598\,
            I => data_in_8_4
        );

    \I__8511\ : CascadeMux
    port map (
            O => \N__34591\,
            I => \N__34588\
        );

    \I__8510\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34584\
        );

    \I__8509\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34581\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__34584\,
            I => \N__34576\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__34581\,
            I => \N__34576\
        );

    \I__8506\ : Span4Mux_v
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__8505\ : Span4Mux_h
    port map (
            O => \N__34573\,
            I => \N__34569\
        );

    \I__8504\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34566\
        );

    \I__8503\ : Odrv4
    port map (
            O => \N__34569\,
            I => data_in_7_4
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__34566\,
            I => data_in_7_4
        );

    \I__8501\ : CascadeMux
    port map (
            O => \N__34561\,
            I => \N__34554\
        );

    \I__8500\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34514\
        );

    \I__8499\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34514\
        );

    \I__8498\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34514\
        );

    \I__8497\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34514\
        );

    \I__8496\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34509\
        );

    \I__8495\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34509\
        );

    \I__8494\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34506\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__34551\,
            I => \N__34502\
        );

    \I__8492\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34487\
        );

    \I__8491\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34482\
        );

    \I__8490\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34482\
        );

    \I__8489\ : CascadeMux
    port map (
            O => \N__34547\,
            I => \N__34479\
        );

    \I__8488\ : CascadeMux
    port map (
            O => \N__34546\,
            I => \N__34475\
        );

    \I__8487\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34468\
        );

    \I__8486\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34468\
        );

    \I__8485\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34461\
        );

    \I__8484\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34455\
        );

    \I__8483\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34452\
        );

    \I__8482\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34441\
        );

    \I__8481\ : InMux
    port map (
            O => \N__34539\,
            I => \N__34441\
        );

    \I__8480\ : InMux
    port map (
            O => \N__34538\,
            I => \N__34438\
        );

    \I__8479\ : CascadeMux
    port map (
            O => \N__34537\,
            I => \N__34435\
        );

    \I__8478\ : CascadeMux
    port map (
            O => \N__34536\,
            I => \N__34432\
        );

    \I__8477\ : CascadeMux
    port map (
            O => \N__34535\,
            I => \N__34418\
        );

    \I__8476\ : CascadeMux
    port map (
            O => \N__34534\,
            I => \N__34409\
        );

    \I__8475\ : InMux
    port map (
            O => \N__34533\,
            I => \N__34403\
        );

    \I__8474\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34398\
        );

    \I__8473\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34398\
        );

    \I__8472\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34391\
        );

    \I__8471\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34391\
        );

    \I__8470\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34391\
        );

    \I__8469\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34386\
        );

    \I__8468\ : InMux
    port map (
            O => \N__34526\,
            I => \N__34386\
        );

    \I__8467\ : InMux
    port map (
            O => \N__34525\,
            I => \N__34383\
        );

    \I__8466\ : InMux
    port map (
            O => \N__34524\,
            I => \N__34380\
        );

    \I__8465\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34375\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__34514\,
            I => \N__34368\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__34509\,
            I => \N__34368\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__34506\,
            I => \N__34368\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__34505\,
            I => \N__34364\
        );

    \I__8460\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34354\
        );

    \I__8459\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34354\
        );

    \I__8458\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34354\
        );

    \I__8457\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34349\
        );

    \I__8456\ : InMux
    port map (
            O => \N__34498\,
            I => \N__34349\
        );

    \I__8455\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34342\
        );

    \I__8454\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34342\
        );

    \I__8453\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34342\
        );

    \I__8452\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34337\
        );

    \I__8451\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34337\
        );

    \I__8450\ : InMux
    port map (
            O => \N__34492\,
            I => \N__34334\
        );

    \I__8449\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34329\
        );

    \I__8448\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34329\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__34487\,
            I => \N__34324\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34324\
        );

    \I__8445\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34321\
        );

    \I__8444\ : InMux
    port map (
            O => \N__34478\,
            I => \N__34310\
        );

    \I__8443\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34310\
        );

    \I__8442\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34310\
        );

    \I__8441\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34310\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__34468\,
            I => \N__34307\
        );

    \I__8439\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34302\
        );

    \I__8438\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34302\
        );

    \I__8437\ : InMux
    port map (
            O => \N__34465\,
            I => \N__34297\
        );

    \I__8436\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34297\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__34461\,
            I => \N__34291\
        );

    \I__8434\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34288\
        );

    \I__8433\ : InMux
    port map (
            O => \N__34459\,
            I => \N__34273\
        );

    \I__8432\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34273\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__34455\,
            I => \N__34268\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__34452\,
            I => \N__34268\
        );

    \I__8429\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34263\
        );

    \I__8428\ : InMux
    port map (
            O => \N__34450\,
            I => \N__34263\
        );

    \I__8427\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34260\
        );

    \I__8426\ : InMux
    port map (
            O => \N__34448\,
            I => \N__34257\
        );

    \I__8425\ : InMux
    port map (
            O => \N__34447\,
            I => \N__34252\
        );

    \I__8424\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34252\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34247\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__34438\,
            I => \N__34247\
        );

    \I__8421\ : InMux
    port map (
            O => \N__34435\,
            I => \N__34232\
        );

    \I__8420\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34232\
        );

    \I__8419\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34232\
        );

    \I__8418\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34232\
        );

    \I__8417\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34232\
        );

    \I__8416\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34232\
        );

    \I__8415\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34232\
        );

    \I__8414\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34221\
        );

    \I__8413\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34221\
        );

    \I__8412\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34221\
        );

    \I__8411\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34221\
        );

    \I__8410\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34221\
        );

    \I__8409\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34212\
        );

    \I__8408\ : InMux
    port map (
            O => \N__34418\,
            I => \N__34203\
        );

    \I__8407\ : InMux
    port map (
            O => \N__34417\,
            I => \N__34203\
        );

    \I__8406\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34203\
        );

    \I__8405\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34203\
        );

    \I__8404\ : InMux
    port map (
            O => \N__34414\,
            I => \N__34196\
        );

    \I__8403\ : InMux
    port map (
            O => \N__34413\,
            I => \N__34196\
        );

    \I__8402\ : InMux
    port map (
            O => \N__34412\,
            I => \N__34196\
        );

    \I__8401\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34189\
        );

    \I__8400\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34189\
        );

    \I__8399\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34189\
        );

    \I__8398\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34186\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34181\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__34398\,
            I => \N__34181\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34172\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__34386\,
            I => \N__34172\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__34383\,
            I => \N__34172\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34172\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__34379\,
            I => \N__34169\
        );

    \I__8390\ : InMux
    port map (
            O => \N__34378\,
            I => \N__34163\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__34375\,
            I => \N__34158\
        );

    \I__8388\ : Span4Mux_v
    port map (
            O => \N__34368\,
            I => \N__34158\
        );

    \I__8387\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34153\
        );

    \I__8386\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34153\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__34363\,
            I => \N__34148\
        );

    \I__8384\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34142\
        );

    \I__8383\ : InMux
    port map (
            O => \N__34361\,
            I => \N__34142\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__34354\,
            I => \N__34135\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34132\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34127\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__34337\,
            I => \N__34127\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34118\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__34329\,
            I => \N__34118\
        );

    \I__8376\ : Span4Mux_h
    port map (
            O => \N__34324\,
            I => \N__34118\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__34321\,
            I => \N__34118\
        );

    \I__8374\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34115\
        );

    \I__8373\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34112\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__34310\,
            I => \N__34103\
        );

    \I__8371\ : Span4Mux_v
    port map (
            O => \N__34307\,
            I => \N__34103\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__34302\,
            I => \N__34103\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__34297\,
            I => \N__34103\
        );

    \I__8368\ : CascadeMux
    port map (
            O => \N__34296\,
            I => \N__34100\
        );

    \I__8367\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34095\
        );

    \I__8366\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34095\
        );

    \I__8365\ : Span4Mux_h
    port map (
            O => \N__34291\,
            I => \N__34090\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34090\
        );

    \I__8363\ : InMux
    port map (
            O => \N__34287\,
            I => \N__34083\
        );

    \I__8362\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34083\
        );

    \I__8361\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34083\
        );

    \I__8360\ : CascadeMux
    port map (
            O => \N__34284\,
            I => \N__34078\
        );

    \I__8359\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34068\
        );

    \I__8358\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34068\
        );

    \I__8357\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34061\
        );

    \I__8356\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34061\
        );

    \I__8355\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34061\
        );

    \I__8354\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34058\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__34273\,
            I => \N__34051\
        );

    \I__8352\ : Span4Mux_v
    port map (
            O => \N__34268\,
            I => \N__34051\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__34263\,
            I => \N__34051\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__34260\,
            I => \N__34038\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__34257\,
            I => \N__34038\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__34252\,
            I => \N__34038\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__34247\,
            I => \N__34038\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__34232\,
            I => \N__34038\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__34221\,
            I => \N__34038\
        );

    \I__8344\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34032\
        );

    \I__8343\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34026\
        );

    \I__8342\ : InMux
    port map (
            O => \N__34218\,
            I => \N__34023\
        );

    \I__8341\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34016\
        );

    \I__8340\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34016\
        );

    \I__8339\ : InMux
    port map (
            O => \N__34215\,
            I => \N__34016\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__34212\,
            I => \N__34000\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34000\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__34196\,
            I => \N__34000\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34000\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__34186\,
            I => \N__33993\
        );

    \I__8333\ : Span4Mux_h
    port map (
            O => \N__34181\,
            I => \N__33993\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__34172\,
            I => \N__33993\
        );

    \I__8331\ : InMux
    port map (
            O => \N__34169\,
            I => \N__33988\
        );

    \I__8330\ : InMux
    port map (
            O => \N__34168\,
            I => \N__33988\
        );

    \I__8329\ : InMux
    port map (
            O => \N__34167\,
            I => \N__33983\
        );

    \I__8328\ : InMux
    port map (
            O => \N__34166\,
            I => \N__33983\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__34163\,
            I => \N__33976\
        );

    \I__8326\ : Span4Mux_h
    port map (
            O => \N__34158\,
            I => \N__33976\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__34153\,
            I => \N__33976\
        );

    \I__8324\ : InMux
    port map (
            O => \N__34152\,
            I => \N__33973\
        );

    \I__8323\ : InMux
    port map (
            O => \N__34151\,
            I => \N__33970\
        );

    \I__8322\ : InMux
    port map (
            O => \N__34148\,
            I => \N__33967\
        );

    \I__8321\ : InMux
    port map (
            O => \N__34147\,
            I => \N__33964\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__34142\,
            I => \N__33961\
        );

    \I__8319\ : InMux
    port map (
            O => \N__34141\,
            I => \N__33954\
        );

    \I__8318\ : InMux
    port map (
            O => \N__34140\,
            I => \N__33954\
        );

    \I__8317\ : InMux
    port map (
            O => \N__34139\,
            I => \N__33954\
        );

    \I__8316\ : InMux
    port map (
            O => \N__34138\,
            I => \N__33951\
        );

    \I__8315\ : Span4Mux_v
    port map (
            O => \N__34135\,
            I => \N__33948\
        );

    \I__8314\ : IoSpan4Mux
    port map (
            O => \N__34132\,
            I => \N__33941\
        );

    \I__8313\ : Span4Mux_v
    port map (
            O => \N__34127\,
            I => \N__33941\
        );

    \I__8312\ : Span4Mux_v
    port map (
            O => \N__34118\,
            I => \N__33941\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__34115\,
            I => \N__33934\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__34112\,
            I => \N__33934\
        );

    \I__8309\ : Span4Mux_v
    port map (
            O => \N__34103\,
            I => \N__33934\
        );

    \I__8308\ : InMux
    port map (
            O => \N__34100\,
            I => \N__33931\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__34095\,
            I => \N__33926\
        );

    \I__8306\ : Span4Mux_v
    port map (
            O => \N__34090\,
            I => \N__33926\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__33923\
        );

    \I__8304\ : InMux
    port map (
            O => \N__34082\,
            I => \N__33907\
        );

    \I__8303\ : InMux
    port map (
            O => \N__34081\,
            I => \N__33907\
        );

    \I__8302\ : InMux
    port map (
            O => \N__34078\,
            I => \N__33907\
        );

    \I__8301\ : InMux
    port map (
            O => \N__34077\,
            I => \N__33907\
        );

    \I__8300\ : InMux
    port map (
            O => \N__34076\,
            I => \N__33907\
        );

    \I__8299\ : InMux
    port map (
            O => \N__34075\,
            I => \N__33904\
        );

    \I__8298\ : InMux
    port map (
            O => \N__34074\,
            I => \N__33901\
        );

    \I__8297\ : InMux
    port map (
            O => \N__34073\,
            I => \N__33898\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__34068\,
            I => \N__33895\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__34061\,
            I => \N__33886\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__34058\,
            I => \N__33886\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__34051\,
            I => \N__33886\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__34038\,
            I => \N__33886\
        );

    \I__8291\ : InMux
    port map (
            O => \N__34037\,
            I => \N__33865\
        );

    \I__8290\ : InMux
    port map (
            O => \N__34036\,
            I => \N__33865\
        );

    \I__8289\ : InMux
    port map (
            O => \N__34035\,
            I => \N__33865\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__34032\,
            I => \N__33862\
        );

    \I__8287\ : InMux
    port map (
            O => \N__34031\,
            I => \N__33855\
        );

    \I__8286\ : InMux
    port map (
            O => \N__34030\,
            I => \N__33855\
        );

    \I__8285\ : InMux
    port map (
            O => \N__34029\,
            I => \N__33855\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__34026\,
            I => \N__33852\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__33847\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__34016\,
            I => \N__33847\
        );

    \I__8281\ : InMux
    port map (
            O => \N__34015\,
            I => \N__33842\
        );

    \I__8280\ : InMux
    port map (
            O => \N__34014\,
            I => \N__33842\
        );

    \I__8279\ : InMux
    port map (
            O => \N__34013\,
            I => \N__33837\
        );

    \I__8278\ : InMux
    port map (
            O => \N__34012\,
            I => \N__33837\
        );

    \I__8277\ : InMux
    port map (
            O => \N__34011\,
            I => \N__33830\
        );

    \I__8276\ : InMux
    port map (
            O => \N__34010\,
            I => \N__33830\
        );

    \I__8275\ : InMux
    port map (
            O => \N__34009\,
            I => \N__33830\
        );

    \I__8274\ : Span4Mux_v
    port map (
            O => \N__34000\,
            I => \N__33827\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__33993\,
            I => \N__33824\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33817\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__33983\,
            I => \N__33817\
        );

    \I__8270\ : Span4Mux_v
    port map (
            O => \N__33976\,
            I => \N__33817\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33812\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__33970\,
            I => \N__33812\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33805\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__33964\,
            I => \N__33805\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__33961\,
            I => \N__33805\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__33954\,
            I => \N__33794\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__33951\,
            I => \N__33794\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__33948\,
            I => \N__33794\
        );

    \I__8261\ : Span4Mux_s0_v
    port map (
            O => \N__33941\,
            I => \N__33794\
        );

    \I__8260\ : Span4Mux_v
    port map (
            O => \N__33934\,
            I => \N__33794\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__33931\,
            I => \N__33787\
        );

    \I__8258\ : Span4Mux_h
    port map (
            O => \N__33926\,
            I => \N__33787\
        );

    \I__8257\ : Span4Mux_v
    port map (
            O => \N__33923\,
            I => \N__33787\
        );

    \I__8256\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33784\
        );

    \I__8255\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33775\
        );

    \I__8254\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33775\
        );

    \I__8253\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33775\
        );

    \I__8252\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33775\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__33907\,
            I => \N__33764\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33764\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__33901\,
            I => \N__33764\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33764\
        );

    \I__8247\ : Sp12to4
    port map (
            O => \N__33895\,
            I => \N__33764\
        );

    \I__8246\ : Span4Mux_v
    port map (
            O => \N__33886\,
            I => \N__33761\
        );

    \I__8245\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33758\
        );

    \I__8244\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33753\
        );

    \I__8243\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33753\
        );

    \I__8242\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33746\
        );

    \I__8241\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33746\
        );

    \I__8240\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33746\
        );

    \I__8239\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33739\
        );

    \I__8238\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33739\
        );

    \I__8237\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33739\
        );

    \I__8236\ : InMux
    port map (
            O => \N__33876\,
            I => \N__33734\
        );

    \I__8235\ : InMux
    port map (
            O => \N__33875\,
            I => \N__33734\
        );

    \I__8234\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33727\
        );

    \I__8233\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33727\
        );

    \I__8232\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33727\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__33865\,
            I => \N__33724\
        );

    \I__8230\ : Span4Mux_h
    port map (
            O => \N__33862\,
            I => \N__33721\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__33855\,
            I => \N__33714\
        );

    \I__8228\ : Span4Mux_v
    port map (
            O => \N__33852\,
            I => \N__33714\
        );

    \I__8227\ : Span4Mux_v
    port map (
            O => \N__33847\,
            I => \N__33714\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__33842\,
            I => \N__33701\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33701\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33701\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__33827\,
            I => \N__33701\
        );

    \I__8222\ : Span4Mux_h
    port map (
            O => \N__33824\,
            I => \N__33701\
        );

    \I__8221\ : Span4Mux_v
    port map (
            O => \N__33817\,
            I => \N__33701\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__33812\,
            I => \N__33692\
        );

    \I__8219\ : Span4Mux_v
    port map (
            O => \N__33805\,
            I => \N__33692\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__33794\,
            I => \N__33692\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__33787\,
            I => \N__33692\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__33784\,
            I => \N__33683\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__33775\,
            I => \N__33683\
        );

    \I__8214\ : Span12Mux_v
    port map (
            O => \N__33764\,
            I => \N__33683\
        );

    \I__8213\ : Sp12to4
    port map (
            O => \N__33761\,
            I => \N__33683\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__33758\,
            I => rx_data_ready
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__33753\,
            I => rx_data_ready
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__33746\,
            I => rx_data_ready
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__33739\,
            I => rx_data_ready
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__33734\,
            I => rx_data_ready
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__33727\,
            I => rx_data_ready
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__33724\,
            I => rx_data_ready
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__33721\,
            I => rx_data_ready
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__33714\,
            I => rx_data_ready
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__33701\,
            I => rx_data_ready
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__33692\,
            I => rx_data_ready
        );

    \I__8201\ : Odrv12
    port map (
            O => \N__33683\,
            I => rx_data_ready
        );

    \I__8200\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33655\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__33655\,
            I => \N__33652\
        );

    \I__8198\ : Span4Mux_h
    port map (
            O => \N__33652\,
            I => \N__33647\
        );

    \I__8197\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33644\
        );

    \I__8196\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33641\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__33647\,
            I => data_in_17_2
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__33644\,
            I => data_in_17_2
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__33641\,
            I => data_in_17_2
        );

    \I__8192\ : CascadeMux
    port map (
            O => \N__33634\,
            I => \N__33631\
        );

    \I__8191\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33627\
        );

    \I__8190\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33624\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33619\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__33624\,
            I => \N__33619\
        );

    \I__8187\ : Span4Mux_v
    port map (
            O => \N__33619\,
            I => \N__33616\
        );

    \I__8186\ : Span4Mux_h
    port map (
            O => \N__33616\,
            I => \N__33612\
        );

    \I__8185\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33609\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__33612\,
            I => data_in_16_2
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__33609\,
            I => data_in_16_2
        );

    \I__8182\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33601\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__33601\,
            I => n26
        );

    \I__8180\ : InMux
    port map (
            O => \N__33598\,
            I => \bfn_15_25_0_\
        );

    \I__8179\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33592\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__33592\,
            I => n25
        );

    \I__8177\ : InMux
    port map (
            O => \N__33589\,
            I => n4437
        );

    \I__8176\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33583\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__33583\,
            I => n24
        );

    \I__8174\ : InMux
    port map (
            O => \N__33580\,
            I => n4438
        );

    \I__8173\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__33574\,
            I => n23
        );

    \I__8171\ : InMux
    port map (
            O => \N__33571\,
            I => n4439
        );

    \I__8170\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33565\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__33565\,
            I => n22
        );

    \I__8168\ : InMux
    port map (
            O => \N__33562\,
            I => n4440
        );

    \I__8167\ : CascadeMux
    port map (
            O => \N__33559\,
            I => \N__33555\
        );

    \I__8166\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33552\
        );

    \I__8165\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33548\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__33552\,
            I => \N__33545\
        );

    \I__8163\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33542\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__33548\,
            I => data_in_9_2
        );

    \I__8161\ : Odrv12
    port map (
            O => \N__33545\,
            I => data_in_9_2
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__33542\,
            I => data_in_9_2
        );

    \I__8159\ : CascadeMux
    port map (
            O => \N__33535\,
            I => \N__33532\
        );

    \I__8158\ : InMux
    port map (
            O => \N__33532\,
            I => \N__33528\
        );

    \I__8157\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33525\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33522\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__33525\,
            I => \N__33519\
        );

    \I__8154\ : Span4Mux_h
    port map (
            O => \N__33522\,
            I => \N__33513\
        );

    \I__8153\ : Span4Mux_h
    port map (
            O => \N__33519\,
            I => \N__33513\
        );

    \I__8152\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33510\
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__33513\,
            I => data_in_8_3
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__33510\,
            I => data_in_8_3
        );

    \I__8149\ : InMux
    port map (
            O => \N__33505\,
            I => \N__33502\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33498\
        );

    \I__8147\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33495\
        );

    \I__8146\ : Span4Mux_s1_v
    port map (
            O => \N__33498\,
            I => \N__33490\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33490\
        );

    \I__8144\ : Span4Mux_h
    port map (
            O => \N__33490\,
            I => \N__33486\
        );

    \I__8143\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33483\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__33486\,
            I => data_in_7_3
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__33483\,
            I => data_in_7_3
        );

    \I__8140\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33473\
        );

    \I__8139\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33470\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__33476\,
            I => \N__33467\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__33473\,
            I => \N__33464\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__33470\,
            I => \N__33461\
        );

    \I__8135\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33458\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__33464\,
            I => \N__33455\
        );

    \I__8133\ : Span4Mux_h
    port map (
            O => \N__33461\,
            I => \N__33449\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__33458\,
            I => \N__33449\
        );

    \I__8131\ : Span4Mux_h
    port map (
            O => \N__33455\,
            I => \N__33446\
        );

    \I__8130\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33443\
        );

    \I__8129\ : Span4Mux_v
    port map (
            O => \N__33449\,
            I => \N__33440\
        );

    \I__8128\ : Odrv4
    port map (
            O => \N__33446\,
            I => data_in_18_0
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__33443\,
            I => data_in_18_0
        );

    \I__8126\ : Odrv4
    port map (
            O => \N__33440\,
            I => data_in_18_0
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__33433\,
            I => \N__33429\
        );

    \I__8124\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33426\
        );

    \I__8123\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33423\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33420\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__33423\,
            I => \N__33416\
        );

    \I__8120\ : Span4Mux_v
    port map (
            O => \N__33420\,
            I => \N__33413\
        );

    \I__8119\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33410\
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__33416\,
            I => data_in_17_0
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__33413\,
            I => data_in_17_0
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__33410\,
            I => data_in_17_0
        );

    \I__8115\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33399\
        );

    \I__8114\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33395\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__33399\,
            I => \N__33390\
        );

    \I__8112\ : InMux
    port map (
            O => \N__33398\,
            I => \N__33387\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__33395\,
            I => \N__33384\
        );

    \I__8110\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33381\
        );

    \I__8109\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33378\
        );

    \I__8108\ : Span4Mux_h
    port map (
            O => \N__33390\,
            I => \N__33375\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__33387\,
            I => \N__33368\
        );

    \I__8106\ : Span4Mux_v
    port map (
            O => \N__33384\,
            I => \N__33368\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__33381\,
            I => \N__33368\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__33378\,
            I => \c0.data_in_field_118\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__33375\,
            I => \c0.data_in_field_118\
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__33368\,
            I => \c0.data_in_field_118\
        );

    \I__8101\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33356\
        );

    \I__8100\ : CascadeMux
    port map (
            O => \N__33360\,
            I => \N__33353\
        );

    \I__8099\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33350\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33347\
        );

    \I__8097\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33343\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33340\
        );

    \I__8095\ : Span12Mux_h
    port map (
            O => \N__33347\,
            I => \N__33336\
        );

    \I__8094\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33333\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__33343\,
            I => \N__33328\
        );

    \I__8092\ : Span4Mux_h
    port map (
            O => \N__33340\,
            I => \N__33328\
        );

    \I__8091\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33325\
        );

    \I__8090\ : Odrv12
    port map (
            O => \N__33336\,
            I => \c0.data_in_field_126\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__33333\,
            I => \c0.data_in_field_126\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__33328\,
            I => \c0.data_in_field_126\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__33325\,
            I => \c0.data_in_field_126\
        );

    \I__8086\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33312\
        );

    \I__8085\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33306\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__33312\,
            I => \N__33303\
        );

    \I__8083\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33300\
        );

    \I__8082\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33295\
        );

    \I__8081\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33291\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__33306\,
            I => \N__33282\
        );

    \I__8079\ : Span4Mux_v
    port map (
            O => \N__33303\,
            I => \N__33277\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__33300\,
            I => \N__33277\
        );

    \I__8077\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33267\
        );

    \I__8076\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33264\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__33295\,
            I => \N__33260\
        );

    \I__8074\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33257\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__33291\,
            I => \N__33253\
        );

    \I__8072\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33250\
        );

    \I__8071\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33247\
        );

    \I__8070\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33241\
        );

    \I__8069\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33241\
        );

    \I__8068\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33238\
        );

    \I__8067\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33233\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__33282\,
            I => \N__33228\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__33277\,
            I => \N__33228\
        );

    \I__8064\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33223\
        );

    \I__8063\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33223\
        );

    \I__8062\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33218\
        );

    \I__8061\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33213\
        );

    \I__8060\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33213\
        );

    \I__8059\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33209\
        );

    \I__8058\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33206\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__33267\,
            I => \N__33203\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__33264\,
            I => \N__33198\
        );

    \I__8055\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33195\
        );

    \I__8054\ : Span4Mux_h
    port map (
            O => \N__33260\,
            I => \N__33190\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__33257\,
            I => \N__33190\
        );

    \I__8052\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33187\
        );

    \I__8051\ : Span4Mux_s2_v
    port map (
            O => \N__33253\,
            I => \N__33174\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__33250\,
            I => \N__33174\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__33247\,
            I => \N__33174\
        );

    \I__8048\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33171\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33168\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33165\
        );

    \I__8045\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33162\
        );

    \I__8044\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33159\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__33233\,
            I => \N__33152\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__33228\,
            I => \N__33152\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__33223\,
            I => \N__33152\
        );

    \I__8040\ : InMux
    port map (
            O => \N__33222\,
            I => \N__33149\
        );

    \I__8039\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33146\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__33218\,
            I => \N__33143\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__33213\,
            I => \N__33140\
        );

    \I__8036\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33135\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__33209\,
            I => \N__33128\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33128\
        );

    \I__8033\ : Span4Mux_v
    port map (
            O => \N__33203\,
            I => \N__33128\
        );

    \I__8032\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33123\
        );

    \I__8031\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33123\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__33198\,
            I => \N__33118\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33118\
        );

    \I__8028\ : Span4Mux_v
    port map (
            O => \N__33190\,
            I => \N__33112\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__33187\,
            I => \N__33109\
        );

    \I__8026\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33104\
        );

    \I__8025\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33104\
        );

    \I__8024\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33101\
        );

    \I__8023\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33096\
        );

    \I__8022\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33096\
        );

    \I__8021\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33093\
        );

    \I__8020\ : Span4Mux_v
    port map (
            O => \N__33174\,
            I => \N__33090\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__33171\,
            I => \N__33079\
        );

    \I__8018\ : Span4Mux_s2_h
    port map (
            O => \N__33168\,
            I => \N__33079\
        );

    \I__8017\ : Span4Mux_h
    port map (
            O => \N__33165\,
            I => \N__33079\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__33162\,
            I => \N__33079\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__33159\,
            I => \N__33079\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__33152\,
            I => \N__33076\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__33149\,
            I => \N__33067\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__33146\,
            I => \N__33067\
        );

    \I__8011\ : Span4Mux_h
    port map (
            O => \N__33143\,
            I => \N__33067\
        );

    \I__8010\ : Span4Mux_v
    port map (
            O => \N__33140\,
            I => \N__33067\
        );

    \I__8009\ : InMux
    port map (
            O => \N__33139\,
            I => \N__33062\
        );

    \I__8008\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33062\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__33135\,
            I => \N__33053\
        );

    \I__8006\ : Span4Mux_h
    port map (
            O => \N__33128\,
            I => \N__33053\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__33123\,
            I => \N__33053\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__33118\,
            I => \N__33053\
        );

    \I__8003\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33050\
        );

    \I__8002\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33047\
        );

    \I__8001\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33044\
        );

    \I__8000\ : Sp12to4
    port map (
            O => \N__33112\,
            I => \N__33033\
        );

    \I__7999\ : Span12Mux_s8_v
    port map (
            O => \N__33109\,
            I => \N__33033\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__33104\,
            I => \N__33033\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__33101\,
            I => \N__33033\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__33096\,
            I => \N__33033\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__33093\,
            I => \N__33024\
        );

    \I__7994\ : Span4Mux_h
    port map (
            O => \N__33090\,
            I => \N__33024\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__33079\,
            I => \N__33024\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__33076\,
            I => \N__33024\
        );

    \I__7991\ : Span4Mux_v
    port map (
            O => \N__33067\,
            I => \N__33017\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33017\
        );

    \I__7989\ : Span4Mux_h
    port map (
            O => \N__33053\,
            I => \N__33017\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__33050\,
            I => \N__33014\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__33047\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__33044\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7985\ : Odrv12
    port map (
            O => \N__33033\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__33024\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__33017\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7982\ : Odrv12
    port map (
            O => \N__33014\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7981\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__32995\,
            I => \N__32991\
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__32994\,
            I => \N__32987\
        );

    \I__7977\ : Sp12to4
    port map (
            O => \N__32991\,
            I => \N__32982\
        );

    \I__7976\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32979\
        );

    \I__7975\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32972\
        );

    \I__7974\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32972\
        );

    \I__7973\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32972\
        );

    \I__7972\ : Odrv12
    port map (
            O => \N__32982\,
            I => \c0.data_in_field_86\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__32979\,
            I => \c0.data_in_field_86\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__32972\,
            I => \c0.data_in_field_86\
        );

    \I__7969\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32961\
        );

    \I__7968\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32957\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__32961\,
            I => \N__32954\
        );

    \I__7966\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32951\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__32957\,
            I => \N__32947\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__32954\,
            I => \N__32942\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__32951\,
            I => \N__32942\
        );

    \I__7962\ : CascadeMux
    port map (
            O => \N__32950\,
            I => \N__32939\
        );

    \I__7961\ : Span4Mux_v
    port map (
            O => \N__32947\,
            I => \N__32933\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__32942\,
            I => \N__32933\
        );

    \I__7959\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32930\
        );

    \I__7958\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32927\
        );

    \I__7957\ : Span4Mux_h
    port map (
            O => \N__32933\,
            I => \N__32924\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__32930\,
            I => \N__32921\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__32927\,
            I => \c0.data_in_field_94\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__32924\,
            I => \c0.data_in_field_94\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__32921\,
            I => \c0.data_in_field_94\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__32914\,
            I => \N__32910\
        );

    \I__7951\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32906\
        );

    \I__7950\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32903\
        );

    \I__7949\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32900\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32897\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__32903\,
            I => \N__32894\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__32900\,
            I => \N__32890\
        );

    \I__7945\ : Span4Mux_v
    port map (
            O => \N__32897\,
            I => \N__32884\
        );

    \I__7944\ : Span4Mux_v
    port map (
            O => \N__32894\,
            I => \N__32884\
        );

    \I__7943\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32881\
        );

    \I__7942\ : Span4Mux_v
    port map (
            O => \N__32890\,
            I => \N__32878\
        );

    \I__7941\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32875\
        );

    \I__7940\ : Sp12to4
    port map (
            O => \N__32884\,
            I => \N__32872\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__32881\,
            I => \c0.data_in_field_70\
        );

    \I__7938\ : Odrv4
    port map (
            O => \N__32878\,
            I => \c0.data_in_field_70\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__32875\,
            I => \c0.data_in_field_70\
        );

    \I__7936\ : Odrv12
    port map (
            O => \N__32872\,
            I => \c0.data_in_field_70\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__32863\,
            I => \c0.n5899_cascade_\
        );

    \I__7934\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32857\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32854\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__32854\,
            I => \N__32849\
        );

    \I__7931\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32844\
        );

    \I__7930\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32844\
        );

    \I__7929\ : Odrv4
    port map (
            O => \N__32849\,
            I => \c0.data_in_field_78\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__32844\,
            I => \c0.data_in_field_78\
        );

    \I__7927\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32836\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32833\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__32833\,
            I => \c0.n5893\
        );

    \I__7924\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32826\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__32829\,
            I => \N__32822\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__32826\,
            I => \N__32819\
        );

    \I__7921\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32816\
        );

    \I__7920\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32813\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__32819\,
            I => \N__32810\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32806\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__32813\,
            I => \N__32801\
        );

    \I__7916\ : Span4Mux_h
    port map (
            O => \N__32810\,
            I => \N__32801\
        );

    \I__7915\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32798\
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__32806\,
            I => \c0.data_in_field_102\
        );

    \I__7913\ : Odrv4
    port map (
            O => \N__32801\,
            I => \c0.data_in_field_102\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__32798\,
            I => \c0.data_in_field_102\
        );

    \I__7911\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32786\
        );

    \I__7910\ : CascadeMux
    port map (
            O => \N__32790\,
            I => \N__32782\
        );

    \I__7909\ : CascadeMux
    port map (
            O => \N__32789\,
            I => \N__32779\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__32786\,
            I => \N__32772\
        );

    \I__7907\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32769\
        );

    \I__7906\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32766\
        );

    \I__7905\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32763\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__32778\,
            I => \N__32760\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__32777\,
            I => \N__32757\
        );

    \I__7902\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32750\
        );

    \I__7901\ : InMux
    port map (
            O => \N__32775\,
            I => \N__32750\
        );

    \I__7900\ : Span4Mux_h
    port map (
            O => \N__32772\,
            I => \N__32741\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__32769\,
            I => \N__32741\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__32766\,
            I => \N__32741\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__32763\,
            I => \N__32741\
        );

    \I__7896\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32736\
        );

    \I__7895\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32736\
        );

    \I__7894\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32730\
        );

    \I__7893\ : InMux
    port map (
            O => \N__32755\,
            I => \N__32727\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__32750\,
            I => \N__32720\
        );

    \I__7891\ : Span4Mux_v
    port map (
            O => \N__32741\,
            I => \N__32720\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__32736\,
            I => \N__32720\
        );

    \I__7889\ : CascadeMux
    port map (
            O => \N__32735\,
            I => \N__32717\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__32734\,
            I => \N__32714\
        );

    \I__7887\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32709\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__32730\,
            I => \N__32702\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32702\
        );

    \I__7884\ : Span4Mux_v
    port map (
            O => \N__32720\,
            I => \N__32702\
        );

    \I__7883\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32699\
        );

    \I__7882\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32691\
        );

    \I__7881\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32691\
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__32712\,
            I => \N__32688\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__32709\,
            I => \N__32685\
        );

    \I__7878\ : Span4Mux_v
    port map (
            O => \N__32702\,
            I => \N__32680\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__32699\,
            I => \N__32680\
        );

    \I__7876\ : CascadeMux
    port map (
            O => \N__32698\,
            I => \N__32675\
        );

    \I__7875\ : CascadeMux
    port map (
            O => \N__32697\,
            I => \N__32671\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__32696\,
            I => \N__32668\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__32691\,
            I => \N__32663\
        );

    \I__7872\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32660\
        );

    \I__7871\ : Span4Mux_s3_v
    port map (
            O => \N__32685\,
            I => \N__32652\
        );

    \I__7870\ : Span4Mux_s3_v
    port map (
            O => \N__32680\,
            I => \N__32652\
        );

    \I__7869\ : CascadeMux
    port map (
            O => \N__32679\,
            I => \N__32649\
        );

    \I__7868\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \N__32646\
        );

    \I__7867\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32643\
        );

    \I__7866\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32634\
        );

    \I__7865\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32634\
        );

    \I__7864\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32634\
        );

    \I__7863\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32634\
        );

    \I__7862\ : CascadeMux
    port map (
            O => \N__32666\,
            I => \N__32631\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__32663\,
            I => \N__32622\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32622\
        );

    \I__7859\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32619\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__32658\,
            I => \N__32616\
        );

    \I__7857\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32613\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__32652\,
            I => \N__32610\
        );

    \I__7855\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32607\
        );

    \I__7854\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32604\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__32643\,
            I => \N__32599\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__32634\,
            I => \N__32599\
        );

    \I__7851\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32596\
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__32630\,
            I => \N__32590\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__32629\,
            I => \N__32583\
        );

    \I__7848\ : CascadeMux
    port map (
            O => \N__32628\,
            I => \N__32577\
        );

    \I__7847\ : CascadeMux
    port map (
            O => \N__32627\,
            I => \N__32573\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__32622\,
            I => \N__32565\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__32619\,
            I => \N__32565\
        );

    \I__7844\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32561\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32554\
        );

    \I__7842\ : Span4Mux_s3_v
    port map (
            O => \N__32610\,
            I => \N__32554\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__32607\,
            I => \N__32554\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32547\
        );

    \I__7839\ : Span4Mux_v
    port map (
            O => \N__32599\,
            I => \N__32547\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32547\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__32595\,
            I => \N__32540\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \N__32537\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__32593\,
            I => \N__32534\
        );

    \I__7834\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32531\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__32589\,
            I => \N__32528\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__32588\,
            I => \N__32519\
        );

    \I__7831\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32513\
        );

    \I__7830\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32508\
        );

    \I__7829\ : InMux
    port map (
            O => \N__32583\,
            I => \N__32508\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__32582\,
            I => \N__32499\
        );

    \I__7827\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32496\
        );

    \I__7826\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32493\
        );

    \I__7825\ : InMux
    port map (
            O => \N__32577\,
            I => \N__32490\
        );

    \I__7824\ : InMux
    port map (
            O => \N__32576\,
            I => \N__32487\
        );

    \I__7823\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32484\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__32572\,
            I => \N__32480\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__32571\,
            I => \N__32477\
        );

    \I__7820\ : CascadeMux
    port map (
            O => \N__32570\,
            I => \N__32472\
        );

    \I__7819\ : Span4Mux_h
    port map (
            O => \N__32565\,
            I => \N__32469\
        );

    \I__7818\ : CascadeMux
    port map (
            O => \N__32564\,
            I => \N__32466\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__32561\,
            I => \N__32461\
        );

    \I__7816\ : Span4Mux_v
    port map (
            O => \N__32554\,
            I => \N__32458\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__32547\,
            I => \N__32455\
        );

    \I__7814\ : CascadeMux
    port map (
            O => \N__32546\,
            I => \N__32451\
        );

    \I__7813\ : CascadeMux
    port map (
            O => \N__32545\,
            I => \N__32448\
        );

    \I__7812\ : CascadeMux
    port map (
            O => \N__32544\,
            I => \N__32440\
        );

    \I__7811\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32437\
        );

    \I__7810\ : InMux
    port map (
            O => \N__32540\,
            I => \N__32434\
        );

    \I__7809\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32429\
        );

    \I__7808\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32429\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32426\
        );

    \I__7806\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32423\
        );

    \I__7805\ : InMux
    port map (
            O => \N__32527\,
            I => \N__32418\
        );

    \I__7804\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32418\
        );

    \I__7803\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32413\
        );

    \I__7802\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32413\
        );

    \I__7801\ : InMux
    port map (
            O => \N__32523\,
            I => \N__32407\
        );

    \I__7800\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32407\
        );

    \I__7799\ : InMux
    port map (
            O => \N__32519\,
            I => \N__32404\
        );

    \I__7798\ : InMux
    port map (
            O => \N__32518\,
            I => \N__32401\
        );

    \I__7797\ : InMux
    port map (
            O => \N__32517\,
            I => \N__32396\
        );

    \I__7796\ : InMux
    port map (
            O => \N__32516\,
            I => \N__32396\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__32513\,
            I => \N__32391\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__32508\,
            I => \N__32391\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__32507\,
            I => \N__32388\
        );

    \I__7792\ : CascadeMux
    port map (
            O => \N__32506\,
            I => \N__32385\
        );

    \I__7791\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32382\
        );

    \I__7790\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32373\
        );

    \I__7789\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32373\
        );

    \I__7788\ : InMux
    port map (
            O => \N__32502\,
            I => \N__32373\
        );

    \I__7787\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32373\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__32496\,
            I => \N__32366\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__32493\,
            I => \N__32366\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__32490\,
            I => \N__32366\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__32487\,
            I => \N__32361\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__32484\,
            I => \N__32361\
        );

    \I__7781\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32356\
        );

    \I__7780\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32356\
        );

    \I__7779\ : InMux
    port map (
            O => \N__32477\,
            I => \N__32351\
        );

    \I__7778\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32351\
        );

    \I__7777\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32346\
        );

    \I__7776\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32346\
        );

    \I__7775\ : Sp12to4
    port map (
            O => \N__32469\,
            I => \N__32343\
        );

    \I__7774\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32340\
        );

    \I__7773\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32337\
        );

    \I__7772\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32334\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__32461\,
            I => \N__32329\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__32458\,
            I => \N__32329\
        );

    \I__7769\ : Span4Mux_v
    port map (
            O => \N__32455\,
            I => \N__32326\
        );

    \I__7768\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32321\
        );

    \I__7767\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32321\
        );

    \I__7766\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32312\
        );

    \I__7765\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32309\
        );

    \I__7764\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32306\
        );

    \I__7763\ : InMux
    port map (
            O => \N__32445\,
            I => \N__32297\
        );

    \I__7762\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32297\
        );

    \I__7761\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32297\
        );

    \I__7760\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32297\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__32437\,
            I => \N__32286\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__32434\,
            I => \N__32286\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__32429\,
            I => \N__32286\
        );

    \I__7756\ : Span4Mux_h
    port map (
            O => \N__32426\,
            I => \N__32286\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32286\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32281\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__32413\,
            I => \N__32281\
        );

    \I__7752\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32278\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32267\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__32404\,
            I => \N__32267\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__32401\,
            I => \N__32267\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__32396\,
            I => \N__32267\
        );

    \I__7747\ : Span4Mux_v
    port map (
            O => \N__32391\,
            I => \N__32267\
        );

    \I__7746\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32262\
        );

    \I__7745\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32262\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__32382\,
            I => \N__32251\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__32373\,
            I => \N__32251\
        );

    \I__7742\ : Span4Mux_v
    port map (
            O => \N__32366\,
            I => \N__32251\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__32361\,
            I => \N__32251\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__32356\,
            I => \N__32251\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32232\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32232\
        );

    \I__7737\ : Span12Mux_s7_v
    port map (
            O => \N__32343\,
            I => \N__32232\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__32340\,
            I => \N__32232\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__32337\,
            I => \N__32232\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__32334\,
            I => \N__32232\
        );

    \I__7733\ : Sp12to4
    port map (
            O => \N__32329\,
            I => \N__32232\
        );

    \I__7732\ : Sp12to4
    port map (
            O => \N__32326\,
            I => \N__32232\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__32321\,
            I => \N__32232\
        );

    \I__7730\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32229\
        );

    \I__7729\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32226\
        );

    \I__7728\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32221\
        );

    \I__7727\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32221\
        );

    \I__7726\ : InMux
    port map (
            O => \N__32316\,
            I => \N__32218\
        );

    \I__7725\ : InMux
    port map (
            O => \N__32315\,
            I => \N__32215\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__32312\,
            I => \N__32212\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32203\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32203\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__32297\,
            I => \N__32203\
        );

    \I__7720\ : Span4Mux_v
    port map (
            O => \N__32286\,
            I => \N__32203\
        );

    \I__7719\ : Span4Mux_v
    port map (
            O => \N__32281\,
            I => \N__32192\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__32278\,
            I => \N__32192\
        );

    \I__7717\ : Span4Mux_v
    port map (
            O => \N__32267\,
            I => \N__32192\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32192\
        );

    \I__7715\ : Span4Mux_h
    port map (
            O => \N__32251\,
            I => \N__32192\
        );

    \I__7714\ : Span12Mux_h
    port map (
            O => \N__32232\,
            I => \N__32189\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__32229\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__32226\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__32221\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__32218\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__32215\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7708\ : Odrv12
    port map (
            O => \N__32212\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7707\ : Odrv4
    port map (
            O => \N__32203\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7706\ : Odrv4
    port map (
            O => \N__32192\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7705\ : Odrv12
    port map (
            O => \N__32189\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7704\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32167\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__32167\,
            I => \N__32163\
        );

    \I__7702\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32158\
        );

    \I__7701\ : Span4Mux_h
    port map (
            O => \N__32163\,
            I => \N__32155\
        );

    \I__7700\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32152\
        );

    \I__7699\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32149\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__32158\,
            I => \c0.data_in_field_110\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__32155\,
            I => \c0.data_in_field_110\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__32152\,
            I => \c0.data_in_field_110\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__32149\,
            I => \c0.data_in_field_110\
        );

    \I__7694\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32137\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__32137\,
            I => \c0.n5384\
        );

    \I__7692\ : CascadeMux
    port map (
            O => \N__32134\,
            I => \c0.n5387_cascade_\
        );

    \I__7691\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32128\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__32128\,
            I => \N__32125\
        );

    \I__7689\ : Span4Mux_v
    port map (
            O => \N__32125\,
            I => \N__32119\
        );

    \I__7688\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32116\
        );

    \I__7687\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32112\
        );

    \I__7686\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32109\
        );

    \I__7685\ : Span4Mux_h
    port map (
            O => \N__32119\,
            I => \N__32103\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__32116\,
            I => \N__32103\
        );

    \I__7683\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32100\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__32112\,
            I => \N__32092\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__32109\,
            I => \N__32092\
        );

    \I__7680\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32089\
        );

    \I__7679\ : Span4Mux_h
    port map (
            O => \N__32103\,
            I => \N__32086\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__32100\,
            I => \N__32083\
        );

    \I__7677\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32080\
        );

    \I__7676\ : InMux
    port map (
            O => \N__32098\,
            I => \N__32076\
        );

    \I__7675\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32073\
        );

    \I__7674\ : Span4Mux_v
    port map (
            O => \N__32092\,
            I => \N__32070\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32061\
        );

    \I__7672\ : Span4Mux_h
    port map (
            O => \N__32086\,
            I => \N__32061\
        );

    \I__7671\ : Span4Mux_s2_h
    port map (
            O => \N__32083\,
            I => \N__32061\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__32080\,
            I => \N__32061\
        );

    \I__7669\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32058\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__32076\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__32073\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__32070\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7665\ : Odrv4
    port map (
            O => \N__32061\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__32058\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7663\ : InMux
    port map (
            O => \N__32047\,
            I => \N__32044\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__32044\,
            I => \N__32041\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__32041\,
            I => \c0.n5378\
        );

    \I__7660\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32035\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__32032\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__32032\,
            I => \N__32029\
        );

    \I__7657\ : Odrv4
    port map (
            O => \N__32029\,
            I => \c0.n5381\
        );

    \I__7656\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32023\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__32023\,
            I => \N__32019\
        );

    \I__7654\ : InMux
    port map (
            O => \N__32022\,
            I => \N__32016\
        );

    \I__7653\ : Span4Mux_s2_h
    port map (
            O => \N__32019\,
            I => \N__32011\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32011\
        );

    \I__7651\ : Span4Mux_v
    port map (
            O => \N__32011\,
            I => \N__32007\
        );

    \I__7650\ : InMux
    port map (
            O => \N__32010\,
            I => \N__32003\
        );

    \I__7649\ : Span4Mux_h
    port map (
            O => \N__32007\,
            I => \N__32000\
        );

    \I__7648\ : InMux
    port map (
            O => \N__32006\,
            I => \N__31996\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__32003\,
            I => \N__31993\
        );

    \I__7646\ : Span4Mux_h
    port map (
            O => \N__32000\,
            I => \N__31990\
        );

    \I__7645\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31987\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__31996\,
            I => \c0.data_in_field_136\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__31993\,
            I => \c0.data_in_field_136\
        );

    \I__7642\ : Odrv4
    port map (
            O => \N__31990\,
            I => \c0.data_in_field_136\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__31987\,
            I => \c0.data_in_field_136\
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__31978\,
            I => \N__31975\
        );

    \I__7639\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31972\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__31972\,
            I => \N__31969\
        );

    \I__7637\ : Span4Mux_v
    port map (
            O => \N__31969\,
            I => \N__31964\
        );

    \I__7636\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31959\
        );

    \I__7635\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31959\
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__31964\,
            I => data_in_15_2
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__31959\,
            I => data_in_15_2
        );

    \I__7632\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31950\
        );

    \I__7631\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31947\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31943\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__31947\,
            I => \N__31940\
        );

    \I__7628\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31937\
        );

    \I__7627\ : Span4Mux_h
    port map (
            O => \N__31943\,
            I => \N__31933\
        );

    \I__7626\ : Span4Mux_v
    port map (
            O => \N__31940\,
            I => \N__31926\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31926\
        );

    \I__7624\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31923\
        );

    \I__7623\ : Span4Mux_h
    port map (
            O => \N__31933\,
            I => \N__31920\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__31932\,
            I => \N__31917\
        );

    \I__7621\ : InMux
    port map (
            O => \N__31931\,
            I => \N__31914\
        );

    \I__7620\ : Span4Mux_h
    port map (
            O => \N__31926\,
            I => \N__31911\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__31923\,
            I => \N__31906\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__31920\,
            I => \N__31906\
        );

    \I__7617\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31903\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__31914\,
            I => \c0.data_in_field_122\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__31911\,
            I => \c0.data_in_field_122\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__31906\,
            I => \c0.data_in_field_122\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__31903\,
            I => \c0.data_in_field_122\
        );

    \I__7612\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31891\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__31891\,
            I => \N__31888\
        );

    \I__7610\ : Span4Mux_h
    port map (
            O => \N__31888\,
            I => \N__31885\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__31885\,
            I => \N__31880\
        );

    \I__7608\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31875\
        );

    \I__7607\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31875\
        );

    \I__7606\ : Odrv4
    port map (
            O => \N__31880\,
            I => data_in_14_3
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__31875\,
            I => data_in_14_3
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__31870\,
            I => \N__31867\
        );

    \I__7603\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31864\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__31864\,
            I => \N__31861\
        );

    \I__7601\ : Span4Mux_h
    port map (
            O => \N__31861\,
            I => \N__31858\
        );

    \I__7600\ : Span4Mux_v
    port map (
            O => \N__31858\,
            I => \N__31855\
        );

    \I__7599\ : Span4Mux_h
    port map (
            O => \N__31855\,
            I => \N__31850\
        );

    \I__7598\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31845\
        );

    \I__7597\ : InMux
    port map (
            O => \N__31853\,
            I => \N__31845\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__31850\,
            I => data_in_13_3
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__31845\,
            I => data_in_13_3
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__31840\,
            I => \N__31837\
        );

    \I__7593\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31834\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__7591\ : Span4Mux_h
    port map (
            O => \N__31831\,
            I => \N__31828\
        );

    \I__7590\ : Span4Mux_h
    port map (
            O => \N__31828\,
            I => \N__31825\
        );

    \I__7589\ : Span4Mux_h
    port map (
            O => \N__31825\,
            I => \N__31820\
        );

    \I__7588\ : InMux
    port map (
            O => \N__31824\,
            I => \N__31815\
        );

    \I__7587\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31815\
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__31820\,
            I => data_in_12_3
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__31815\,
            I => data_in_12_3
        );

    \I__7584\ : InMux
    port map (
            O => \N__31810\,
            I => \N__31807\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__31807\,
            I => \N__31803\
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__31806\,
            I => \N__31800\
        );

    \I__7581\ : Span4Mux_h
    port map (
            O => \N__31803\,
            I => \N__31796\
        );

    \I__7580\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31791\
        );

    \I__7579\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31791\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__31796\,
            I => data_in_11_3
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__31791\,
            I => data_in_11_3
        );

    \I__7576\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31782\
        );

    \I__7575\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31779\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__31782\,
            I => \N__31776\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31772\
        );

    \I__7572\ : Span4Mux_h
    port map (
            O => \N__31776\,
            I => \N__31769\
        );

    \I__7571\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31764\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__31772\,
            I => \N__31759\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__31769\,
            I => \N__31759\
        );

    \I__7568\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31756\
        );

    \I__7567\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31753\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__31764\,
            I => \c0.data_in_field_91\
        );

    \I__7565\ : Odrv4
    port map (
            O => \N__31759\,
            I => \c0.data_in_field_91\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__31756\,
            I => \c0.data_in_field_91\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__31753\,
            I => \c0.data_in_field_91\
        );

    \I__7562\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31741\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__31741\,
            I => \N__31738\
        );

    \I__7560\ : Span4Mux_v
    port map (
            O => \N__31738\,
            I => \N__31735\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__31735\,
            I => \N__31732\
        );

    \I__7558\ : Span4Mux_h
    port map (
            O => \N__31732\,
            I => \N__31727\
        );

    \I__7557\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31724\
        );

    \I__7556\ : InMux
    port map (
            O => \N__31730\,
            I => \N__31721\
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__31727\,
            I => data_in_0_3
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__31724\,
            I => data_in_0_3
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__31721\,
            I => data_in_0_3
        );

    \I__7552\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31711\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__31711\,
            I => \N__31706\
        );

    \I__7550\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31703\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__31709\,
            I => \N__31700\
        );

    \I__7548\ : Span4Mux_h
    port map (
            O => \N__31706\,
            I => \N__31697\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__31703\,
            I => \N__31694\
        );

    \I__7546\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31690\
        );

    \I__7545\ : Span4Mux_h
    port map (
            O => \N__31697\,
            I => \N__31687\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__31694\,
            I => \N__31684\
        );

    \I__7543\ : InMux
    port map (
            O => \N__31693\,
            I => \N__31681\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__31690\,
            I => \c0.data_in_field_3\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__31687\,
            I => \c0.data_in_field_3\
        );

    \I__7540\ : Odrv4
    port map (
            O => \N__31684\,
            I => \c0.data_in_field_3\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__31681\,
            I => \c0.data_in_field_3\
        );

    \I__7538\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31668\
        );

    \I__7537\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31665\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31662\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__31665\,
            I => \N__31659\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__31662\,
            I => \N__31656\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__31659\,
            I => \N__31653\
        );

    \I__7532\ : Span4Mux_h
    port map (
            O => \N__31656\,
            I => \N__31647\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__31653\,
            I => \N__31647\
        );

    \I__7530\ : InMux
    port map (
            O => \N__31652\,
            I => \N__31644\
        );

    \I__7529\ : Odrv4
    port map (
            O => \N__31647\,
            I => data_in_11_2
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__31644\,
            I => data_in_11_2
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__31639\,
            I => \N__31636\
        );

    \I__7526\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__31633\,
            I => \N__31630\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__31630\,
            I => \N__31627\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__31627\,
            I => \N__31624\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__31624\,
            I => \N__31619\
        );

    \I__7521\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31614\
        );

    \I__7520\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31614\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__31619\,
            I => data_in_10_2
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__31614\,
            I => data_in_10_2
        );

    \I__7517\ : CascadeMux
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__7516\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__7514\ : Span4Mux_v
    port map (
            O => \N__31600\,
            I => \N__31595\
        );

    \I__7513\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31590\
        );

    \I__7512\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31590\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__31595\,
            I => data_in_5_4
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__31590\,
            I => data_in_5_4
        );

    \I__7509\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31582\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__7507\ : Span4Mux_v
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__7506\ : Span4Mux_h
    port map (
            O => \N__31576\,
            I => \N__31571\
        );

    \I__7505\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31568\
        );

    \I__7504\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31565\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__31571\,
            I => \N__31560\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31560\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__31565\,
            I => \c0.data_in_field_44\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__31560\,
            I => \c0.data_in_field_44\
        );

    \I__7499\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31551\
        );

    \I__7498\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31548\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31543\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__31548\,
            I => \N__31543\
        );

    \I__7495\ : Span4Mux_v
    port map (
            O => \N__31543\,
            I => \N__31539\
        );

    \I__7494\ : InMux
    port map (
            O => \N__31542\,
            I => \N__31536\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__31539\,
            I => \N__31531\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__31536\,
            I => \N__31531\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__31531\,
            I => \c0.n1962\
        );

    \I__7490\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31525\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__31525\,
            I => \N__31521\
        );

    \I__7488\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31518\
        );

    \I__7487\ : Span4Mux_s3_v
    port map (
            O => \N__31521\,
            I => \N__31514\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31510\
        );

    \I__7485\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31507\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__31514\,
            I => \N__31504\
        );

    \I__7483\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31501\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__31510\,
            I => \N__31496\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__31507\,
            I => \N__31496\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__31504\,
            I => data_in_3_0
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__31501\,
            I => data_in_3_0
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__31496\,
            I => data_in_3_0
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__31489\,
            I => \N__31485\
        );

    \I__7476\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31482\
        );

    \I__7475\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31477\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__31482\,
            I => \N__31474\
        );

    \I__7473\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31471\
        );

    \I__7472\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31468\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__31477\,
            I => \c0.data_in_field_24\
        );

    \I__7470\ : Odrv4
    port map (
            O => \N__31474\,
            I => \c0.data_in_field_24\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__31471\,
            I => \c0.data_in_field_24\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__31468\,
            I => \c0.data_in_field_24\
        );

    \I__7467\ : CascadeMux
    port map (
            O => \N__31459\,
            I => \N__31455\
        );

    \I__7466\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31452\
        );

    \I__7465\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31449\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N__31446\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__31449\,
            I => \N__31441\
        );

    \I__7462\ : Span4Mux_h
    port map (
            O => \N__31446\,
            I => \N__31441\
        );

    \I__7461\ : Span4Mux_h
    port map (
            O => \N__31441\,
            I => \N__31436\
        );

    \I__7460\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31433\
        );

    \I__7459\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31430\
        );

    \I__7458\ : Span4Mux_h
    port map (
            O => \N__31436\,
            I => \N__31427\
        );

    \I__7457\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31424\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__31430\,
            I => data_in_2_0
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__31427\,
            I => data_in_2_0
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__31424\,
            I => data_in_2_0
        );

    \I__7453\ : InMux
    port map (
            O => \N__31417\,
            I => \N__31413\
        );

    \I__7452\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31410\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31406\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31403\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__31409\,
            I => \N__31399\
        );

    \I__7448\ : Span4Mux_v
    port map (
            O => \N__31406\,
            I => \N__31394\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__31403\,
            I => \N__31394\
        );

    \I__7446\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31391\
        );

    \I__7445\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31388\
        );

    \I__7444\ : Span4Mux_h
    port map (
            O => \N__31394\,
            I => \N__31385\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__31391\,
            I => data_in_1_0
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__31388\,
            I => data_in_1_0
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__31385\,
            I => data_in_1_0
        );

    \I__7440\ : CascadeMux
    port map (
            O => \N__31378\,
            I => \N__31375\
        );

    \I__7439\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__31372\,
            I => \N__31368\
        );

    \I__7437\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31365\
        );

    \I__7436\ : Span4Mux_h
    port map (
            O => \N__31368\,
            I => \N__31361\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31358\
        );

    \I__7434\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31355\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__31361\,
            I => data_in_15_3
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__31358\,
            I => data_in_15_3
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__31355\,
            I => data_in_15_3
        );

    \I__7430\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31345\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__31345\,
            I => \N__31341\
        );

    \I__7428\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31338\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__31341\,
            I => \N__31335\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__31338\,
            I => \N__31332\
        );

    \I__7425\ : Span4Mux_v
    port map (
            O => \N__31335\,
            I => \N__31327\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__31332\,
            I => \N__31324\
        );

    \I__7423\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31321\
        );

    \I__7422\ : InMux
    port map (
            O => \N__31330\,
            I => \N__31318\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__31327\,
            I => \N__31313\
        );

    \I__7420\ : Span4Mux_h
    port map (
            O => \N__31324\,
            I => \N__31313\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__31321\,
            I => \c0.data_in_field_123\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__31318\,
            I => \c0.data_in_field_123\
        );

    \I__7417\ : Odrv4
    port map (
            O => \N__31313\,
            I => \c0.data_in_field_123\
        );

    \I__7416\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31300\
        );

    \I__7415\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31300\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__31300\,
            I => \N__31296\
        );

    \I__7413\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31293\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__31296\,
            I => data_in_12_6
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__31293\,
            I => data_in_12_6
        );

    \I__7410\ : CascadeMux
    port map (
            O => \N__31288\,
            I => \N__31285\
        );

    \I__7409\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31281\
        );

    \I__7408\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31278\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31275\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__31278\,
            I => \N__31271\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__31275\,
            I => \N__31268\
        );

    \I__7404\ : InMux
    port map (
            O => \N__31274\,
            I => \N__31265\
        );

    \I__7403\ : Span12Mux_v
    port map (
            O => \N__31271\,
            I => \N__31262\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__31268\,
            I => \N__31259\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__31265\,
            I => data_in_11_6
        );

    \I__7400\ : Odrv12
    port map (
            O => \N__31262\,
            I => data_in_11_6
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__31259\,
            I => data_in_11_6
        );

    \I__7398\ : CascadeMux
    port map (
            O => \N__31252\,
            I => \N__31248\
        );

    \I__7397\ : CascadeMux
    port map (
            O => \N__31251\,
            I => \N__31244\
        );

    \I__7396\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31241\
        );

    \I__7395\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31238\
        );

    \I__7394\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31234\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31229\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__31238\,
            I => \N__31229\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__31237\,
            I => \N__31226\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__31234\,
            I => \N__31223\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__31229\,
            I => \N__31220\
        );

    \I__7388\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31217\
        );

    \I__7387\ : Sp12to4
    port map (
            O => \N__31223\,
            I => \N__31214\
        );

    \I__7386\ : Span4Mux_h
    port map (
            O => \N__31220\,
            I => \N__31211\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__31217\,
            I => data_in_18_2
        );

    \I__7384\ : Odrv12
    port map (
            O => \N__31214\,
            I => data_in_18_2
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__31211\,
            I => data_in_18_2
        );

    \I__7382\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31200\
        );

    \I__7381\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31197\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31194\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31191\
        );

    \I__7378\ : Span4Mux_v
    port map (
            O => \N__31194\,
            I => \N__31185\
        );

    \I__7377\ : Span4Mux_h
    port map (
            O => \N__31191\,
            I => \N__31185\
        );

    \I__7376\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31181\
        );

    \I__7375\ : Span4Mux_h
    port map (
            O => \N__31185\,
            I => \N__31178\
        );

    \I__7374\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31175\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__31181\,
            I => \c0.data_in_field_74\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__31178\,
            I => \c0.data_in_field_74\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__31175\,
            I => \c0.data_in_field_74\
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__31168\,
            I => \N__31165\
        );

    \I__7369\ : InMux
    port map (
            O => \N__31165\,
            I => \N__31162\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__31162\,
            I => \N__31159\
        );

    \I__7367\ : Span4Mux_s2_v
    port map (
            O => \N__31159\,
            I => \N__31156\
        );

    \I__7366\ : Span4Mux_v
    port map (
            O => \N__31156\,
            I => \N__31151\
        );

    \I__7365\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31146\
        );

    \I__7364\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31146\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__31151\,
            I => data_in_15_1
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__31146\,
            I => data_in_15_1
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__31141\,
            I => \N__31138\
        );

    \I__7360\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31134\
        );

    \I__7359\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31131\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31127\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__31124\
        );

    \I__7356\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31121\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__31127\,
            I => data_in_14_4
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__31124\,
            I => data_in_14_4
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__31121\,
            I => data_in_14_4
        );

    \I__7352\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31111\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__31111\,
            I => \N__31108\
        );

    \I__7350\ : Span12Mux_h
    port map (
            O => \N__31108\,
            I => \N__31103\
        );

    \I__7349\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31098\
        );

    \I__7348\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31098\
        );

    \I__7347\ : Odrv12
    port map (
            O => \N__31103\,
            I => \c0.data_in_field_116\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__31098\,
            I => \c0.data_in_field_116\
        );

    \I__7345\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31090\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31087\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__31087\,
            I => \N__31084\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__31084\,
            I => \N__31080\
        );

    \I__7341\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31077\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__31080\,
            I => \c0.n1815\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__31077\,
            I => \c0.n1815\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__31072\,
            I => \c0.n1815_cascade_\
        );

    \I__7337\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31065\
        );

    \I__7336\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31062\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__31065\,
            I => \N__31059\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31056\
        );

    \I__7333\ : Span4Mux_h
    port map (
            O => \N__31059\,
            I => \N__31053\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__31056\,
            I => \N__31050\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__31053\,
            I => \N__31045\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__31050\,
            I => \N__31042\
        );

    \I__7329\ : InMux
    port map (
            O => \N__31049\,
            I => \N__31037\
        );

    \I__7328\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31037\
        );

    \I__7327\ : Odrv4
    port map (
            O => \N__31045\,
            I => \c0.data_in_field_52\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__31042\,
            I => \c0.data_in_field_52\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__31037\,
            I => \c0.data_in_field_52\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__31030\,
            I => \N__31027\
        );

    \I__7323\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31024\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__31024\,
            I => \N__31021\
        );

    \I__7321\ : Span4Mux_h
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__31018\,
            I => \N__31015\
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__31015\,
            I => \c0.n27\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__31012\,
            I => \N__31009\
        );

    \I__7317\ : InMux
    port map (
            O => \N__31009\,
            I => \N__31006\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__31006\,
            I => \N__31003\
        );

    \I__7315\ : Span4Mux_h
    port map (
            O => \N__31003\,
            I => \N__31000\
        );

    \I__7314\ : Span4Mux_h
    port map (
            O => \N__31000\,
            I => \N__30996\
        );

    \I__7313\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30993\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__30996\,
            I => \N__30987\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30987\
        );

    \I__7310\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30984\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__30987\,
            I => data_in_14_1
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__30984\,
            I => data_in_14_1
        );

    \I__7307\ : InMux
    port map (
            O => \N__30979\,
            I => \N__30976\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__30976\,
            I => \N__30972\
        );

    \I__7305\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30969\
        );

    \I__7304\ : Span4Mux_v
    port map (
            O => \N__30972\,
            I => \N__30966\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__30969\,
            I => \N__30963\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__30966\,
            I => \N__30960\
        );

    \I__7301\ : Span4Mux_v
    port map (
            O => \N__30963\,
            I => \N__30957\
        );

    \I__7300\ : Span4Mux_h
    port map (
            O => \N__30960\,
            I => \N__30953\
        );

    \I__7299\ : Span4Mux_h
    port map (
            O => \N__30957\,
            I => \N__30950\
        );

    \I__7298\ : InMux
    port map (
            O => \N__30956\,
            I => \N__30947\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__30953\,
            I => data_in_13_1
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__30950\,
            I => data_in_13_1
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__30947\,
            I => data_in_13_1
        );

    \I__7294\ : CascadeMux
    port map (
            O => \N__30940\,
            I => \N__30937\
        );

    \I__7293\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30934\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__30934\,
            I => \N__30931\
        );

    \I__7291\ : Span4Mux_h
    port map (
            O => \N__30931\,
            I => \N__30926\
        );

    \I__7290\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30921\
        );

    \I__7289\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30921\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__30926\,
            I => data_in_7_0
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__30921\,
            I => data_in_7_0
        );

    \I__7286\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30912\
        );

    \I__7285\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30909\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30904\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__30909\,
            I => \N__30901\
        );

    \I__7282\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30896\
        );

    \I__7281\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30896\
        );

    \I__7280\ : Span4Mux_h
    port map (
            O => \N__30904\,
            I => \N__30893\
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__30901\,
            I => \c0.data_in_field_56\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__30896\,
            I => \c0.data_in_field_56\
        );

    \I__7277\ : Odrv4
    port map (
            O => \N__30893\,
            I => \c0.data_in_field_56\
        );

    \I__7276\ : InMux
    port map (
            O => \N__30886\,
            I => \N__30882\
        );

    \I__7275\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30879\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__30882\,
            I => \N__30876\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__30879\,
            I => \N__30873\
        );

    \I__7272\ : Span4Mux_v
    port map (
            O => \N__30876\,
            I => \N__30869\
        );

    \I__7271\ : Span4Mux_v
    port map (
            O => \N__30873\,
            I => \N__30866\
        );

    \I__7270\ : InMux
    port map (
            O => \N__30872\,
            I => \N__30862\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__30869\,
            I => \N__30857\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__30866\,
            I => \N__30857\
        );

    \I__7267\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30854\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__30862\,
            I => \N__30851\
        );

    \I__7265\ : Span4Mux_h
    port map (
            O => \N__30857\,
            I => \N__30844\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__30854\,
            I => \N__30844\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__30851\,
            I => \N__30841\
        );

    \I__7262\ : InMux
    port map (
            O => \N__30850\,
            I => \N__30836\
        );

    \I__7261\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30836\
        );

    \I__7260\ : Span4Mux_v
    port map (
            O => \N__30844\,
            I => \N__30833\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__30841\,
            I => \c0.data_in_field_129\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__30836\,
            I => \c0.data_in_field_129\
        );

    \I__7257\ : Odrv4
    port map (
            O => \N__30833\,
            I => \c0.data_in_field_129\
        );

    \I__7256\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30823\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__30823\,
            I => \N__30820\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__30820\,
            I => \N__30817\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__30817\,
            I => \c0.n15_adj_1923\
        );

    \I__7252\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30811\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30808\
        );

    \I__7250\ : Span4Mux_v
    port map (
            O => \N__30808\,
            I => \N__30803\
        );

    \I__7249\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30798\
        );

    \I__7248\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30798\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__30803\,
            I => data_in_6_2
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__30798\,
            I => data_in_6_2
        );

    \I__7245\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30789\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__30792\,
            I => \N__30784\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__30789\,
            I => \N__30781\
        );

    \I__7242\ : CascadeMux
    port map (
            O => \N__30788\,
            I => \N__30778\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__30787\,
            I => \N__30775\
        );

    \I__7240\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30772\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__30781\,
            I => \N__30769\
        );

    \I__7238\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30764\
        );

    \I__7237\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30764\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__30772\,
            I => \c0.data_in_field_50\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__30769\,
            I => \c0.data_in_field_50\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__30764\,
            I => \c0.data_in_field_50\
        );

    \I__7233\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30754\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__30754\,
            I => \N__30750\
        );

    \I__7231\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30746\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__30750\,
            I => \N__30743\
        );

    \I__7229\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30739\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30736\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__30743\,
            I => \N__30733\
        );

    \I__7226\ : InMux
    port map (
            O => \N__30742\,
            I => \N__30730\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__30739\,
            I => \c0.data_in_field_8\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__30736\,
            I => \c0.data_in_field_8\
        );

    \I__7223\ : Odrv4
    port map (
            O => \N__30733\,
            I => \c0.data_in_field_8\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__30730\,
            I => \c0.data_in_field_8\
        );

    \I__7221\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30718\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__30718\,
            I => \N__30715\
        );

    \I__7219\ : Span4Mux_h
    port map (
            O => \N__30715\,
            I => \N__30710\
        );

    \I__7218\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30705\
        );

    \I__7217\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30705\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__30710\,
            I => data_in_8_2
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__30705\,
            I => data_in_8_2
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__30700\,
            I => \N__30696\
        );

    \I__7213\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30693\
        );

    \I__7212\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30690\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__30693\,
            I => \N__30687\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30681\
        );

    \I__7209\ : Span4Mux_h
    port map (
            O => \N__30687\,
            I => \N__30681\
        );

    \I__7208\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30678\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__30681\,
            I => data_in_14_2
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__30678\,
            I => data_in_14_2
        );

    \I__7205\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30669\
        );

    \I__7204\ : CascadeMux
    port map (
            O => \N__30672\,
            I => \N__30665\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__30669\,
            I => \N__30661\
        );

    \I__7202\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30658\
        );

    \I__7201\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30655\
        );

    \I__7200\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30652\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__30661\,
            I => \N__30649\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N__30645\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30642\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30639\
        );

    \I__7195\ : Span4Mux_h
    port map (
            O => \N__30649\,
            I => \N__30636\
        );

    \I__7194\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30633\
        );

    \I__7193\ : Span12Mux_v
    port map (
            O => \N__30645\,
            I => \N__30626\
        );

    \I__7192\ : Span12Mux_s6_v
    port map (
            O => \N__30642\,
            I => \N__30626\
        );

    \I__7191\ : Span12Mux_s8_h
    port map (
            O => \N__30639\,
            I => \N__30626\
        );

    \I__7190\ : Span4Mux_h
    port map (
            O => \N__30636\,
            I => \N__30623\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__30633\,
            I => \c0.data_in_field_114\
        );

    \I__7188\ : Odrv12
    port map (
            O => \N__30626\,
            I => \c0.data_in_field_114\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__30623\,
            I => \c0.data_in_field_114\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__30616\,
            I => \N__30612\
        );

    \I__7185\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30609\
        );

    \I__7184\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30606\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30603\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__30606\,
            I => \N__30600\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__30603\,
            I => \N__30597\
        );

    \I__7180\ : Span4Mux_v
    port map (
            O => \N__30600\,
            I => \N__30593\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__30597\,
            I => \N__30590\
        );

    \I__7178\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30587\
        );

    \I__7177\ : Odrv4
    port map (
            O => \N__30593\,
            I => data_in_4_2
        );

    \I__7176\ : Odrv4
    port map (
            O => \N__30590\,
            I => data_in_4_2
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__30587\,
            I => data_in_4_2
        );

    \I__7174\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30576\
        );

    \I__7173\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30573\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__30576\,
            I => \N__30567\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30564\
        );

    \I__7170\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30561\
        );

    \I__7169\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30556\
        );

    \I__7168\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30556\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__30567\,
            I => \c0.data_in_field_66\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__30564\,
            I => \c0.data_in_field_66\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__30561\,
            I => \c0.data_in_field_66\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__30556\,
            I => \c0.data_in_field_66\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__30547\,
            I => \N__30543\
        );

    \I__7162\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30540\
        );

    \I__7161\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30537\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30534\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30531\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__30534\,
            I => \N__30526\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__30531\,
            I => \N__30523\
        );

    \I__7156\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30518\
        );

    \I__7155\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30518\
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__30526\,
            I => \c0.data_in_field_84\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__30523\,
            I => \c0.data_in_field_84\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__30518\,
            I => \c0.data_in_field_84\
        );

    \I__7151\ : InMux
    port map (
            O => \N__30511\,
            I => \N__30508\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__30508\,
            I => \N__30505\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__30505\,
            I => \N__30501\
        );

    \I__7148\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30498\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__30501\,
            I => \N__30494\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N__30491\
        );

    \I__7145\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30488\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__30494\,
            I => \c0.n1969\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__30491\,
            I => \c0.n1969\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__30488\,
            I => \c0.n1969\
        );

    \I__7141\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30478\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__30478\,
            I => \N__30475\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__30475\,
            I => \N__30472\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__30472\,
            I => \c0.n25\
        );

    \I__7137\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30463\
        );

    \I__7136\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30463\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__30463\,
            I => \N__30459\
        );

    \I__7134\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30456\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__30459\,
            I => data_in_5_2
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__30456\,
            I => data_in_5_2
        );

    \I__7131\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30445\
        );

    \I__7130\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30442\
        );

    \I__7129\ : CascadeMux
    port map (
            O => \N__30449\,
            I => \N__30439\
        );

    \I__7128\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30436\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__30445\,
            I => \N__30433\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__30442\,
            I => \N__30430\
        );

    \I__7125\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30427\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30424\
        );

    \I__7123\ : Span4Mux_h
    port map (
            O => \N__30433\,
            I => \N__30421\
        );

    \I__7122\ : Span4Mux_v
    port map (
            O => \N__30430\,
            I => \N__30418\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__30427\,
            I => \c0.data_in_field_42\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__30424\,
            I => \c0.data_in_field_42\
        );

    \I__7119\ : Odrv4
    port map (
            O => \N__30421\,
            I => \c0.data_in_field_42\
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__30418\,
            I => \c0.data_in_field_42\
        );

    \I__7117\ : CascadeMux
    port map (
            O => \N__30409\,
            I => \N__30406\
        );

    \I__7116\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30401\
        );

    \I__7115\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30398\
        );

    \I__7114\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30395\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__30401\,
            I => \N__30392\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__30398\,
            I => \N__30389\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__30395\,
            I => \N__30386\
        );

    \I__7110\ : Span4Mux_v
    port map (
            O => \N__30392\,
            I => \N__30383\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__30389\,
            I => \N__30378\
        );

    \I__7108\ : Span4Mux_v
    port map (
            O => \N__30386\,
            I => \N__30375\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__30383\,
            I => \N__30372\
        );

    \I__7106\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30367\
        );

    \I__7105\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30367\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__30378\,
            I => \c0.data_in_field_107\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__30375\,
            I => \c0.data_in_field_107\
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__30372\,
            I => \c0.data_in_field_107\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__30367\,
            I => \c0.data_in_field_107\
        );

    \I__7100\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30355\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__30355\,
            I => \N__30350\
        );

    \I__7098\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30347\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__30353\,
            I => \N__30344\
        );

    \I__7096\ : Sp12to4
    port map (
            O => \N__30350\,
            I => \N__30341\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30338\
        );

    \I__7094\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30334\
        );

    \I__7093\ : Span12Mux_v
    port map (
            O => \N__30341\,
            I => \N__30331\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__30338\,
            I => \N__30328\
        );

    \I__7091\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30325\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__30334\,
            I => \c0.data_in_field_15\
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__30331\,
            I => \c0.data_in_field_15\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__30328\,
            I => \c0.data_in_field_15\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__30325\,
            I => \c0.data_in_field_15\
        );

    \I__7086\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30313\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30310\
        );

    \I__7084\ : Span4Mux_h
    port map (
            O => \N__30310\,
            I => \N__30307\
        );

    \I__7083\ : Span4Mux_h
    port map (
            O => \N__30307\,
            I => \N__30304\
        );

    \I__7082\ : Odrv4
    port map (
            O => \N__30304\,
            I => \c0.n20_adj_1916\
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__30301\,
            I => \N__30298\
        );

    \I__7080\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30294\
        );

    \I__7079\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30291\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30288\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__30291\,
            I => \N__30285\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__30288\,
            I => \N__30279\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__30285\,
            I => \N__30279\
        );

    \I__7074\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30276\
        );

    \I__7073\ : Odrv4
    port map (
            O => \N__30279\,
            I => data_in_8_1
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__30276\,
            I => data_in_8_1
        );

    \I__7071\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30268\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30264\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__30267\,
            I => \N__30261\
        );

    \I__7068\ : Sp12to4
    port map (
            O => \N__30264\,
            I => \N__30254\
        );

    \I__7067\ : InMux
    port map (
            O => \N__30261\,
            I => \N__30251\
        );

    \I__7066\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30248\
        );

    \I__7065\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30243\
        );

    \I__7064\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30243\
        );

    \I__7063\ : InMux
    port map (
            O => \N__30257\,
            I => \N__30240\
        );

    \I__7062\ : Span12Mux_s6_v
    port map (
            O => \N__30254\,
            I => \N__30233\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__30251\,
            I => \N__30233\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__30248\,
            I => \N__30233\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__30243\,
            I => \N__30230\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__30240\,
            I => \c0.data_in_field_65\
        );

    \I__7057\ : Odrv12
    port map (
            O => \N__30233\,
            I => \c0.data_in_field_65\
        );

    \I__7056\ : Odrv4
    port map (
            O => \N__30230\,
            I => \c0.data_in_field_65\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__7054\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30217\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__30217\,
            I => \N__30213\
        );

    \I__7052\ : InMux
    port map (
            O => \N__30216\,
            I => \N__30210\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__30213\,
            I => \N__30207\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__30210\,
            I => \N__30204\
        );

    \I__7049\ : Span4Mux_v
    port map (
            O => \N__30207\,
            I => \N__30200\
        );

    \I__7048\ : Span12Mux_h
    port map (
            O => \N__30204\,
            I => \N__30197\
        );

    \I__7047\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30194\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__30200\,
            I => data_in_16_1
        );

    \I__7045\ : Odrv12
    port map (
            O => \N__30197\,
            I => data_in_16_1
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__30194\,
            I => data_in_16_1
        );

    \I__7043\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30182\
        );

    \I__7042\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30178\
        );

    \I__7041\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30175\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30172\
        );

    \I__7039\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30169\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30164\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__30175\,
            I => \N__30164\
        );

    \I__7036\ : Odrv4
    port map (
            O => \N__30172\,
            I => data_in_2_1
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__30169\,
            I => data_in_2_1
        );

    \I__7034\ : Odrv12
    port map (
            O => \N__30164\,
            I => data_in_2_1
        );

    \I__7033\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30150\
        );

    \I__7031\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30145\
        );

    \I__7030\ : Span4Mux_h
    port map (
            O => \N__30150\,
            I => \N__30142\
        );

    \I__7029\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30137\
        );

    \I__7028\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30137\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__30145\,
            I => \N__30134\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__30142\,
            I => data_in_1_1
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__30137\,
            I => data_in_1_1
        );

    \I__7024\ : Odrv12
    port map (
            O => \N__30134\,
            I => data_in_1_1
        );

    \I__7023\ : CascadeMux
    port map (
            O => \N__30127\,
            I => \N__30124\
        );

    \I__7022\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30120\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__30123\,
            I => \N__30116\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__30120\,
            I => \N__30113\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__30119\,
            I => \N__30110\
        );

    \I__7018\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30107\
        );

    \I__7017\ : Span4Mux_h
    port map (
            O => \N__30113\,
            I => \N__30104\
        );

    \I__7016\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30101\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30097\
        );

    \I__7014\ : Sp12to4
    port map (
            O => \N__30104\,
            I => \N__30092\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__30101\,
            I => \N__30092\
        );

    \I__7012\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30089\
        );

    \I__7011\ : Odrv4
    port map (
            O => \N__30097\,
            I => \c0.data_in_field_48\
        );

    \I__7010\ : Odrv12
    port map (
            O => \N__30092\,
            I => \c0.data_in_field_48\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__30089\,
            I => \c0.data_in_field_48\
        );

    \I__7008\ : CascadeMux
    port map (
            O => \N__30082\,
            I => \N__30079\
        );

    \I__7007\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30076\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__30076\,
            I => \c0.n5701\
        );

    \I__7005\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30069\
        );

    \I__7004\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30066\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__30063\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30060\
        );

    \I__7001\ : Sp12to4
    port map (
            O => \N__30063\,
            I => \N__30057\
        );

    \I__7000\ : Span4Mux_h
    port map (
            O => \N__30060\,
            I => \N__30054\
        );

    \I__6999\ : Span12Mux_s7_v
    port map (
            O => \N__30057\,
            I => \N__30050\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__30054\,
            I => \N__30047\
        );

    \I__6997\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30044\
        );

    \I__6996\ : Odrv12
    port map (
            O => \N__30050\,
            I => data_in_4_4
        );

    \I__6995\ : Odrv4
    port map (
            O => \N__30047\,
            I => data_in_4_4
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__30044\,
            I => data_in_4_4
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__30037\,
            I => \N__30034\
        );

    \I__6992\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__30027\
        );

    \I__6990\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30024\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__30027\,
            I => \N__30021\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30018\
        );

    \I__6987\ : Span4Mux_h
    port map (
            O => \N__30021\,
            I => \N__30013\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__30018\,
            I => \N__30013\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__30013\,
            I => \N__30009\
        );

    \I__6984\ : InMux
    port map (
            O => \N__30012\,
            I => \N__30006\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__30009\,
            I => data_in_6_4
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__30006\,
            I => data_in_6_4
        );

    \I__6981\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29998\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__29998\,
            I => \N__29995\
        );

    \I__6979\ : Span4Mux_h
    port map (
            O => \N__29995\,
            I => \N__29990\
        );

    \I__6978\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29987\
        );

    \I__6977\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29984\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__29990\,
            I => data_in_7_2
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__29987\,
            I => data_in_7_2
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__29984\,
            I => data_in_7_2
        );

    \I__6973\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29974\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__29974\,
            I => \N__29971\
        );

    \I__6971\ : Span4Mux_v
    port map (
            O => \N__29971\,
            I => \N__29967\
        );

    \I__6970\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29964\
        );

    \I__6969\ : Sp12to4
    port map (
            O => \N__29967\,
            I => \N__29961\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__29964\,
            I => \N__29958\
        );

    \I__6967\ : Span12Mux_s10_h
    port map (
            O => \N__29961\,
            I => \N__29954\
        );

    \I__6966\ : Span4Mux_h
    port map (
            O => \N__29958\,
            I => \N__29951\
        );

    \I__6965\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29948\
        );

    \I__6964\ : Odrv12
    port map (
            O => \N__29954\,
            I => data_in_10_6
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__29951\,
            I => data_in_10_6
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__29948\,
            I => data_in_10_6
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__29941\,
            I => \N__29938\
        );

    \I__6960\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29935\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__29935\,
            I => \N__29932\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__29932\,
            I => \N__29929\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__29929\,
            I => \N__29924\
        );

    \I__6956\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29921\
        );

    \I__6955\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29918\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__29924\,
            I => data_in_9_6
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__29921\,
            I => data_in_9_6
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__29918\,
            I => data_in_9_6
        );

    \I__6951\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29907\
        );

    \I__6950\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29903\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__29907\,
            I => \N__29900\
        );

    \I__6948\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29897\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__29903\,
            I => data_in_10_0
        );

    \I__6946\ : Odrv12
    port map (
            O => \N__29900\,
            I => data_in_10_0
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__29897\,
            I => data_in_10_0
        );

    \I__6944\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29886\
        );

    \I__6943\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29882\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__29886\,
            I => \N__29879\
        );

    \I__6941\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29876\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__29882\,
            I => \N__29870\
        );

    \I__6939\ : Span4Mux_v
    port map (
            O => \N__29879\,
            I => \N__29870\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29867\
        );

    \I__6937\ : CascadeMux
    port map (
            O => \N__29875\,
            I => \N__29864\
        );

    \I__6936\ : Span4Mux_h
    port map (
            O => \N__29870\,
            I => \N__29861\
        );

    \I__6935\ : Span4Mux_h
    port map (
            O => \N__29867\,
            I => \N__29858\
        );

    \I__6934\ : InMux
    port map (
            O => \N__29864\,
            I => \N__29854\
        );

    \I__6933\ : Span4Mux_h
    port map (
            O => \N__29861\,
            I => \N__29849\
        );

    \I__6932\ : Span4Mux_h
    port map (
            O => \N__29858\,
            I => \N__29849\
        );

    \I__6931\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29846\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__29854\,
            I => \c0.data_in_field_80\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__29849\,
            I => \c0.data_in_field_80\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__29846\,
            I => \c0.data_in_field_80\
        );

    \I__6927\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29834\
        );

    \I__6926\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29829\
        );

    \I__6925\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29829\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__29834\,
            I => data_in_13_6
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__29829\,
            I => data_in_13_6
        );

    \I__6922\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29821\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__29821\,
            I => n5332
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__29818\,
            I => \n5331_cascade_\
        );

    \I__6919\ : IoInMux
    port map (
            O => \N__29815\,
            I => \N__29812\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__29812\,
            I => \N__29809\
        );

    \I__6917\ : IoSpan4Mux
    port map (
            O => \N__29809\,
            I => \N__29806\
        );

    \I__6916\ : IoSpan4Mux
    port map (
            O => \N__29806\,
            I => \N__29803\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__29803\,
            I => \LED_c\
        );

    \I__6914\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29796\
        );

    \I__6913\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29791\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29787\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__29795\,
            I => \N__29783\
        );

    \I__6910\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29780\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__29791\,
            I => \N__29777\
        );

    \I__6908\ : InMux
    port map (
            O => \N__29790\,
            I => \N__29774\
        );

    \I__6907\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29771\
        );

    \I__6906\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29768\
        );

    \I__6905\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29765\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__29780\,
            I => \N__29762\
        );

    \I__6903\ : Span4Mux_h
    port map (
            O => \N__29777\,
            I => \N__29757\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29757\
        );

    \I__6901\ : Span4Mux_h
    port map (
            O => \N__29771\,
            I => \N__29752\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29752\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__29765\,
            I => \c0.data_in_field_97\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__29762\,
            I => \c0.data_in_field_97\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__29757\,
            I => \c0.data_in_field_97\
        );

    \I__6896\ : Odrv4
    port map (
            O => \N__29752\,
            I => \c0.data_in_field_97\
        );

    \I__6895\ : CascadeMux
    port map (
            O => \N__29743\,
            I => \N__29740\
        );

    \I__6894\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29736\
        );

    \I__6893\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29733\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__29736\,
            I => \N__29730\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__29733\,
            I => \N__29727\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__29730\,
            I => \N__29724\
        );

    \I__6889\ : Span12Mux_v
    port map (
            O => \N__29727\,
            I => \N__29721\
        );

    \I__6888\ : Span4Mux_h
    port map (
            O => \N__29724\,
            I => \N__29718\
        );

    \I__6887\ : Odrv12
    port map (
            O => \N__29721\,
            I => \c0.n1972\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__29718\,
            I => \c0.n1972\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__29713\,
            I => \N__29710\
        );

    \I__6884\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29707\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29704\
        );

    \I__6882\ : Span4Mux_v
    port map (
            O => \N__29704\,
            I => \N__29699\
        );

    \I__6881\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29696\
        );

    \I__6880\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29693\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__29699\,
            I => data_in_9_4
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__29696\,
            I => data_in_9_4
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__29693\,
            I => data_in_9_4
        );

    \I__6876\ : InMux
    port map (
            O => \N__29686\,
            I => \N__29683\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__29683\,
            I => \N__29680\
        );

    \I__6874\ : Span4Mux_v
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__6873\ : Span4Mux_h
    port map (
            O => \N__29677\,
            I => \N__29671\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29666\
        );

    \I__6871\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29666\
        );

    \I__6870\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29663\
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__29671\,
            I => \c0.data_in_field_76\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__29666\,
            I => \c0.data_in_field_76\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__29663\,
            I => \c0.data_in_field_76\
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__29656\,
            I => \N__29652\
        );

    \I__6865\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29649\
        );

    \I__6864\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29646\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__29649\,
            I => \N__29640\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__29646\,
            I => \N__29640\
        );

    \I__6861\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29637\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__29640\,
            I => \N__29634\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__29637\,
            I => data_in_0_1
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__29634\,
            I => data_in_0_1
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__29629\,
            I => \N__29626\
        );

    \I__6856\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29621\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29618\
        );

    \I__6854\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29615\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__29621\,
            I => data_in_5_5
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__29618\,
            I => data_in_5_5
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__29615\,
            I => data_in_5_5
        );

    \I__6850\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29604\
        );

    \I__6849\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29601\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__29604\,
            I => \N__29598\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__29601\,
            I => \N__29594\
        );

    \I__6846\ : Span4Mux_h
    port map (
            O => \N__29598\,
            I => \N__29591\
        );

    \I__6845\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29587\
        );

    \I__6844\ : Span4Mux_h
    port map (
            O => \N__29594\,
            I => \N__29584\
        );

    \I__6843\ : Span4Mux_h
    port map (
            O => \N__29591\,
            I => \N__29581\
        );

    \I__6842\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29578\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__29587\,
            I => \c0.data_in_field_45\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__29584\,
            I => \c0.data_in_field_45\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__29581\,
            I => \c0.data_in_field_45\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__29578\,
            I => \c0.data_in_field_45\
        );

    \I__6837\ : CascadeMux
    port map (
            O => \N__29569\,
            I => \N__29566\
        );

    \I__6836\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29563\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__29563\,
            I => \N__29559\
        );

    \I__6834\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29556\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__29559\,
            I => \N__29551\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29551\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__29551\,
            I => \N__29547\
        );

    \I__6830\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29544\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__29547\,
            I => data_in_9_0
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__29544\,
            I => data_in_9_0
        );

    \I__6827\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29536\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__29536\,
            I => \N__29531\
        );

    \I__6825\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29528\
        );

    \I__6824\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29524\
        );

    \I__6823\ : Span4Mux_v
    port map (
            O => \N__29531\,
            I => \N__29519\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__29528\,
            I => \N__29519\
        );

    \I__6821\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29516\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29512\
        );

    \I__6819\ : Span4Mux_h
    port map (
            O => \N__29519\,
            I => \N__29509\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29506\
        );

    \I__6817\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29503\
        );

    \I__6816\ : Span12Mux_s9_h
    port map (
            O => \N__29512\,
            I => \N__29500\
        );

    \I__6815\ : Span4Mux_h
    port map (
            O => \N__29509\,
            I => \N__29495\
        );

    \I__6814\ : Span4Mux_h
    port map (
            O => \N__29506\,
            I => \N__29495\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__29503\,
            I => \c0.data_in_field_128\
        );

    \I__6812\ : Odrv12
    port map (
            O => \N__29500\,
            I => \c0.data_in_field_128\
        );

    \I__6811\ : Odrv4
    port map (
            O => \N__29495\,
            I => \c0.data_in_field_128\
        );

    \I__6810\ : CascadeMux
    port map (
            O => \N__29488\,
            I => \N__29485\
        );

    \I__6809\ : InMux
    port map (
            O => \N__29485\,
            I => \N__29480\
        );

    \I__6808\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29475\
        );

    \I__6807\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29475\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__29480\,
            I => \N__29472\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__29475\,
            I => \c0.data_in_field_16\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__29472\,
            I => \c0.data_in_field_16\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__29467\,
            I => \N__29464\
        );

    \I__6802\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29461\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__29461\,
            I => \N__29458\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__29458\,
            I => \N__29452\
        );

    \I__6799\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29447\
        );

    \I__6798\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29447\
        );

    \I__6797\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29444\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__29452\,
            I => \c0.data_in_field_72\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__29447\,
            I => \c0.data_in_field_72\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__29444\,
            I => \c0.data_in_field_72\
        );

    \I__6793\ : InMux
    port map (
            O => \N__29437\,
            I => \N__29433\
        );

    \I__6792\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29430\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__29433\,
            I => \c0.n5188\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__29430\,
            I => \c0.n5188\
        );

    \I__6789\ : CascadeMux
    port map (
            O => \N__29425\,
            I => \c0.n5138_cascade_\
        );

    \I__6788\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29419\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__29419\,
            I => \N__29416\
        );

    \I__6786\ : Odrv12
    port map (
            O => \N__29416\,
            I => \c0.n15_adj_1968\
        );

    \I__6785\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29409\
        );

    \I__6784\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29406\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29403\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__29406\,
            I => \N__29400\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__29403\,
            I => \N__29393\
        );

    \I__6780\ : Span4Mux_h
    port map (
            O => \N__29400\,
            I => \N__29393\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__29399\,
            I => \N__29390\
        );

    \I__6778\ : InMux
    port map (
            O => \N__29398\,
            I => \N__29387\
        );

    \I__6777\ : Span4Mux_v
    port map (
            O => \N__29393\,
            I => \N__29384\
        );

    \I__6776\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29381\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__29387\,
            I => data_in_3_2
        );

    \I__6774\ : Odrv4
    port map (
            O => \N__29384\,
            I => data_in_3_2
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__29381\,
            I => data_in_3_2
        );

    \I__6772\ : InMux
    port map (
            O => \N__29374\,
            I => \N__29371\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__6770\ : Span4Mux_h
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__6769\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29356\
        );

    \I__6768\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29356\
        );

    \I__6767\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29353\
        );

    \I__6766\ : Span4Mux_v
    port map (
            O => \N__29362\,
            I => \N__29350\
        );

    \I__6765\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29347\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__29356\,
            I => \N__29344\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__29353\,
            I => \c0.data_in_field_26\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__29350\,
            I => \c0.data_in_field_26\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__29347\,
            I => \c0.data_in_field_26\
        );

    \I__6760\ : Odrv12
    port map (
            O => \N__29344\,
            I => \c0.data_in_field_26\
        );

    \I__6759\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29331\
        );

    \I__6758\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29328\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__29331\,
            I => \N__29325\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__29328\,
            I => \N__29321\
        );

    \I__6755\ : Span4Mux_s3_v
    port map (
            O => \N__29325\,
            I => \N__29318\
        );

    \I__6754\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29315\
        );

    \I__6753\ : Span12Mux_h
    port map (
            O => \N__29321\,
            I => \N__29312\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__29318\,
            I => \N__29309\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__29315\,
            I => data_in_4_1
        );

    \I__6750\ : Odrv12
    port map (
            O => \N__29312\,
            I => data_in_4_1
        );

    \I__6749\ : Odrv4
    port map (
            O => \N__29309\,
            I => data_in_4_1
        );

    \I__6748\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29299\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__29299\,
            I => \N__29295\
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__29298\,
            I => \N__29291\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__29295\,
            I => \N__29288\
        );

    \I__6744\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29285\
        );

    \I__6743\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29281\
        );

    \I__6742\ : Span4Mux_h
    port map (
            O => \N__29288\,
            I => \N__29276\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29276\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__29284\,
            I => \N__29273\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__29281\,
            I => \N__29270\
        );

    \I__6738\ : Span4Mux_h
    port map (
            O => \N__29276\,
            I => \N__29267\
        );

    \I__6737\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29264\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__29270\,
            I => \c0.data_in_field_33\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__29267\,
            I => \c0.data_in_field_33\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__29264\,
            I => \c0.data_in_field_33\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__6732\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29251\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29247\
        );

    \I__6730\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29243\
        );

    \I__6729\ : Span4Mux_h
    port map (
            O => \N__29247\,
            I => \N__29240\
        );

    \I__6728\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29236\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__29243\,
            I => \N__29233\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__29240\,
            I => \N__29230\
        );

    \I__6725\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29227\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__29236\,
            I => data_in_2_2
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__29233\,
            I => data_in_2_2
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__29230\,
            I => data_in_2_2
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__29227\,
            I => data_in_2_2
        );

    \I__6720\ : CascadeMux
    port map (
            O => \N__29218\,
            I => \N__29214\
        );

    \I__6719\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29211\
        );

    \I__6718\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__29211\,
            I => \N__29205\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29202\
        );

    \I__6715\ : Span4Mux_h
    port map (
            O => \N__29205\,
            I => \N__29199\
        );

    \I__6714\ : Span4Mux_h
    port map (
            O => \N__29202\,
            I => \N__29196\
        );

    \I__6713\ : Span4Mux_v
    port map (
            O => \N__29199\,
            I => \N__29191\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__29196\,
            I => \N__29188\
        );

    \I__6711\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29183\
        );

    \I__6710\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29183\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__29191\,
            I => \c0.data_in_field_18\
        );

    \I__6708\ : Odrv4
    port map (
            O => \N__29188\,
            I => \c0.data_in_field_18\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__29183\,
            I => \c0.data_in_field_18\
        );

    \I__6706\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29173\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__29173\,
            I => \c0.n6\
        );

    \I__6704\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29166\
        );

    \I__6703\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29163\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__29166\,
            I => \N__29160\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29157\
        );

    \I__6700\ : Span4Mux_v
    port map (
            O => \N__29160\,
            I => \N__29152\
        );

    \I__6699\ : Span4Mux_v
    port map (
            O => \N__29157\,
            I => \N__29152\
        );

    \I__6698\ : Sp12to4
    port map (
            O => \N__29152\,
            I => \N__29148\
        );

    \I__6697\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29145\
        );

    \I__6696\ : Odrv12
    port map (
            O => \N__29148\,
            I => data_in_4_0
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__29145\,
            I => data_in_4_0
        );

    \I__6694\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29136\
        );

    \I__6693\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29133\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29130\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29126\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__29130\,
            I => \N__29123\
        );

    \I__6689\ : InMux
    port map (
            O => \N__29129\,
            I => \N__29120\
        );

    \I__6688\ : Span4Mux_v
    port map (
            O => \N__29126\,
            I => \N__29115\
        );

    \I__6687\ : Span4Mux_v
    port map (
            O => \N__29123\,
            I => \N__29115\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__29120\,
            I => \N__29110\
        );

    \I__6685\ : Span4Mux_h
    port map (
            O => \N__29115\,
            I => \N__29107\
        );

    \I__6684\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29102\
        );

    \I__6683\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29102\
        );

    \I__6682\ : Odrv12
    port map (
            O => \N__29110\,
            I => \c0.data_in_field_32\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__29107\,
            I => \c0.data_in_field_32\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__29102\,
            I => \c0.data_in_field_32\
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__29095\,
            I => \N__29092\
        );

    \I__6678\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29088\
        );

    \I__6677\ : InMux
    port map (
            O => \N__29091\,
            I => \N__29085\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29082\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__29085\,
            I => \N__29079\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__29082\,
            I => \N__29073\
        );

    \I__6673\ : Span4Mux_h
    port map (
            O => \N__29079\,
            I => \N__29073\
        );

    \I__6672\ : InMux
    port map (
            O => \N__29078\,
            I => \N__29070\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__29073\,
            I => data_in_13_2
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__29070\,
            I => data_in_13_2
        );

    \I__6669\ : CascadeMux
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__6668\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29059\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__29059\,
            I => \N__29056\
        );

    \I__6666\ : Span4Mux_h
    port map (
            O => \N__29056\,
            I => \N__29052\
        );

    \I__6665\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29049\
        );

    \I__6664\ : Span4Mux_v
    port map (
            O => \N__29052\,
            I => \N__29044\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29044\
        );

    \I__6662\ : Span4Mux_h
    port map (
            O => \N__29044\,
            I => \N__29040\
        );

    \I__6661\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29037\
        );

    \I__6660\ : Odrv4
    port map (
            O => \N__29040\,
            I => data_in_12_2
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__29037\,
            I => data_in_12_2
        );

    \I__6658\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29026\
        );

    \I__6657\ : InMux
    port map (
            O => \N__29031\,
            I => \N__29023\
        );

    \I__6656\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29020\
        );

    \I__6655\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29016\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__29026\,
            I => \N__29012\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__29023\,
            I => \N__29009\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__29020\,
            I => \N__29006\
        );

    \I__6651\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29003\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29000\
        );

    \I__6649\ : InMux
    port map (
            O => \N__29015\,
            I => \N__28997\
        );

    \I__6648\ : Span4Mux_h
    port map (
            O => \N__29012\,
            I => \N__28994\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__29009\,
            I => \N__28991\
        );

    \I__6646\ : Span12Mux_v
    port map (
            O => \N__29006\,
            I => \N__28984\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__29003\,
            I => \N__28984\
        );

    \I__6644\ : Sp12to4
    port map (
            O => \N__29000\,
            I => \N__28984\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__28997\,
            I => \c0.data_in_field_64\
        );

    \I__6642\ : Odrv4
    port map (
            O => \N__28994\,
            I => \c0.data_in_field_64\
        );

    \I__6641\ : Odrv4
    port map (
            O => \N__28991\,
            I => \c0.data_in_field_64\
        );

    \I__6640\ : Odrv12
    port map (
            O => \N__28984\,
            I => \c0.data_in_field_64\
        );

    \I__6639\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28970\
        );

    \I__6638\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28965\
        );

    \I__6637\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28965\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__28970\,
            I => \c0.n5179\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__28965\,
            I => \c0.n5179\
        );

    \I__6634\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28956\
        );

    \I__6633\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28951\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28948\
        );

    \I__6631\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28945\
        );

    \I__6630\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28942\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28939\
        );

    \I__6628\ : Span4Mux_h
    port map (
            O => \N__28948\,
            I => \N__28936\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28933\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__28942\,
            I => \c0.data_in_field_46\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__28939\,
            I => \c0.data_in_field_46\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__28936\,
            I => \c0.data_in_field_46\
        );

    \I__6623\ : Odrv4
    port map (
            O => \N__28933\,
            I => \c0.data_in_field_46\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__28924\,
            I => \N__28921\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28918\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__28918\,
            I => \N__28911\
        );

    \I__6619\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28908\
        );

    \I__6618\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28905\
        );

    \I__6617\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28902\
        );

    \I__6616\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28899\
        );

    \I__6615\ : Span12Mux_s6_v
    port map (
            O => \N__28911\,
            I => \N__28896\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__28908\,
            I => \c0.data_in_field_4\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__28905\,
            I => \c0.data_in_field_4\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28902\,
            I => \c0.data_in_field_4\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__28899\,
            I => \c0.data_in_field_4\
        );

    \I__6610\ : Odrv12
    port map (
            O => \N__28896\,
            I => \c0.data_in_field_4\
        );

    \I__6609\ : CascadeMux
    port map (
            O => \N__28885\,
            I => \c0.n1767_cascade_\
        );

    \I__6608\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28879\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__28879\,
            I => \N__28875\
        );

    \I__6606\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28872\
        );

    \I__6605\ : Odrv4
    port map (
            O => \N__28875\,
            I => \c0.n1899\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__28872\,
            I => \c0.n1899\
        );

    \I__6603\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28864\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__28864\,
            I => \c0.n5126\
        );

    \I__6601\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__28855\,
            I => \N__28850\
        );

    \I__6598\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28845\
        );

    \I__6597\ : InMux
    port map (
            O => \N__28853\,
            I => \N__28841\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__28850\,
            I => \N__28838\
        );

    \I__6595\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28835\
        );

    \I__6594\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28832\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__28845\,
            I => \N__28829\
        );

    \I__6592\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28826\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__28841\,
            I => \c0.data_in_field_140\
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__28838\,
            I => \c0.data_in_field_140\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__28835\,
            I => \c0.data_in_field_140\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__28832\,
            I => \c0.data_in_field_140\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__28829\,
            I => \c0.data_in_field_140\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__28826\,
            I => \c0.data_in_field_140\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__28813\,
            I => \c0.n5126_cascade_\
        );

    \I__6584\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28805\
        );

    \I__6583\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28802\
        );

    \I__6582\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28799\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__28805\,
            I => \N__28796\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28793\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__28799\,
            I => \N__28790\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__28796\,
            I => \N__28783\
        );

    \I__6577\ : Span4Mux_v
    port map (
            O => \N__28793\,
            I => \N__28783\
        );

    \I__6576\ : Span4Mux_h
    port map (
            O => \N__28790\,
            I => \N__28780\
        );

    \I__6575\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28777\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__28788\,
            I => \N__28774\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__28783\,
            I => \N__28769\
        );

    \I__6572\ : Span4Mux_v
    port map (
            O => \N__28780\,
            I => \N__28769\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28766\
        );

    \I__6570\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28763\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__28769\,
            I => \c0.data_in_field_125\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__28766\,
            I => \c0.data_in_field_125\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__28763\,
            I => \c0.data_in_field_125\
        );

    \I__6566\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28753\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__6564\ : Span4Mux_h
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__28744\,
            I => \c0.n20_adj_1899\
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__28741\,
            I => \N__28738\
        );

    \I__6560\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28734\
        );

    \I__6559\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28731\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__28734\,
            I => \N__28726\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__28731\,
            I => \N__28726\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__28726\,
            I => \N__28722\
        );

    \I__6555\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28719\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__28722\,
            I => data_in_14_6
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__28719\,
            I => data_in_14_6
        );

    \I__6552\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28711\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__28711\,
            I => \c0.n10_adj_1872\
        );

    \I__6550\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28704\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__28707\,
            I => \N__28701\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__28704\,
            I => \N__28698\
        );

    \I__6547\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28695\
        );

    \I__6546\ : Span4Mux_h
    port map (
            O => \N__28698\,
            I => \N__28692\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__28695\,
            I => \N__28689\
        );

    \I__6544\ : Span4Mux_v
    port map (
            O => \N__28692\,
            I => \N__28686\
        );

    \I__6543\ : Span4Mux_h
    port map (
            O => \N__28689\,
            I => \N__28682\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__28686\,
            I => \N__28679\
        );

    \I__6541\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28676\
        );

    \I__6540\ : Odrv4
    port map (
            O => \N__28682\,
            I => data_in_12_4
        );

    \I__6539\ : Odrv4
    port map (
            O => \N__28679\,
            I => data_in_12_4
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__28676\,
            I => data_in_12_4
        );

    \I__6537\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28666\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28662\
        );

    \I__6535\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28659\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__28662\,
            I => \N__28656\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__28659\,
            I => \N__28651\
        );

    \I__6532\ : Span4Mux_h
    port map (
            O => \N__28656\,
            I => \N__28648\
        );

    \I__6531\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28643\
        );

    \I__6530\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28643\
        );

    \I__6529\ : Odrv4
    port map (
            O => \N__28651\,
            I => \c0.data_in_field_100\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__28648\,
            I => \c0.data_in_field_100\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__28643\,
            I => \c0.data_in_field_100\
        );

    \I__6526\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28632\
        );

    \I__6525\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28627\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__28632\,
            I => \N__28624\
        );

    \I__6523\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28621\
        );

    \I__6522\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28618\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__28627\,
            I => \c0.data_in_field_40\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__28624\,
            I => \c0.data_in_field_40\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__28621\,
            I => \c0.data_in_field_40\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__28618\,
            I => \c0.data_in_field_40\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__28609\,
            I => \N__28605\
        );

    \I__6516\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28602\
        );

    \I__6515\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28599\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__28602\,
            I => \N__28596\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28593\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__28596\,
            I => \N__28590\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__28593\,
            I => \N__28586\
        );

    \I__6510\ : Span4Mux_h
    port map (
            O => \N__28590\,
            I => \N__28583\
        );

    \I__6509\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28580\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__28586\,
            I => data_in_11_1
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__28583\,
            I => data_in_11_1
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__28580\,
            I => data_in_11_1
        );

    \I__6505\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28570\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__28570\,
            I => \N__28567\
        );

    \I__6503\ : Span4Mux_h
    port map (
            O => \N__28567\,
            I => \N__28564\
        );

    \I__6502\ : Span4Mux_h
    port map (
            O => \N__28564\,
            I => \N__28559\
        );

    \I__6501\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28556\
        );

    \I__6500\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28553\
        );

    \I__6499\ : Span4Mux_v
    port map (
            O => \N__28559\,
            I => \N__28550\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__28556\,
            I => data_in_10_1
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__28553\,
            I => data_in_10_1
        );

    \I__6496\ : Odrv4
    port map (
            O => \N__28550\,
            I => data_in_10_1
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__28543\,
            I => \N__28540\
        );

    \I__6494\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__28537\,
            I => \N__28533\
        );

    \I__6492\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28530\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__28533\,
            I => \N__28527\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__28530\,
            I => \N__28524\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__28527\,
            I => \N__28518\
        );

    \I__6488\ : Span4Mux_h
    port map (
            O => \N__28524\,
            I => \N__28518\
        );

    \I__6487\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28515\
        );

    \I__6486\ : Odrv4
    port map (
            O => \N__28518\,
            I => data_in_11_0
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__28515\,
            I => data_in_11_0
        );

    \I__6484\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28506\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__28509\,
            I => \N__28502\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__28506\,
            I => \N__28499\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__28505\,
            I => \N__28496\
        );

    \I__6480\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28493\
        );

    \I__6479\ : Span4Mux_h
    port map (
            O => \N__28499\,
            I => \N__28490\
        );

    \I__6478\ : InMux
    port map (
            O => \N__28496\,
            I => \N__28487\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__28493\,
            I => \c0.data_in_field_14\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__28490\,
            I => \c0.data_in_field_14\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__28487\,
            I => \c0.data_in_field_14\
        );

    \I__6474\ : CascadeMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__6473\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__6471\ : Span4Mux_h
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__6470\ : Span4Mux_h
    port map (
            O => \N__28468\,
            I => \N__28465\
        );

    \I__6469\ : Odrv4
    port map (
            O => \N__28465\,
            I => \c0.n5911\
        );

    \I__6468\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28459\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28453\
        );

    \I__6466\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28448\
        );

    \I__6465\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28448\
        );

    \I__6464\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28445\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__28453\,
            I => \c0.data_in_field_6\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__28448\,
            I => \c0.data_in_field_6\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__28445\,
            I => \c0.data_in_field_6\
        );

    \I__6460\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28434\
        );

    \I__6459\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28431\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28428\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__28431\,
            I => \N__28425\
        );

    \I__6456\ : Span4Mux_v
    port map (
            O => \N__28428\,
            I => \N__28419\
        );

    \I__6455\ : Span4Mux_s3_h
    port map (
            O => \N__28425\,
            I => \N__28419\
        );

    \I__6454\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28416\
        );

    \I__6453\ : Span4Mux_h
    port map (
            O => \N__28419\,
            I => \N__28411\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__28416\,
            I => \N__28411\
        );

    \I__6451\ : Span4Mux_h
    port map (
            O => \N__28411\,
            I => \N__28406\
        );

    \I__6450\ : InMux
    port map (
            O => \N__28410\,
            I => \N__28401\
        );

    \I__6449\ : InMux
    port map (
            O => \N__28409\,
            I => \N__28401\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__28406\,
            I => \c0.data_in_field_138\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__28401\,
            I => \c0.data_in_field_138\
        );

    \I__6446\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28392\
        );

    \I__6445\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28389\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__28392\,
            I => \N__28386\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28383\
        );

    \I__6442\ : Span4Mux_s3_h
    port map (
            O => \N__28386\,
            I => \N__28377\
        );

    \I__6441\ : Span4Mux_v
    port map (
            O => \N__28383\,
            I => \N__28377\
        );

    \I__6440\ : CascadeMux
    port map (
            O => \N__28382\,
            I => \N__28374\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__28377\,
            I => \N__28371\
        );

    \I__6438\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28368\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__28371\,
            I => \N__28361\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28361\
        );

    \I__6435\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28356\
        );

    \I__6434\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28356\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__28361\,
            I => \c0.data_in_field_130\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__28356\,
            I => \c0.data_in_field_130\
        );

    \I__6431\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28348\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__28348\,
            I => \N__28345\
        );

    \I__6429\ : Span4Mux_h
    port map (
            O => \N__28345\,
            I => \N__28342\
        );

    \I__6428\ : Span4Mux_h
    port map (
            O => \N__28342\,
            I => \N__28339\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__28339\,
            I => \c0.n5123\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__28336\,
            I => \c0.n5123_cascade_\
        );

    \I__6425\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__28330\,
            I => \N__28327\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__28327\,
            I => \N__28323\
        );

    \I__6422\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28320\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__28323\,
            I => \N__28317\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__28320\,
            I => \N__28314\
        );

    \I__6419\ : Span4Mux_h
    port map (
            O => \N__28317\,
            I => \N__28311\
        );

    \I__6418\ : Odrv12
    port map (
            O => \N__28314\,
            I => \c0.n5231\
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__28311\,
            I => \c0.n5231\
        );

    \I__6416\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28301\
        );

    \I__6415\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28298\
        );

    \I__6414\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28295\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__28301\,
            I => \N__28291\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28288\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28285\
        );

    \I__6410\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28281\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__28291\,
            I => \N__28278\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__28288\,
            I => \N__28273\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__28285\,
            I => \N__28273\
        );

    \I__6406\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28270\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__28281\,
            I => \c0.data_in_field_58\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__28278\,
            I => \c0.data_in_field_58\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__28273\,
            I => \c0.data_in_field_58\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__28270\,
            I => \c0.data_in_field_58\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__28261\,
            I => \c0.n5773_cascade_\
        );

    \I__6400\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28254\
        );

    \I__6399\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28251\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__28254\,
            I => \N__28246\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28243\
        );

    \I__6396\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28240\
        );

    \I__6395\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28237\
        );

    \I__6394\ : Span4Mux_v
    port map (
            O => \N__28246\,
            I => \N__28234\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__28243\,
            I => \N__28231\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28228\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__28237\,
            I => \c0.data_in_field_34\
        );

    \I__6390\ : Odrv4
    port map (
            O => \N__28234\,
            I => \c0.data_in_field_34\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__28231\,
            I => \c0.data_in_field_34\
        );

    \I__6388\ : Odrv12
    port map (
            O => \N__28228\,
            I => \c0.data_in_field_34\
        );

    \I__6387\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28216\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__6385\ : Span4Mux_h
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__6384\ : Odrv4
    port map (
            O => \N__28210\,
            I => \c0.n5441\
        );

    \I__6383\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28201\
        );

    \I__6381\ : Span12Mux_v
    port map (
            O => \N__28201\,
            I => \N__28198\
        );

    \I__6380\ : Odrv12
    port map (
            O => \N__28198\,
            I => \c0.n5477\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__28195\,
            I => \N__28192\
        );

    \I__6378\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28189\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__28189\,
            I => \N__28185\
        );

    \I__6376\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28182\
        );

    \I__6375\ : Span4Mux_h
    port map (
            O => \N__28185\,
            I => \N__28179\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__28182\,
            I => \N__28173\
        );

    \I__6373\ : Span4Mux_h
    port map (
            O => \N__28179\,
            I => \N__28173\
        );

    \I__6372\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28170\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__28173\,
            I => \N__28167\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__28170\,
            I => data_in_16_4
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__28167\,
            I => data_in_16_4
        );

    \I__6368\ : CascadeMux
    port map (
            O => \N__28162\,
            I => \N__28159\
        );

    \I__6367\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28156\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__28156\,
            I => \N__28152\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__28155\,
            I => \N__28149\
        );

    \I__6364\ : Span4Mux_h
    port map (
            O => \N__28152\,
            I => \N__28145\
        );

    \I__6363\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28140\
        );

    \I__6362\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28140\
        );

    \I__6361\ : Span4Mux_h
    port map (
            O => \N__28145\,
            I => \N__28137\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__28140\,
            I => data_in_15_4
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__28137\,
            I => data_in_15_4
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__28132\,
            I => \N__28127\
        );

    \I__6357\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28124\
        );

    \I__6356\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28121\
        );

    \I__6355\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28118\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__28124\,
            I => \N__28115\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__28121\,
            I => data_in_8_6
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__28118\,
            I => data_in_8_6
        );

    \I__6351\ : Odrv4
    port map (
            O => \N__28115\,
            I => data_in_8_6
        );

    \I__6350\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28104\
        );

    \I__6349\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28101\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__28104\,
            I => \N__28097\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__28101\,
            I => \N__28094\
        );

    \I__6346\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28091\
        );

    \I__6345\ : Span4Mux_h
    port map (
            O => \N__28097\,
            I => \N__28088\
        );

    \I__6344\ : Span4Mux_h
    port map (
            O => \N__28094\,
            I => \N__28085\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__28091\,
            I => data_in_6_5
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__28088\,
            I => data_in_6_5
        );

    \I__6341\ : Odrv4
    port map (
            O => \N__28085\,
            I => data_in_6_5
        );

    \I__6340\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28075\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__28075\,
            I => \N__28070\
        );

    \I__6338\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28067\
        );

    \I__6337\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28064\
        );

    \I__6336\ : Odrv4
    port map (
            O => \N__28070\,
            I => data_in_4_6
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__28067\,
            I => data_in_4_6
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__28064\,
            I => data_in_4_6
        );

    \I__6333\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28054\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__28054\,
            I => \N__28051\
        );

    \I__6331\ : Span4Mux_h
    port map (
            O => \N__28051\,
            I => \N__28047\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__28050\,
            I => \N__28043\
        );

    \I__6329\ : Sp12to4
    port map (
            O => \N__28047\,
            I => \N__28040\
        );

    \I__6328\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28035\
        );

    \I__6327\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28035\
        );

    \I__6326\ : Odrv12
    port map (
            O => \N__28040\,
            I => data_in_6_0
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__28035\,
            I => data_in_6_0
        );

    \I__6324\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28026\
        );

    \I__6323\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28021\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28018\
        );

    \I__6321\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28015\
        );

    \I__6320\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28012\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__28021\,
            I => \N__28009\
        );

    \I__6318\ : Span4Mux_v
    port map (
            O => \N__28018\,
            I => \N__28004\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__28015\,
            I => \N__28004\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__28012\,
            I => \N__28000\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__28009\,
            I => \N__27995\
        );

    \I__6314\ : Span4Mux_h
    port map (
            O => \N__28004\,
            I => \N__27995\
        );

    \I__6313\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27991\
        );

    \I__6312\ : Span12Mux_v
    port map (
            O => \N__28000\,
            I => \N__27988\
        );

    \I__6311\ : Span4Mux_h
    port map (
            O => \N__27995\,
            I => \N__27985\
        );

    \I__6310\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27982\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__27991\,
            I => \c0.data_in_field_60\
        );

    \I__6308\ : Odrv12
    port map (
            O => \N__27988\,
            I => \c0.data_in_field_60\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__27985\,
            I => \c0.data_in_field_60\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__27982\,
            I => \c0.data_in_field_60\
        );

    \I__6305\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27970\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__27970\,
            I => \c0.n6_adj_1875\
        );

    \I__6303\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27963\
        );

    \I__6302\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27960\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__27963\,
            I => \N__27957\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__27960\,
            I => \N__27953\
        );

    \I__6299\ : Span4Mux_s2_v
    port map (
            O => \N__27957\,
            I => \N__27950\
        );

    \I__6298\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27946\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__27953\,
            I => \N__27943\
        );

    \I__6296\ : Span4Mux_h
    port map (
            O => \N__27950\,
            I => \N__27940\
        );

    \I__6295\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27937\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__27946\,
            I => data_in_3_5
        );

    \I__6293\ : Odrv4
    port map (
            O => \N__27943\,
            I => data_in_3_5
        );

    \I__6292\ : Odrv4
    port map (
            O => \N__27940\,
            I => data_in_3_5
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__27937\,
            I => data_in_3_5
        );

    \I__6290\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27923\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__27927\,
            I => \N__27920\
        );

    \I__6288\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27916\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27913\
        );

    \I__6286\ : InMux
    port map (
            O => \N__27920\,
            I => \N__27910\
        );

    \I__6285\ : InMux
    port map (
            O => \N__27919\,
            I => \N__27907\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27904\
        );

    \I__6283\ : Span4Mux_v
    port map (
            O => \N__27913\,
            I => \N__27899\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__27910\,
            I => \N__27899\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__27907\,
            I => data_in_3_4
        );

    \I__6280\ : Odrv12
    port map (
            O => \N__27904\,
            I => data_in_3_4
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__27899\,
            I => data_in_3_4
        );

    \I__6278\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27888\
        );

    \I__6277\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27885\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__27888\,
            I => \N__27882\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__27885\,
            I => \N__27879\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__27882\,
            I => \N__27876\
        );

    \I__6273\ : Span4Mux_h
    port map (
            O => \N__27879\,
            I => \N__27873\
        );

    \I__6272\ : Span4Mux_h
    port map (
            O => \N__27876\,
            I => \N__27870\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__27873\,
            I => \N__27865\
        );

    \I__6270\ : Sp12to4
    port map (
            O => \N__27870\,
            I => \N__27862\
        );

    \I__6269\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27857\
        );

    \I__6268\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27857\
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__27865\,
            I => data_in_2_6
        );

    \I__6266\ : Odrv12
    port map (
            O => \N__27862\,
            I => data_in_2_6
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__27857\,
            I => data_in_2_6
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__27850\,
            I => \N__27847\
        );

    \I__6263\ : InMux
    port map (
            O => \N__27847\,
            I => \N__27844\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__27844\,
            I => \N__27841\
        );

    \I__6261\ : Span4Mux_h
    port map (
            O => \N__27841\,
            I => \N__27838\
        );

    \I__6260\ : Span4Mux_h
    port map (
            O => \N__27838\,
            I => \N__27832\
        );

    \I__6259\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27825\
        );

    \I__6258\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27825\
        );

    \I__6257\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27825\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__27832\,
            I => data_in_3_6
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__27825\,
            I => data_in_3_6
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__27820\,
            I => \c0.n28_adj_1953_cascade_\
        );

    \I__6253\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27814\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__27814\,
            I => \c0.n22_adj_1952\
        );

    \I__6251\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__6249\ : Odrv12
    port map (
            O => \N__27805\,
            I => \c0.n30_adj_1959\
        );

    \I__6248\ : CascadeMux
    port map (
            O => \N__27802\,
            I => \N__27799\
        );

    \I__6247\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27792\
        );

    \I__6245\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27789\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__27792\,
            I => \N__27785\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27782\
        );

    \I__6242\ : InMux
    port map (
            O => \N__27788\,
            I => \N__27779\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__27785\,
            I => data_in_4_5
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__27782\,
            I => data_in_4_5
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__27779\,
            I => data_in_4_5
        );

    \I__6238\ : CascadeMux
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__6237\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27763\
        );

    \I__6236\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27763\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27760\
        );

    \I__6234\ : Span4Mux_h
    port map (
            O => \N__27760\,
            I => \N__27756\
        );

    \I__6233\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27753\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__27756\,
            I => data_in_8_0
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__27753\,
            I => data_in_8_0
        );

    \I__6230\ : CascadeMux
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__6229\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27741\
        );

    \I__6228\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27738\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27734\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__27738\,
            I => \N__27731\
        );

    \I__6225\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27728\
        );

    \I__6224\ : Odrv12
    port map (
            O => \N__27734\,
            I => data_in_5_7
        );

    \I__6223\ : Odrv4
    port map (
            O => \N__27731\,
            I => data_in_5_7
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__27728\,
            I => data_in_5_7
        );

    \I__6221\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27717\
        );

    \I__6220\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27714\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__27717\,
            I => \N__27710\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__27714\,
            I => \N__27707\
        );

    \I__6217\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27703\
        );

    \I__6216\ : Span4Mux_h
    port map (
            O => \N__27710\,
            I => \N__27698\
        );

    \I__6215\ : Span4Mux_v
    port map (
            O => \N__27707\,
            I => \N__27698\
        );

    \I__6214\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27695\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__27703\,
            I => \c0.data_in_field_47\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__27698\,
            I => \c0.data_in_field_47\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__27695\,
            I => \c0.data_in_field_47\
        );

    \I__6210\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27684\
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__27687\,
            I => \N__27681\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27678\
        );

    \I__6207\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27674\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__27678\,
            I => \N__27671\
        );

    \I__6205\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27668\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__27674\,
            I => data_in_15_7
        );

    \I__6203\ : Odrv4
    port map (
            O => \N__27671\,
            I => data_in_15_7
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__27668\,
            I => data_in_15_7
        );

    \I__6201\ : InMux
    port map (
            O => \N__27661\,
            I => \N__27658\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__27658\,
            I => \N__27654\
        );

    \I__6199\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27651\
        );

    \I__6198\ : Span4Mux_h
    port map (
            O => \N__27654\,
            I => \N__27645\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27645\
        );

    \I__6196\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27642\
        );

    \I__6195\ : Span4Mux_v
    port map (
            O => \N__27645\,
            I => \N__27637\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27634\
        );

    \I__6193\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27631\
        );

    \I__6192\ : InMux
    port map (
            O => \N__27640\,
            I => \N__27628\
        );

    \I__6191\ : Span4Mux_h
    port map (
            O => \N__27637\,
            I => \N__27625\
        );

    \I__6190\ : Span4Mux_h
    port map (
            O => \N__27634\,
            I => \N__27622\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__27631\,
            I => \c0.data_in_field_127\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__27628\,
            I => \c0.data_in_field_127\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__27625\,
            I => \c0.data_in_field_127\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__27622\,
            I => \c0.data_in_field_127\
        );

    \I__6185\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27609\
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__27612\,
            I => \N__27605\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__27609\,
            I => \N__27602\
        );

    \I__6182\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27599\
        );

    \I__6181\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27596\
        );

    \I__6180\ : Span4Mux_h
    port map (
            O => \N__27602\,
            I => \N__27593\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__27599\,
            I => data_in_16_0
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__27596\,
            I => data_in_16_0
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__27593\,
            I => data_in_16_0
        );

    \I__6176\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27582\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__27585\,
            I => \N__27579\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__27582\,
            I => \N__27574\
        );

    \I__6173\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27571\
        );

    \I__6172\ : InMux
    port map (
            O => \N__27578\,
            I => \N__27568\
        );

    \I__6171\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27565\
        );

    \I__6170\ : Span12Mux_h
    port map (
            O => \N__27574\,
            I => \N__27562\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__27571\,
            I => \N__27559\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__27568\,
            I => data_in_1_7
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__27565\,
            I => data_in_1_7
        );

    \I__6166\ : Odrv12
    port map (
            O => \N__27562\,
            I => data_in_1_7
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__27559\,
            I => data_in_1_7
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__27550\,
            I => \N__27547\
        );

    \I__6163\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27543\
        );

    \I__6162\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27540\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__27543\,
            I => \N__27537\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27534\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__27537\,
            I => \N__27529\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__27534\,
            I => \N__27529\
        );

    \I__6157\ : Sp12to4
    port map (
            O => \N__27529\,
            I => \N__27525\
        );

    \I__6156\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27522\
        );

    \I__6155\ : Odrv12
    port map (
            O => \N__27525\,
            I => data_in_10_5
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__27522\,
            I => data_in_10_5
        );

    \I__6153\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27514\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27510\
        );

    \I__6151\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27506\
        );

    \I__6150\ : Span4Mux_h
    port map (
            O => \N__27510\,
            I => \N__27503\
        );

    \I__6149\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27500\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__27506\,
            I => data_in_9_5
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__27503\,
            I => data_in_9_5
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__27500\,
            I => data_in_9_5
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__27493\,
            I => \N__27490\
        );

    \I__6144\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27485\
        );

    \I__6143\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27482\
        );

    \I__6142\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27479\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__27485\,
            I => \N__27476\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__27482\,
            I => \N__27473\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__27479\,
            I => data_in_0_5
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__27476\,
            I => data_in_0_5
        );

    \I__6137\ : Odrv12
    port map (
            O => \N__27473\,
            I => data_in_0_5
        );

    \I__6136\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27463\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__27463\,
            I => \N__27460\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__27460\,
            I => \N__27457\
        );

    \I__6133\ : Span4Mux_h
    port map (
            O => \N__27457\,
            I => \N__27451\
        );

    \I__6132\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27446\
        );

    \I__6131\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27446\
        );

    \I__6130\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27443\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__27451\,
            I => data_in_1_2
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__27446\,
            I => data_in_1_2
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__27443\,
            I => data_in_1_2
        );

    \I__6126\ : CascadeMux
    port map (
            O => \N__27436\,
            I => \c0.n6_adj_1876_cascade_\
        );

    \I__6125\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27430\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27427\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__27427\,
            I => \N__27421\
        );

    \I__6122\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27418\
        );

    \I__6121\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27415\
        );

    \I__6120\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27411\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__27421\,
            I => \N__27406\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27406\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__27415\,
            I => \N__27403\
        );

    \I__6116\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27400\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__27411\,
            I => \c0.data_in_field_132\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__27406\,
            I => \c0.data_in_field_132\
        );

    \I__6113\ : Odrv12
    port map (
            O => \N__27403\,
            I => \c0.data_in_field_132\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__27400\,
            I => \c0.data_in_field_132\
        );

    \I__6111\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__27388\,
            I => \N__27385\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__27385\,
            I => \N__27382\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__27382\,
            I => \N__27378\
        );

    \I__6107\ : InMux
    port map (
            O => \N__27381\,
            I => \N__27375\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__27378\,
            I => \c0.n5129\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__27375\,
            I => \c0.n5129\
        );

    \I__6104\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__27367\,
            I => \N__27364\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__27364\,
            I => \c0.n6_adj_1874\
        );

    \I__6101\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27358\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__27358\,
            I => \N__27355\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__27355\,
            I => \N__27350\
        );

    \I__6098\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27345\
        );

    \I__6097\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27345\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__27350\,
            I => data_in_0_0
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__27345\,
            I => data_in_0_0
        );

    \I__6094\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27337\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27331\
        );

    \I__6092\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27324\
        );

    \I__6091\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27324\
        );

    \I__6090\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27324\
        );

    \I__6089\ : Odrv4
    port map (
            O => \N__27331\,
            I => \c0.data_in_field_0\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__27324\,
            I => \c0.data_in_field_0\
        );

    \I__6087\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27315\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__27318\,
            I => \N__27312\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__27315\,
            I => \N__27307\
        );

    \I__6084\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27304\
        );

    \I__6083\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27301\
        );

    \I__6082\ : CascadeMux
    port map (
            O => \N__27310\,
            I => \N__27298\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__27307\,
            I => \N__27291\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27291\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__27301\,
            I => \N__27288\
        );

    \I__6078\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27285\
        );

    \I__6077\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27282\
        );

    \I__6076\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27279\
        );

    \I__6075\ : Span4Mux_h
    port map (
            O => \N__27291\,
            I => \N__27276\
        );

    \I__6074\ : Span4Mux_h
    port map (
            O => \N__27288\,
            I => \N__27273\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__27285\,
            I => \c0.data_in_field_90\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__27282\,
            I => \c0.data_in_field_90\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__27279\,
            I => \c0.data_in_field_90\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__27276\,
            I => \c0.data_in_field_90\
        );

    \I__6069\ : Odrv4
    port map (
            O => \N__27273\,
            I => \c0.data_in_field_90\
        );

    \I__6068\ : InMux
    port map (
            O => \N__27262\,
            I => \N__27259\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__27259\,
            I => \N__27256\
        );

    \I__6066\ : Span4Mux_h
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__27253\,
            I => \c0.n22_adj_1935\
        );

    \I__6064\ : CascadeMux
    port map (
            O => \N__27250\,
            I => \N__27247\
        );

    \I__6063\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27244\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__27244\,
            I => \N__27241\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__27241\,
            I => \N__27236\
        );

    \I__6060\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27231\
        );

    \I__6059\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27231\
        );

    \I__6058\ : Odrv4
    port map (
            O => \N__27236\,
            I => data_in_5_6
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__27231\,
            I => data_in_5_6
        );

    \I__6056\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27222\
        );

    \I__6055\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27219\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__27222\,
            I => \N__27214\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__27219\,
            I => \N__27211\
        );

    \I__6052\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27208\
        );

    \I__6051\ : InMux
    port map (
            O => \N__27217\,
            I => \N__27205\
        );

    \I__6050\ : Span4Mux_v
    port map (
            O => \N__27214\,
            I => \N__27202\
        );

    \I__6049\ : Span12Mux_s9_h
    port map (
            O => \N__27211\,
            I => \N__27199\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__27208\,
            I => \N__27196\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__27205\,
            I => \c0.data_in_field_2\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__27202\,
            I => \c0.data_in_field_2\
        );

    \I__6045\ : Odrv12
    port map (
            O => \N__27199\,
            I => \c0.data_in_field_2\
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__27196\,
            I => \c0.data_in_field_2\
        );

    \I__6043\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__27184\,
            I => \N__27181\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__27181\,
            I => \N__27175\
        );

    \I__6040\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27172\
        );

    \I__6039\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27169\
        );

    \I__6038\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27166\
        );

    \I__6037\ : Span4Mux_h
    port map (
            O => \N__27175\,
            I => \N__27161\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__27172\,
            I => \N__27161\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__27169\,
            I => \c0.data_in_field_108\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__27166\,
            I => \c0.data_in_field_108\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__27161\,
            I => \c0.data_in_field_108\
        );

    \I__6032\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27151\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__27151\,
            I => \N__27147\
        );

    \I__6030\ : InMux
    port map (
            O => \N__27150\,
            I => \N__27144\
        );

    \I__6029\ : Odrv12
    port map (
            O => \N__27147\,
            I => \c0.n5102\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__27144\,
            I => \c0.n5102\
        );

    \I__6027\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27134\
        );

    \I__6026\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27131\
        );

    \I__6025\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27127\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27123\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__27131\,
            I => \N__27120\
        );

    \I__6022\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27117\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__27127\,
            I => \N__27114\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__27126\,
            I => \N__27110\
        );

    \I__6019\ : Span12Mux_v
    port map (
            O => \N__27123\,
            I => \N__27107\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__27120\,
            I => \N__27104\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27099\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__27114\,
            I => \N__27099\
        );

    \I__6015\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27094\
        );

    \I__6014\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27094\
        );

    \I__6013\ : Odrv12
    port map (
            O => \N__27107\,
            I => \c0.data_in_field_142\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__27104\,
            I => \c0.data_in_field_142\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__27099\,
            I => \c0.data_in_field_142\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__27094\,
            I => \c0.data_in_field_142\
        );

    \I__6009\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27082\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27078\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__27081\,
            I => \N__27075\
        );

    \I__6006\ : Span12Mux_v
    port map (
            O => \N__27078\,
            I => \N__27072\
        );

    \I__6005\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27069\
        );

    \I__6004\ : Odrv12
    port map (
            O => \N__27072\,
            I => \c0.n1795\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__27069\,
            I => \c0.n1795\
        );

    \I__6002\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__27061\,
            I => \N__27058\
        );

    \I__6000\ : Odrv12
    port map (
            O => \N__27058\,
            I => \c0.n11_adj_1913\
        );

    \I__5999\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27051\
        );

    \I__5998\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27048\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27051\,
            I => \N__27045\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__27048\,
            I => \N__27042\
        );

    \I__5995\ : Span4Mux_v
    port map (
            O => \N__27045\,
            I => \N__27039\
        );

    \I__5994\ : Span4Mux_h
    port map (
            O => \N__27042\,
            I => \N__27035\
        );

    \I__5993\ : Span4Mux_h
    port map (
            O => \N__27039\,
            I => \N__27032\
        );

    \I__5992\ : InMux
    port map (
            O => \N__27038\,
            I => \N__27029\
        );

    \I__5991\ : Span4Mux_h
    port map (
            O => \N__27035\,
            I => \N__27026\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__27032\,
            I => \N__27023\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__27029\,
            I => data_in_11_4
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__27026\,
            I => data_in_11_4
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__27023\,
            I => data_in_11_4
        );

    \I__5986\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__27009\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27012\,
            I => \N__27006\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__27009\,
            I => \N__27003\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__27006\,
            I => \N__27000\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__27003\,
            I => \N__26993\
        );

    \I__5980\ : Span4Mux_v
    port map (
            O => \N__27000\,
            I => \N__26993\
        );

    \I__5979\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26988\
        );

    \I__5978\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26988\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__26993\,
            I => \c0.data_in_field_92\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__26988\,
            I => \c0.data_in_field_92\
        );

    \I__5975\ : CascadeMux
    port map (
            O => \N__26983\,
            I => \N__26979\
        );

    \I__5974\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26975\
        );

    \I__5973\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26970\
        );

    \I__5972\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26970\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__26975\,
            I => \N__26967\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__26970\,
            I => \N__26964\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__26967\,
            I => \N__26961\
        );

    \I__5968\ : Span4Mux_v
    port map (
            O => \N__26964\,
            I => \N__26956\
        );

    \I__5967\ : Span4Mux_h
    port map (
            O => \N__26961\,
            I => \N__26956\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__26956\,
            I => data_in_11_5
        );

    \I__5965\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__26950\,
            I => \N__26947\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__26947\,
            I => \N__26942\
        );

    \I__5962\ : InMux
    port map (
            O => \N__26946\,
            I => \N__26937\
        );

    \I__5961\ : InMux
    port map (
            O => \N__26945\,
            I => \N__26937\
        );

    \I__5960\ : Span4Mux_h
    port map (
            O => \N__26942\,
            I => \N__26931\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26931\
        );

    \I__5958\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26927\
        );

    \I__5957\ : Span4Mux_h
    port map (
            O => \N__26931\,
            I => \N__26924\
        );

    \I__5956\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26921\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__26927\,
            I => \c0.data_in_field_93\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__26924\,
            I => \c0.data_in_field_93\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__26921\,
            I => \c0.data_in_field_93\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__5951\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__26908\,
            I => \c0.n5707\
        );

    \I__5949\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26902\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__26902\,
            I => \N__26898\
        );

    \I__5947\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26895\
        );

    \I__5946\ : Span4Mux_v
    port map (
            O => \N__26898\,
            I => \N__26891\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26888\
        );

    \I__5944\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26885\
        );

    \I__5943\ : Odrv4
    port map (
            O => \N__26891\,
            I => \c0.n1838\
        );

    \I__5942\ : Odrv12
    port map (
            O => \N__26888\,
            I => \c0.n1838\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__26885\,
            I => \c0.n1838\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__26878\,
            I => \N__26875\
        );

    \I__5939\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26871\
        );

    \I__5938\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26868\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__26871\,
            I => \N__26865\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26862\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__26865\,
            I => \N__26858\
        );

    \I__5934\ : Span4Mux_s3_v
    port map (
            O => \N__26862\,
            I => \N__26855\
        );

    \I__5933\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26852\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__26858\,
            I => data_in_5_0
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__26855\,
            I => data_in_5_0
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__26852\,
            I => data_in_5_0
        );

    \I__5929\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26842\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__26842\,
            I => \N__26839\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__26839\,
            I => \N__26836\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__26836\,
            I => \N__26832\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__26835\,
            I => \N__26828\
        );

    \I__5924\ : Span4Mux_h
    port map (
            O => \N__26832\,
            I => \N__26825\
        );

    \I__5923\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26822\
        );

    \I__5922\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26819\
        );

    \I__5921\ : Span4Mux_h
    port map (
            O => \N__26825\,
            I => \N__26816\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__26822\,
            I => data_in_16_3
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__26819\,
            I => data_in_16_3
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__26816\,
            I => data_in_16_3
        );

    \I__5917\ : CascadeMux
    port map (
            O => \N__26809\,
            I => \N__26804\
        );

    \I__5916\ : CascadeMux
    port map (
            O => \N__26808\,
            I => \N__26801\
        );

    \I__5915\ : InMux
    port map (
            O => \N__26807\,
            I => \N__26796\
        );

    \I__5914\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26796\
        );

    \I__5913\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26792\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__26796\,
            I => \N__26789\
        );

    \I__5911\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26786\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__26792\,
            I => \N__26783\
        );

    \I__5909\ : Sp12to4
    port map (
            O => \N__26789\,
            I => \N__26780\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__26786\,
            I => \N__26777\
        );

    \I__5907\ : Span4Mux_h
    port map (
            O => \N__26783\,
            I => \N__26774\
        );

    \I__5906\ : Span12Mux_v
    port map (
            O => \N__26780\,
            I => \N__26771\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__26777\,
            I => data_in_18_4
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__26774\,
            I => data_in_18_4
        );

    \I__5903\ : Odrv12
    port map (
            O => \N__26771\,
            I => data_in_18_4
        );

    \I__5902\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26760\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__26763\,
            I => \N__26756\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26753\
        );

    \I__5899\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26748\
        );

    \I__5898\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26748\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__26753\,
            I => \N__26745\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__26748\,
            I => data_in_17_4
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__26745\,
            I => data_in_17_4
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__26740\,
            I => \N__26737\
        );

    \I__5893\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26734\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__26734\,
            I => \N__26731\
        );

    \I__5891\ : Span4Mux_h
    port map (
            O => \N__26731\,
            I => \N__26725\
        );

    \I__5890\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26722\
        );

    \I__5889\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26719\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26716\
        );

    \I__5887\ : Span4Mux_v
    port map (
            O => \N__26725\,
            I => \N__26712\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__26722\,
            I => \N__26709\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26706\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__26716\,
            I => \N__26703\
        );

    \I__5883\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26699\
        );

    \I__5882\ : IoSpan4Mux
    port map (
            O => \N__26712\,
            I => \N__26696\
        );

    \I__5881\ : Span4Mux_h
    port map (
            O => \N__26709\,
            I => \N__26693\
        );

    \I__5880\ : Span4Mux_v
    port map (
            O => \N__26706\,
            I => \N__26690\
        );

    \I__5879\ : Span4Mux_h
    port map (
            O => \N__26703\,
            I => \N__26687\
        );

    \I__5878\ : InMux
    port map (
            O => \N__26702\,
            I => \N__26684\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__26699\,
            I => \c0.data_in_field_63\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__26696\,
            I => \c0.data_in_field_63\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__26693\,
            I => \c0.data_in_field_63\
        );

    \I__5874\ : Odrv4
    port map (
            O => \N__26690\,
            I => \c0.data_in_field_63\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__26687\,
            I => \c0.data_in_field_63\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__26684\,
            I => \c0.data_in_field_63\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__26671\,
            I => \N__26668\
        );

    \I__5870\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__26665\,
            I => \N__26660\
        );

    \I__5868\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26657\
        );

    \I__5867\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26652\
        );

    \I__5866\ : Span4Mux_h
    port map (
            O => \N__26660\,
            I => \N__26647\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__26657\,
            I => \N__26647\
        );

    \I__5864\ : InMux
    port map (
            O => \N__26656\,
            I => \N__26644\
        );

    \I__5863\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26641\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__26652\,
            I => \c0.data_in_field_62\
        );

    \I__5861\ : Odrv4
    port map (
            O => \N__26647\,
            I => \c0.data_in_field_62\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__26644\,
            I => \c0.data_in_field_62\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__26641\,
            I => \c0.data_in_field_62\
        );

    \I__5858\ : CascadeMux
    port map (
            O => \N__26632\,
            I => \c0.n1795_cascade_\
        );

    \I__5857\ : InMux
    port map (
            O => \N__26629\,
            I => \N__26626\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__5855\ : Odrv12
    port map (
            O => \N__26623\,
            I => \c0.n6097\
        );

    \I__5854\ : CascadeMux
    port map (
            O => \N__26620\,
            I => \N__26616\
        );

    \I__5853\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26613\
        );

    \I__5852\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26610\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__26613\,
            I => \N__26607\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__26610\,
            I => \N__26604\
        );

    \I__5849\ : Span4Mux_h
    port map (
            O => \N__26607\,
            I => \N__26601\
        );

    \I__5848\ : Span12Mux_h
    port map (
            O => \N__26604\,
            I => \N__26597\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__26601\,
            I => \N__26594\
        );

    \I__5846\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26591\
        );

    \I__5845\ : Odrv12
    port map (
            O => \N__26597\,
            I => data_in_6_3
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__26594\,
            I => data_in_6_3
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__26591\,
            I => data_in_6_3
        );

    \I__5842\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26581\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__5840\ : Span4Mux_s1_v
    port map (
            O => \N__26578\,
            I => \N__26575\
        );

    \I__5839\ : Sp12to4
    port map (
            O => \N__26575\,
            I => \N__26571\
        );

    \I__5838\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26567\
        );

    \I__5837\ : Span12Mux_s10_h
    port map (
            O => \N__26571\,
            I => \N__26564\
        );

    \I__5836\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26561\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__26567\,
            I => data_in_5_3
        );

    \I__5834\ : Odrv12
    port map (
            O => \N__26564\,
            I => data_in_5_3
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__26561\,
            I => data_in_5_3
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__26554\,
            I => \N__26551\
        );

    \I__5831\ : InMux
    port map (
            O => \N__26551\,
            I => \N__26548\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__26548\,
            I => \N__26545\
        );

    \I__5829\ : Span4Mux_h
    port map (
            O => \N__26545\,
            I => \N__26542\
        );

    \I__5828\ : Span4Mux_h
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__26539\,
            I => \N__26534\
        );

    \I__5826\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26529\
        );

    \I__5825\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26529\
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__26534\,
            I => data_in_9_1
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__26529\,
            I => data_in_9_1
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__26524\,
            I => \N__26520\
        );

    \I__5821\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26517\
        );

    \I__5820\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26514\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__26517\,
            I => \N__26511\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__26514\,
            I => \N__26505\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__26511\,
            I => \N__26505\
        );

    \I__5816\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26502\
        );

    \I__5815\ : Odrv4
    port map (
            O => \N__26505\,
            I => data_in_7_6
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__26502\,
            I => data_in_7_6
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__26497\,
            I => \N__26493\
        );

    \I__5812\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26490\
        );

    \I__5811\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26486\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__26490\,
            I => \N__26483\
        );

    \I__5809\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26480\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__26486\,
            I => data_in_10_4
        );

    \I__5807\ : Odrv12
    port map (
            O => \N__26483\,
            I => data_in_10_4
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__26480\,
            I => data_in_10_4
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__26473\,
            I => \N__26470\
        );

    \I__5804\ : InMux
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__26467\,
            I => \N__26464\
        );

    \I__5802\ : Span4Mux_h
    port map (
            O => \N__26464\,
            I => \N__26461\
        );

    \I__5801\ : Span4Mux_h
    port map (
            O => \N__26461\,
            I => \N__26458\
        );

    \I__5800\ : Span4Mux_v
    port map (
            O => \N__26458\,
            I => \N__26453\
        );

    \I__5799\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26448\
        );

    \I__5798\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26448\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__26453\,
            I => data_in_10_3
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__26448\,
            I => data_in_10_3
        );

    \I__5795\ : InMux
    port map (
            O => \N__26443\,
            I => \N__26439\
        );

    \I__5794\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26436\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__26439\,
            I => \N__26433\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__26436\,
            I => \N__26429\
        );

    \I__5791\ : Sp12to4
    port map (
            O => \N__26433\,
            I => \N__26426\
        );

    \I__5790\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26423\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__26429\,
            I => data_in_9_3
        );

    \I__5788\ : Odrv12
    port map (
            O => \N__26426\,
            I => data_in_9_3
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__26423\,
            I => data_in_9_3
        );

    \I__5786\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26413\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26410\
        );

    \I__5784\ : Span4Mux_h
    port map (
            O => \N__26410\,
            I => \N__26407\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__26407\,
            I => \c0.n26_adj_1878\
        );

    \I__5782\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26401\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__26401\,
            I => \N__26398\
        );

    \I__5780\ : Span4Mux_h
    port map (
            O => \N__26398\,
            I => \N__26395\
        );

    \I__5779\ : Span4Mux_v
    port map (
            O => \N__26395\,
            I => \N__26390\
        );

    \I__5778\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26385\
        );

    \I__5777\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26385\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__26390\,
            I => data_in_0_4
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__26385\,
            I => data_in_0_4
        );

    \I__5774\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26376\
        );

    \I__5773\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26372\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__26376\,
            I => \N__26369\
        );

    \I__5771\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26366\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26361\
        );

    \I__5769\ : Span4Mux_h
    port map (
            O => \N__26369\,
            I => \N__26356\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__26366\,
            I => \N__26356\
        );

    \I__5767\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26352\
        );

    \I__5766\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26349\
        );

    \I__5765\ : Span4Mux_v
    port map (
            O => \N__26361\,
            I => \N__26344\
        );

    \I__5764\ : Span4Mux_v
    port map (
            O => \N__26356\,
            I => \N__26344\
        );

    \I__5763\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26341\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__26352\,
            I => \N__26338\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__26349\,
            I => \c0.data_in_field_68\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__26344\,
            I => \c0.data_in_field_68\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__26341\,
            I => \c0.data_in_field_68\
        );

    \I__5758\ : Odrv12
    port map (
            O => \N__26338\,
            I => \c0.data_in_field_68\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__5756\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26322\
        );

    \I__5755\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26319\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N__26316\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__26319\,
            I => \N__26313\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__26316\,
            I => \N__26310\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__26313\,
            I => \N__26307\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__26310\,
            I => \c0.n5105\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__26307\,
            I => \c0.n5105\
        );

    \I__5748\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26299\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__26299\,
            I => \N__26296\
        );

    \I__5746\ : Span4Mux_v
    port map (
            O => \N__26296\,
            I => \N__26292\
        );

    \I__5745\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26289\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__26292\,
            I => \c0.n5111\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__26289\,
            I => \c0.n5111\
        );

    \I__5742\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26281\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__26281\,
            I => \N__26278\
        );

    \I__5740\ : Span12Mux_s10_h
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__5739\ : Odrv12
    port map (
            O => \N__26275\,
            I => \c0.n35\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__26272\,
            I => \N__26268\
        );

    \I__5737\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26265\
        );

    \I__5736\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26261\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__26265\,
            I => \N__26257\
        );

    \I__5734\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26254\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26251\
        );

    \I__5732\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26248\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__26257\,
            I => \N__26242\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26242\
        );

    \I__5729\ : Span4Mux_h
    port map (
            O => \N__26251\,
            I => \N__26237\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__26248\,
            I => \N__26237\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__26247\,
            I => \N__26234\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__26242\,
            I => \N__26229\
        );

    \I__5725\ : Span4Mux_v
    port map (
            O => \N__26237\,
            I => \N__26229\
        );

    \I__5724\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26226\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__26229\,
            I => \N__26223\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__26226\,
            I => \c0.data_in_field_59\
        );

    \I__5721\ : Odrv4
    port map (
            O => \N__26223\,
            I => \c0.data_in_field_59\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__26218\,
            I => \N__26215\
        );

    \I__5719\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26211\
        );

    \I__5718\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26208\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__26211\,
            I => \N__26205\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26202\
        );

    \I__5715\ : Span4Mux_v
    port map (
            O => \N__26205\,
            I => \N__26199\
        );

    \I__5714\ : Span4Mux_s1_v
    port map (
            O => \N__26202\,
            I => \N__26196\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__26199\,
            I => \N__26190\
        );

    \I__5712\ : Span4Mux_v
    port map (
            O => \N__26196\,
            I => \N__26190\
        );

    \I__5711\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26187\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__26190\,
            I => data_in_6_6
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__26187\,
            I => data_in_6_6
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__26182\,
            I => \N__26179\
        );

    \I__5707\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26175\
        );

    \I__5706\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26172\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__26175\,
            I => \N__26167\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26167\
        );

    \I__5703\ : Span12Mux_s10_v
    port map (
            O => \N__26167\,
            I => \N__26163\
        );

    \I__5702\ : InMux
    port map (
            O => \N__26166\,
            I => \N__26160\
        );

    \I__5701\ : Odrv12
    port map (
            O => \N__26163\,
            I => data_in_13_4
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__26160\,
            I => data_in_13_4
        );

    \I__5699\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26151\
        );

    \I__5698\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26147\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__26151\,
            I => \N__26144\
        );

    \I__5696\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26140\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__26147\,
            I => \N__26137\
        );

    \I__5694\ : Span4Mux_v
    port map (
            O => \N__26144\,
            I => \N__26134\
        );

    \I__5693\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26131\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__26140\,
            I => \N__26128\
        );

    \I__5691\ : Span12Mux_s8_v
    port map (
            O => \N__26137\,
            I => \N__26125\
        );

    \I__5690\ : Span4Mux_h
    port map (
            O => \N__26134\,
            I => \N__26118\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26118\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__26128\,
            I => \N__26118\
        );

    \I__5687\ : Odrv12
    port map (
            O => \N__26125\,
            I => data_in_2_4
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__26118\,
            I => data_in_2_4
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__26113\,
            I => \N__26108\
        );

    \I__5684\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26105\
        );

    \I__5683\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26102\
        );

    \I__5682\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26098\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__26105\,
            I => \N__26095\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26092\
        );

    \I__5679\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26088\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__26098\,
            I => \N__26085\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__26095\,
            I => \N__26082\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__26092\,
            I => \N__26079\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__26091\,
            I => \N__26076\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26071\
        );

    \I__5673\ : Span4Mux_v
    port map (
            O => \N__26085\,
            I => \N__26071\
        );

    \I__5672\ : Span4Mux_h
    port map (
            O => \N__26082\,
            I => \N__26066\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__26079\,
            I => \N__26066\
        );

    \I__5670\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26063\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__26071\,
            I => \N__26060\
        );

    \I__5668\ : Span4Mux_v
    port map (
            O => \N__26066\,
            I => \N__26057\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__26063\,
            I => \c0.data_in_field_115\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__26060\,
            I => \c0.data_in_field_115\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__26057\,
            I => \c0.data_in_field_115\
        );

    \I__5664\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26047\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__5662\ : Span4Mux_s2_v
    port map (
            O => \N__26044\,
            I => \N__26040\
        );

    \I__5661\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26035\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__26040\,
            I => \N__26032\
        );

    \I__5659\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26027\
        );

    \I__5658\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26027\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__26035\,
            I => data_in_18_7
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__26032\,
            I => data_in_18_7
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__26027\,
            I => data_in_18_7
        );

    \I__5654\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26013\
        );

    \I__5653\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26013\
        );

    \I__5652\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26010\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__26013\,
            I => data_in_17_7
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__26010\,
            I => data_in_17_7
        );

    \I__5649\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25999\
        );

    \I__5648\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25999\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__25999\,
            I => \N__25994\
        );

    \I__5646\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25991\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__25997\,
            I => \N__25988\
        );

    \I__5644\ : Span4Mux_v
    port map (
            O => \N__25994\,
            I => \N__25985\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25982\
        );

    \I__5642\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25978\
        );

    \I__5641\ : Span4Mux_s2_v
    port map (
            O => \N__25985\,
            I => \N__25975\
        );

    \I__5640\ : Span12Mux_v
    port map (
            O => \N__25982\,
            I => \N__25972\
        );

    \I__5639\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25969\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__25978\,
            I => \c0.data_in_field_49\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__25975\,
            I => \c0.data_in_field_49\
        );

    \I__5636\ : Odrv12
    port map (
            O => \N__25972\,
            I => \c0.data_in_field_49\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__25969\,
            I => \c0.data_in_field_49\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__25960\,
            I => \c0.n2092_cascade_\
        );

    \I__5633\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25953\
        );

    \I__5632\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25950\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__25953\,
            I => \N__25947\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25944\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__25947\,
            I => \c0.n2043\
        );

    \I__5628\ : Odrv12
    port map (
            O => \N__25944\,
            I => \c0.n2043\
        );

    \I__5627\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25935\
        );

    \I__5626\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25932\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25929\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__25932\,
            I => \N__25926\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__25929\,
            I => \N__25923\
        );

    \I__5622\ : Span4Mux_v
    port map (
            O => \N__25926\,
            I => \N__25920\
        );

    \I__5621\ : Span4Mux_h
    port map (
            O => \N__25923\,
            I => \N__25917\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__25920\,
            I => \c0.n5246\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__25917\,
            I => \c0.n5246\
        );

    \I__5618\ : CascadeMux
    port map (
            O => \N__25912\,
            I => \N__25908\
        );

    \I__5617\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25904\
        );

    \I__5616\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25901\
        );

    \I__5615\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25898\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__25904\,
            I => \N__25895\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__25901\,
            I => \N__25892\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__25898\,
            I => data_in_0_2
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__25895\,
            I => data_in_0_2
        );

    \I__5610\ : Odrv12
    port map (
            O => \N__25892\,
            I => data_in_0_2
        );

    \I__5609\ : InMux
    port map (
            O => \N__25885\,
            I => \N__25882\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__25882\,
            I => \N__25878\
        );

    \I__5607\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25875\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__25878\,
            I => \N__25872\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__25875\,
            I => \N__25867\
        );

    \I__5604\ : Span4Mux_h
    port map (
            O => \N__25872\,
            I => \N__25864\
        );

    \I__5603\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25859\
        );

    \I__5602\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25859\
        );

    \I__5601\ : Odrv4
    port map (
            O => \N__25867\,
            I => \c0.data_in_field_9\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__25864\,
            I => \c0.data_in_field_9\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25859\,
            I => \c0.data_in_field_9\
        );

    \I__5598\ : CascadeMux
    port map (
            O => \N__25852\,
            I => \N__25849\
        );

    \I__5597\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25846\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__25846\,
            I => \N__25843\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__25843\,
            I => \N__25840\
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__25840\,
            I => \c0.n5749\
        );

    \I__5593\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25832\
        );

    \I__5592\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25827\
        );

    \I__5591\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25827\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__25832\,
            I => \c0.data_in_field_1\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__25827\,
            I => \c0.data_in_field_1\
        );

    \I__5588\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25819\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__5586\ : Span12Mux_v
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__5585\ : Odrv12
    port map (
            O => \N__25813\,
            I => \c0.n5453\
        );

    \I__5584\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25806\
        );

    \I__5583\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25803\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__25806\,
            I => \N__25800\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__25803\,
            I => \N__25797\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__25800\,
            I => \N__25792\
        );

    \I__5579\ : Span4Mux_v
    port map (
            O => \N__25797\,
            I => \N__25792\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__25792\,
            I => \N__25788\
        );

    \I__5577\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25785\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__25788\,
            I => \c0.n1830\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__25785\,
            I => \c0.n1830\
        );

    \I__5574\ : InMux
    port map (
            O => \N__25780\,
            I => \N__25777\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__25777\,
            I => \c0.n5141\
        );

    \I__5572\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25771\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__25771\,
            I => \N__25767\
        );

    \I__5570\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25764\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__25767\,
            I => \N__25760\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__25764\,
            I => \N__25756\
        );

    \I__5567\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25753\
        );

    \I__5566\ : Span4Mux_v
    port map (
            O => \N__25760\,
            I => \N__25750\
        );

    \I__5565\ : InMux
    port map (
            O => \N__25759\,
            I => \N__25746\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__25756\,
            I => \N__25741\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25741\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__25750\,
            I => \N__25738\
        );

    \I__5561\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25735\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__25746\,
            I => \c0.data_in_field_106\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__25741\,
            I => \c0.data_in_field_106\
        );

    \I__5558\ : Odrv4
    port map (
            O => \N__25738\,
            I => \c0.data_in_field_106\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__25735\,
            I => \c0.data_in_field_106\
        );

    \I__5556\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25722\
        );

    \I__5555\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25719\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__25722\,
            I => \N__25715\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__25719\,
            I => \N__25712\
        );

    \I__5552\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25709\
        );

    \I__5551\ : Odrv12
    port map (
            O => \N__25715\,
            I => data_in_13_7
        );

    \I__5550\ : Odrv4
    port map (
            O => \N__25712\,
            I => data_in_13_7
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__25709\,
            I => data_in_13_7
        );

    \I__5548\ : InMux
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__25696\,
            I => \N__25693\
        );

    \I__5545\ : Span4Mux_h
    port map (
            O => \N__25693\,
            I => \N__25688\
        );

    \I__5544\ : InMux
    port map (
            O => \N__25692\,
            I => \N__25683\
        );

    \I__5543\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25683\
        );

    \I__5542\ : Odrv4
    port map (
            O => \N__25688\,
            I => \c0.data_in_field_111\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__25683\,
            I => \c0.data_in_field_111\
        );

    \I__5540\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25673\
        );

    \I__5539\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25669\
        );

    \I__5538\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25665\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25662\
        );

    \I__5536\ : CascadeMux
    port map (
            O => \N__25672\,
            I => \N__25659\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25656\
        );

    \I__5534\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25653\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25649\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__25662\,
            I => \N__25646\
        );

    \I__5531\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25643\
        );

    \I__5530\ : Span12Mux_v
    port map (
            O => \N__25656\,
            I => \N__25640\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__25653\,
            I => \N__25637\
        );

    \I__5528\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25634\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__25649\,
            I => \N__25629\
        );

    \I__5526\ : Span4Mux_v
    port map (
            O => \N__25646\,
            I => \N__25629\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__25643\,
            I => \c0.data_in_field_143\
        );

    \I__5524\ : Odrv12
    port map (
            O => \N__25640\,
            I => \c0.data_in_field_143\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__25637\,
            I => \c0.data_in_field_143\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__25634\,
            I => \c0.data_in_field_143\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__25629\,
            I => \c0.data_in_field_143\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__25618\,
            I => \N__25615\
        );

    \I__5519\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25612\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__25612\,
            I => \N__25609\
        );

    \I__5517\ : Span4Mux_h
    port map (
            O => \N__25609\,
            I => \N__25605\
        );

    \I__5516\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25602\
        );

    \I__5515\ : Span4Mux_s0_v
    port map (
            O => \N__25605\,
            I => \N__25596\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__25602\,
            I => \N__25596\
        );

    \I__5513\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25593\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__25596\,
            I => data_in_16_7
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__25593\,
            I => data_in_16_7
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \N__25585\
        );

    \I__5509\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25582\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__25582\,
            I => \N__25579\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__25579\,
            I => \N__25574\
        );

    \I__5506\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25569\
        );

    \I__5505\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25569\
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__25574\,
            I => data_in_4_7
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__25569\,
            I => data_in_4_7
        );

    \I__5502\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25561\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__25561\,
            I => \N__25557\
        );

    \I__5500\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25554\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__25557\,
            I => \N__25549\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__25554\,
            I => \N__25546\
        );

    \I__5497\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25541\
        );

    \I__5496\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25541\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__25549\,
            I => \c0.data_in_field_39\
        );

    \I__5494\ : Odrv4
    port map (
            O => \N__25546\,
            I => \c0.data_in_field_39\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__25541\,
            I => \c0.data_in_field_39\
        );

    \I__5492\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25530\
        );

    \I__5491\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25527\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__25530\,
            I => \N__25523\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__25527\,
            I => \N__25520\
        );

    \I__5488\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25516\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__25523\,
            I => \N__25511\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__25520\,
            I => \N__25511\
        );

    \I__5485\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25508\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__25516\,
            I => \c0.data_in_field_5\
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__25511\,
            I => \c0.data_in_field_5\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__25508\,
            I => \c0.data_in_field_5\
        );

    \I__5481\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25498\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25494\
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__25497\,
            I => \N__25488\
        );

    \I__5478\ : Span4Mux_v
    port map (
            O => \N__25494\,
            I => \N__25485\
        );

    \I__5477\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25480\
        );

    \I__5476\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25480\
        );

    \I__5475\ : CascadeMux
    port map (
            O => \N__25491\,
            I => \N__25477\
        );

    \I__5474\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25474\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__25485\,
            I => \N__25469\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25469\
        );

    \I__5471\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25466\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__25474\,
            I => \c0.data_in_field_79\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__25469\,
            I => \c0.data_in_field_79\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__25466\,
            I => \c0.data_in_field_79\
        );

    \I__5467\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25456\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25453\
        );

    \I__5465\ : Span4Mux_s1_h
    port map (
            O => \N__25453\,
            I => \N__25448\
        );

    \I__5464\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25445\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__25451\,
            I => \N__25442\
        );

    \I__5462\ : Span4Mux_h
    port map (
            O => \N__25448\,
            I => \N__25439\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__25445\,
            I => \N__25436\
        );

    \I__5460\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25432\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__25439\,
            I => \N__25427\
        );

    \I__5458\ : Span4Mux_h
    port map (
            O => \N__25436\,
            I => \N__25427\
        );

    \I__5457\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25424\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__25432\,
            I => \c0.data_in_field_77\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__25427\,
            I => \c0.data_in_field_77\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__25424\,
            I => \c0.data_in_field_77\
        );

    \I__5453\ : CascadeMux
    port map (
            O => \N__25417\,
            I => \c0.n10_adj_1871_cascade_\
        );

    \I__5452\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25411\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__25411\,
            I => \N__25407\
        );

    \I__5450\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25404\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__25407\,
            I => \N__25399\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__25404\,
            I => \N__25399\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__25399\,
            I => \c0.n5234\
        );

    \I__5446\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__25393\,
            I => \N__25389\
        );

    \I__5444\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25386\
        );

    \I__5443\ : Odrv12
    port map (
            O => \N__25389\,
            I => \c0.n1975\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__25386\,
            I => \c0.n1975\
        );

    \I__5441\ : InMux
    port map (
            O => \N__25381\,
            I => \N__25378\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__25378\,
            I => \N__25374\
        );

    \I__5439\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25371\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__25374\,
            I => \N__25368\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__25371\,
            I => \N__25362\
        );

    \I__5436\ : Span4Mux_h
    port map (
            O => \N__25368\,
            I => \N__25359\
        );

    \I__5435\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25356\
        );

    \I__5434\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25351\
        );

    \I__5433\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25351\
        );

    \I__5432\ : Odrv12
    port map (
            O => \N__25362\,
            I => \c0.data_in_field_38\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__25359\,
            I => \c0.data_in_field_38\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__25356\,
            I => \c0.data_in_field_38\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__25351\,
            I => \c0.data_in_field_38\
        );

    \I__5428\ : InMux
    port map (
            O => \N__25342\,
            I => \N__25339\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__25339\,
            I => \N__25336\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__25336\,
            I => \N__25333\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__25333\,
            I => \N__25328\
        );

    \I__5424\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25325\
        );

    \I__5423\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25322\
        );

    \I__5422\ : Odrv4
    port map (
            O => \N__25328\,
            I => data_in_12_1
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__25325\,
            I => data_in_12_1
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__25322\,
            I => data_in_12_1
        );

    \I__5419\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25312\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__25312\,
            I => \N__25308\
        );

    \I__5417\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25305\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__25308\,
            I => \N__25302\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__25305\,
            I => \N__25299\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__25302\,
            I => \c0.n2062\
        );

    \I__5413\ : Odrv12
    port map (
            O => \N__25299\,
            I => \c0.n2062\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__25294\,
            I => \N__25289\
        );

    \I__5411\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25286\
        );

    \I__5410\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25283\
        );

    \I__5409\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25279\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25276\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__25283\,
            I => \N__25273\
        );

    \I__5406\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25270\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__25279\,
            I => \c0.data_in_field_61\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__25276\,
            I => \c0.data_in_field_61\
        );

    \I__5403\ : Odrv12
    port map (
            O => \N__25273\,
            I => \c0.data_in_field_61\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__25270\,
            I => \c0.data_in_field_61\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__25261\,
            I => \c0.n5875_cascade_\
        );

    \I__5400\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25255\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__25252\,
            I => \N__25246\
        );

    \I__5397\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25243\
        );

    \I__5396\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25240\
        );

    \I__5395\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25237\
        );

    \I__5394\ : Span4Mux_h
    port map (
            O => \N__25246\,
            I => \N__25234\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__25243\,
            I => \N__25231\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__25240\,
            I => \N__25228\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__25237\,
            I => \c0.data_in_field_37\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__25234\,
            I => \c0.data_in_field_37\
        );

    \I__5389\ : Odrv12
    port map (
            O => \N__25231\,
            I => \c0.data_in_field_37\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__25228\,
            I => \c0.data_in_field_37\
        );

    \I__5387\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25216\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__25213\,
            I => \N__25210\
        );

    \I__5384\ : Sp12to4
    port map (
            O => \N__25210\,
            I => \N__25207\
        );

    \I__5383\ : Span12Mux_s4_v
    port map (
            O => \N__25207\,
            I => \N__25204\
        );

    \I__5382\ : Odrv12
    port map (
            O => \N__25204\,
            I => \c0.n5396\
        );

    \I__5381\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25197\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__25200\,
            I => \N__25193\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__25197\,
            I => \N__25189\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__25196\,
            I => \N__25186\
        );

    \I__5377\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25182\
        );

    \I__5376\ : InMux
    port map (
            O => \N__25192\,
            I => \N__25179\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__25189\,
            I => \N__25176\
        );

    \I__5374\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25171\
        );

    \I__5373\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25171\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__25182\,
            I => \c0.data_in_field_53\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__25179\,
            I => \c0.data_in_field_53\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__25176\,
            I => \c0.data_in_field_53\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__25171\,
            I => \c0.data_in_field_53\
        );

    \I__5368\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25157\
        );

    \I__5367\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25154\
        );

    \I__5366\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25151\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25147\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__25154\,
            I => \N__25144\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__25151\,
            I => \N__25140\
        );

    \I__5362\ : InMux
    port map (
            O => \N__25150\,
            I => \N__25137\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__25147\,
            I => \N__25132\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__25144\,
            I => \N__25132\
        );

    \I__5359\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25129\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__25140\,
            I => \N__25126\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__25137\,
            I => \c0.data_in_field_88\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__25132\,
            I => \c0.data_in_field_88\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__25129\,
            I => \c0.data_in_field_88\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__25126\,
            I => \c0.data_in_field_88\
        );

    \I__5353\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25114\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__25114\,
            I => \N__25111\
        );

    \I__5351\ : Span4Mux_v
    port map (
            O => \N__25111\,
            I => \N__25108\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__25108\,
            I => \N__25101\
        );

    \I__5349\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25096\
        );

    \I__5348\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25096\
        );

    \I__5347\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25091\
        );

    \I__5346\ : InMux
    port map (
            O => \N__25104\,
            I => \N__25091\
        );

    \I__5345\ : Odrv4
    port map (
            O => \N__25101\,
            I => \c0.data_in_field_124\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__25096\,
            I => \c0.data_in_field_124\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__25091\,
            I => \c0.data_in_field_124\
        );

    \I__5342\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25077\
        );

    \I__5340\ : CascadeMux
    port map (
            O => \N__25080\,
            I => \N__25074\
        );

    \I__5339\ : Span4Mux_h
    port map (
            O => \N__25077\,
            I => \N__25071\
        );

    \I__5338\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25068\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__25071\,
            I => \c0.n1944\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__25068\,
            I => \c0.n1944\
        );

    \I__5335\ : CascadeMux
    port map (
            O => \N__25063\,
            I => \c0.n1944_cascade_\
        );

    \I__5334\ : CascadeMux
    port map (
            O => \N__25060\,
            I => \c0.n20_cascade_\
        );

    \I__5333\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25053\
        );

    \I__5332\ : InMux
    port map (
            O => \N__25056\,
            I => \N__25049\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__25053\,
            I => \N__25046\
        );

    \I__5330\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25043\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__25049\,
            I => \N__25040\
        );

    \I__5328\ : Span12Mux_s2_h
    port map (
            O => \N__25046\,
            I => \N__25033\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__25043\,
            I => \N__25033\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__25040\,
            I => \N__25030\
        );

    \I__5325\ : InMux
    port map (
            O => \N__25039\,
            I => \N__25025\
        );

    \I__5324\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25025\
        );

    \I__5323\ : Odrv12
    port map (
            O => \N__25033\,
            I => \c0.data_in_field_43\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__25030\,
            I => \c0.data_in_field_43\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__25025\,
            I => \c0.data_in_field_43\
        );

    \I__5320\ : InMux
    port map (
            O => \N__25018\,
            I => \N__25015\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__25015\,
            I => \N__25012\
        );

    \I__5318\ : Odrv12
    port map (
            O => \N__25012\,
            I => \c0.n24\
        );

    \I__5317\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25005\
        );

    \I__5316\ : CascadeMux
    port map (
            O => \N__25008\,
            I => \N__25000\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24997\
        );

    \I__5314\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24994\
        );

    \I__5313\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24991\
        );

    \I__5312\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24988\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__24997\,
            I => \N__24983\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__24994\,
            I => \N__24983\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__24991\,
            I => \N__24980\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__24988\,
            I => \c0.data_in_field_139\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__24983\,
            I => \c0.data_in_field_139\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__24980\,
            I => \c0.data_in_field_139\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__24973\,
            I => \c0.n1947_cascade_\
        );

    \I__5304\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24967\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__24967\,
            I => \c0.n10\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__5301\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24957\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__24960\,
            I => \N__24953\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__24957\,
            I => \N__24950\
        );

    \I__5298\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24947\
        );

    \I__5297\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24944\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__24950\,
            I => \N__24939\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24939\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__24944\,
            I => \N__24936\
        );

    \I__5293\ : Span4Mux_h
    port map (
            O => \N__24939\,
            I => \N__24933\
        );

    \I__5292\ : Span12Mux_s9_h
    port map (
            O => \N__24936\,
            I => \N__24928\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__24933\,
            I => \N__24925\
        );

    \I__5290\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24920\
        );

    \I__5289\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24920\
        );

    \I__5288\ : Odrv12
    port map (
            O => \N__24928\,
            I => \c0.data_in_field_51\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__24925\,
            I => \c0.data_in_field_51\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__24920\,
            I => \c0.data_in_field_51\
        );

    \I__5285\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__24910\,
            I => \N__24906\
        );

    \I__5283\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24903\
        );

    \I__5282\ : Odrv12
    port map (
            O => \N__24906\,
            I => \c0.n1922\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__24903\,
            I => \c0.n1922\
        );

    \I__5280\ : InMux
    port map (
            O => \N__24898\,
            I => \N__24895\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__24895\,
            I => \N__24891\
        );

    \I__5278\ : InMux
    port map (
            O => \N__24894\,
            I => \N__24888\
        );

    \I__5277\ : Span4Mux_h
    port map (
            O => \N__24891\,
            I => \N__24880\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__24888\,
            I => \N__24880\
        );

    \I__5275\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24877\
        );

    \I__5274\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24872\
        );

    \I__5273\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24872\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__24880\,
            I => \c0.data_in_field_75\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__24877\,
            I => \c0.data_in_field_75\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__24872\,
            I => \c0.data_in_field_75\
        );

    \I__5269\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24862\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__24862\,
            I => \N__24859\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__24859\,
            I => \N__24856\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__24856\,
            I => \c0.n5474\
        );

    \I__5265\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24850\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24847\
        );

    \I__5263\ : Span12Mux_s9_h
    port map (
            O => \N__24847\,
            I => \N__24844\
        );

    \I__5262\ : Odrv12
    port map (
            O => \N__24844\,
            I => \c0.n26_adj_1884\
        );

    \I__5261\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24837\
        );

    \I__5260\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24833\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24830\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__24836\,
            I => \N__24825\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24822\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__24830\,
            I => \N__24819\
        );

    \I__5255\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24816\
        );

    \I__5254\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24813\
        );

    \I__5253\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24810\
        );

    \I__5252\ : Span4Mux_v
    port map (
            O => \N__24822\,
            I => \N__24805\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__24819\,
            I => \N__24805\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__24816\,
            I => \N__24802\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__24813\,
            I => \c0.data_in_field_98\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__24810\,
            I => \c0.data_in_field_98\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__24805\,
            I => \c0.data_in_field_98\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__24802\,
            I => \c0.data_in_field_98\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__24793\,
            I => \N__24790\
        );

    \I__5244\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24786\
        );

    \I__5243\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24783\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24780\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__24783\,
            I => \N__24776\
        );

    \I__5240\ : Span4Mux_v
    port map (
            O => \N__24780\,
            I => \N__24773\
        );

    \I__5239\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24770\
        );

    \I__5238\ : Span4Mux_v
    port map (
            O => \N__24776\,
            I => \N__24767\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__24773\,
            I => \N__24764\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__24770\,
            I => data_in_12_7
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__24767\,
            I => data_in_12_7
        );

    \I__5234\ : Odrv4
    port map (
            O => \N__24764\,
            I => data_in_12_7
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__24757\,
            I => \N__24753\
        );

    \I__5232\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24750\
        );

    \I__5231\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24747\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24744\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24741\
        );

    \I__5228\ : Span4Mux_v
    port map (
            O => \N__24744\,
            I => \N__24736\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__24741\,
            I => \N__24733\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__24740\,
            I => \N__24730\
        );

    \I__5225\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24727\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__24736\,
            I => \N__24724\
        );

    \I__5223\ : Sp12to4
    port map (
            O => \N__24733\,
            I => \N__24721\
        );

    \I__5222\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24718\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__24727\,
            I => \c0.data_in_field_103\
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__24724\,
            I => \c0.data_in_field_103\
        );

    \I__5219\ : Odrv12
    port map (
            O => \N__24721\,
            I => \c0.data_in_field_103\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__24718\,
            I => \c0.data_in_field_103\
        );

    \I__5217\ : InMux
    port map (
            O => \N__24709\,
            I => \N__24706\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__24706\,
            I => \N__24703\
        );

    \I__5215\ : Span4Mux_v
    port map (
            O => \N__24703\,
            I => \N__24700\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__24700\,
            I => \N__24694\
        );

    \I__5213\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24687\
        );

    \I__5212\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24687\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24687\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__24694\,
            I => \c0.data_in_field_28\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__24687\,
            I => \c0.data_in_field_28\
        );

    \I__5208\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24679\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__24679\,
            I => \N__24676\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__24676\,
            I => \N__24672\
        );

    \I__5205\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24669\
        );

    \I__5204\ : Span4Mux_v
    port map (
            O => \N__24672\,
            I => \N__24665\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24662\
        );

    \I__5202\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24658\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__24665\,
            I => \N__24655\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__24662\,
            I => \N__24652\
        );

    \I__5199\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24649\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__24658\,
            I => \c0.data_in_field_20\
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__24655\,
            I => \c0.data_in_field_20\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__24652\,
            I => \c0.data_in_field_20\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__24649\,
            I => \c0.data_in_field_20\
        );

    \I__5194\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24636\
        );

    \I__5193\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24632\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__24636\,
            I => \N__24629\
        );

    \I__5191\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24626\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__24632\,
            I => \N__24623\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__24629\,
            I => \N__24618\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__24626\,
            I => \N__24618\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__24623\,
            I => \N__24613\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__24618\,
            I => \N__24610\
        );

    \I__5185\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24605\
        );

    \I__5184\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24605\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__24613\,
            I => \c0.data_in_field_12\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__24610\,
            I => \c0.data_in_field_12\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__24605\,
            I => \c0.data_in_field_12\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__24598\,
            I => \c0.n5851_cascade_\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__24595\,
            I => \N__24592\
        );

    \I__5178\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24589\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__24583\,
            I => \c0.n5408\
        );

    \I__5174\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24576\
        );

    \I__5173\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24573\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__24576\,
            I => \N__24570\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__24573\,
            I => \N__24567\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__24570\,
            I => \N__24564\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__24567\,
            I => \N__24561\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__24564\,
            I => \N__24558\
        );

    \I__5167\ : Span4Mux_v
    port map (
            O => \N__24561\,
            I => \N__24555\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__24558\,
            I => \c0.n5267\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__24555\,
            I => \c0.n5267\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__5163\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24544\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__24541\,
            I => \N__24538\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__24538\,
            I => \c0.n5905\
        );

    \I__5159\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24532\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__24532\,
            I => \c0.n2074\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__24529\,
            I => \N__24525\
        );

    \I__5156\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24521\
        );

    \I__5155\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24518\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__24524\,
            I => \N__24515\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24512\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24509\
        );

    \I__5151\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24506\
        );

    \I__5150\ : Span4Mux_v
    port map (
            O => \N__24512\,
            I => \N__24500\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__24509\,
            I => \N__24500\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24497\
        );

    \I__5147\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24494\
        );

    \I__5146\ : Sp12to4
    port map (
            O => \N__24500\,
            I => \N__24489\
        );

    \I__5145\ : Span12Mux_h
    port map (
            O => \N__24497\,
            I => \N__24489\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__24494\,
            I => data_in_19_5
        );

    \I__5143\ : Odrv12
    port map (
            O => \N__24489\,
            I => data_in_19_5
        );

    \I__5142\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__5140\ : Odrv12
    port map (
            O => \N__24478\,
            I => \c0.n22_adj_1914\
        );

    \I__5139\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24471\
        );

    \I__5138\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24468\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__24471\,
            I => \N__24465\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__24468\,
            I => \N__24462\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__24465\,
            I => \N__24458\
        );

    \I__5134\ : Span4Mux_s2_v
    port map (
            O => \N__24462\,
            I => \N__24455\
        );

    \I__5133\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24452\
        );

    \I__5132\ : Span4Mux_h
    port map (
            O => \N__24458\,
            I => \N__24447\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__24455\,
            I => \N__24447\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__24452\,
            I => data_in_16_5
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__24447\,
            I => data_in_16_5
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__5127\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24436\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__24436\,
            I => \N__24431\
        );

    \I__5125\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24428\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__24434\,
            I => \N__24425\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__24431\,
            I => \N__24420\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__24428\,
            I => \N__24420\
        );

    \I__5121\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24417\
        );

    \I__5120\ : Span4Mux_h
    port map (
            O => \N__24420\,
            I => \N__24413\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__24417\,
            I => \N__24410\
        );

    \I__5118\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24407\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__24413\,
            I => \N__24404\
        );

    \I__5116\ : Span12Mux_s5_h
    port map (
            O => \N__24410\,
            I => \N__24401\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__24407\,
            I => data_in_19_2
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__24404\,
            I => data_in_19_2
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__24401\,
            I => data_in_19_2
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__5111\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24388\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__5109\ : Odrv4
    port map (
            O => \N__24385\,
            I => \c0.n5779\
        );

    \I__5108\ : InMux
    port map (
            O => \N__24382\,
            I => \N__24376\
        );

    \I__5107\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24376\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24372\
        );

    \I__5105\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24369\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__24372\,
            I => data_in_13_0
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__24369\,
            I => data_in_13_0
        );

    \I__5102\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24358\
        );

    \I__5101\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24358\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__5098\ : Span4Mux_h
    port map (
            O => \N__24352\,
            I => \N__24348\
        );

    \I__5097\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24345\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__24348\,
            I => data_in_14_0
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__24345\,
            I => data_in_14_0
        );

    \I__5094\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24337\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__24337\,
            I => \N__24334\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__24334\,
            I => \N__24331\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__24331\,
            I => \c0.n1929\
        );

    \I__5090\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24324\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__24327\,
            I => \N__24320\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__24324\,
            I => \N__24317\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \N__24313\
        );

    \I__5086\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24310\
        );

    \I__5085\ : Span4Mux_v
    port map (
            O => \N__24317\,
            I => \N__24307\
        );

    \I__5084\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24304\
        );

    \I__5083\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24301\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__24310\,
            I => \N__24298\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__24307\,
            I => \N__24293\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__24304\,
            I => \N__24293\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__24301\,
            I => \c0.data_in_field_112\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__24298\,
            I => \c0.data_in_field_112\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__24293\,
            I => \c0.data_in_field_112\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__24286\,
            I => \c0.n1929_cascade_\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__24283\,
            I => \c0.n10_adj_1870_cascade_\
        );

    \I__5074\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24276\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__24279\,
            I => \N__24273\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24270\
        );

    \I__5071\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24267\
        );

    \I__5070\ : Span4Mux_v
    port map (
            O => \N__24270\,
            I => \N__24264\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24261\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__24264\,
            I => \N__24258\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__24261\,
            I => \N__24255\
        );

    \I__5066\ : Odrv4
    port map (
            O => \N__24258\,
            I => \c0.n5204\
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__24255\,
            I => \c0.n5204\
        );

    \I__5064\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24243\
        );

    \I__5062\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24240\
        );

    \I__5061\ : Span4Mux_s2_v
    port map (
            O => \N__24243\,
            I => \N__24235\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24235\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__24235\,
            I => \N__24231\
        );

    \I__5058\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24228\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__24231\,
            I => data_in_7_5
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__24228\,
            I => data_in_7_5
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__24223\,
            I => \N__24219\
        );

    \I__5054\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24216\
        );

    \I__5053\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24213\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__24216\,
            I => \N__24208\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__24213\,
            I => \N__24205\
        );

    \I__5050\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24202\
        );

    \I__5049\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24199\
        );

    \I__5048\ : Span12Mux_s2_v
    port map (
            O => \N__24208\,
            I => \N__24196\
        );

    \I__5047\ : Span4Mux_v
    port map (
            O => \N__24205\,
            I => \N__24193\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__24202\,
            I => data_in_18_6
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__24199\,
            I => data_in_18_6
        );

    \I__5044\ : Odrv12
    port map (
            O => \N__24196\,
            I => data_in_18_6
        );

    \I__5043\ : Odrv4
    port map (
            O => \N__24193\,
            I => data_in_18_6
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__24184\,
            I => \N__24180\
        );

    \I__5041\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24177\
        );

    \I__5040\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24174\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__24177\,
            I => \N__24171\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24167\
        );

    \I__5037\ : Span4Mux_h
    port map (
            O => \N__24171\,
            I => \N__24164\
        );

    \I__5036\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24161\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__24167\,
            I => data_in_17_6
        );

    \I__5034\ : Odrv4
    port map (
            O => \N__24164\,
            I => data_in_17_6
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__24161\,
            I => data_in_17_6
        );

    \I__5032\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24151\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__24151\,
            I => \N__24147\
        );

    \I__5030\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24143\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__24147\,
            I => \N__24140\
        );

    \I__5028\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24136\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__24143\,
            I => \N__24133\
        );

    \I__5026\ : Sp12to4
    port map (
            O => \N__24140\,
            I => \N__24130\
        );

    \I__5025\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24127\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__24136\,
            I => data_in_1_5
        );

    \I__5023\ : Odrv12
    port map (
            O => \N__24133\,
            I => data_in_1_5
        );

    \I__5022\ : Odrv12
    port map (
            O => \N__24130\,
            I => data_in_1_5
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__24127\,
            I => data_in_1_5
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__24118\,
            I => \N__24115\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24111\
        );

    \I__5018\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24108\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__24111\,
            I => \N__24105\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24102\
        );

    \I__5015\ : Span4Mux_v
    port map (
            O => \N__24105\,
            I => \N__24098\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__24102\,
            I => \N__24095\
        );

    \I__5013\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24092\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__24098\,
            I => data_in_7_7
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__24095\,
            I => data_in_7_7
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__24092\,
            I => data_in_7_7
        );

    \I__5009\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24082\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__24082\,
            I => \N__24078\
        );

    \I__5007\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24075\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__24078\,
            I => \N__24072\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__24069\
        );

    \I__5004\ : Sp12to4
    port map (
            O => \N__24072\,
            I => \N__24062\
        );

    \I__5003\ : Span12Mux_v
    port map (
            O => \N__24069\,
            I => \N__24062\
        );

    \I__5002\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24057\
        );

    \I__5001\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24057\
        );

    \I__5000\ : Odrv12
    port map (
            O => \N__24062\,
            I => \c0.data_in_field_121\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__24057\,
            I => \c0.data_in_field_121\
        );

    \I__4998\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24049\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24044\
        );

    \I__4996\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24040\
        );

    \I__4995\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24037\
        );

    \I__4994\ : Span4Mux_h
    port map (
            O => \N__24044\,
            I => \N__24034\
        );

    \I__4993\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24031\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__24040\,
            I => \N__24026\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__24037\,
            I => \N__24026\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__24034\,
            I => data_in_3_7
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__24031\,
            I => data_in_3_7
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__24026\,
            I => data_in_3_7
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__4986\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24012\
        );

    \I__4985\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24009\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__24012\,
            I => \N__24004\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__24009\,
            I => \N__24004\
        );

    \I__4982\ : Span4Mux_s3_v
    port map (
            O => \N__24004\,
            I => \N__24000\
        );

    \I__4981\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23997\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__24000\,
            I => \N__23994\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__23997\,
            I => \N__23991\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__23994\,
            I => data_in_17_5
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__23991\,
            I => data_in_17_5
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__23986\,
            I => \N__23983\
        );

    \I__4975\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23980\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__23980\,
            I => \N__23976\
        );

    \I__4973\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23973\
        );

    \I__4972\ : Span4Mux_h
    port map (
            O => \N__23976\,
            I => \N__23969\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N__23966\
        );

    \I__4970\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23963\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__23969\,
            I => data_in_7_1
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__23966\,
            I => data_in_7_1
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__23963\,
            I => data_in_7_1
        );

    \I__4966\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23953\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__4964\ : Span4Mux_s2_v
    port map (
            O => \N__23950\,
            I => \N__23945\
        );

    \I__4963\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23940\
        );

    \I__4962\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23940\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__23945\,
            I => \N__23937\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__23940\,
            I => data_in_6_1
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__23937\,
            I => data_in_6_1
        );

    \I__4958\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23929\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23925\
        );

    \I__4956\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23922\
        );

    \I__4955\ : Span4Mux_h
    port map (
            O => \N__23925\,
            I => \N__23915\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23915\
        );

    \I__4953\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23912\
        );

    \I__4952\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23908\
        );

    \I__4951\ : Span4Mux_v
    port map (
            O => \N__23915\,
            I => \N__23903\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23903\
        );

    \I__4949\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23900\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__23908\,
            I => \c0.data_in_field_141\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__23903\,
            I => \c0.data_in_field_141\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__23900\,
            I => \c0.data_in_field_141\
        );

    \I__4945\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23888\
        );

    \I__4944\ : InMux
    port map (
            O => \N__23892\,
            I => \N__23885\
        );

    \I__4943\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23882\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23879\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__23885\,
            I => \N__23876\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23873\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__23879\,
            I => \N__23868\
        );

    \I__4938\ : Span4Mux_s2_v
    port map (
            O => \N__23876\,
            I => \N__23868\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__23873\,
            I => \N__23865\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__23868\,
            I => \N__23861\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__23865\,
            I => \N__23858\
        );

    \I__4934\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23855\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__23861\,
            I => \N__23852\
        );

    \I__4932\ : Odrv4
    port map (
            O => \N__23858\,
            I => data_in_1_6
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__23855\,
            I => data_in_1_6
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__23852\,
            I => data_in_1_6
        );

    \I__4929\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23841\
        );

    \I__4928\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23838\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__23841\,
            I => \N__23835\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__23838\,
            I => \N__23832\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__23835\,
            I => \N__23829\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__23832\,
            I => \N__23825\
        );

    \I__4923\ : Span4Mux_s0_v
    port map (
            O => \N__23829\,
            I => \N__23822\
        );

    \I__4922\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23819\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__23825\,
            I => data_in_9_7
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__23822\,
            I => data_in_9_7
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__23819\,
            I => data_in_9_7
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__23812\,
            I => \N__23809\
        );

    \I__4917\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__4915\ : Span12Mux_v
    port map (
            O => \N__23803\,
            I => \N__23798\
        );

    \I__4914\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23793\
        );

    \I__4913\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23793\
        );

    \I__4912\ : Odrv12
    port map (
            O => \N__23798\,
            I => data_in_6_7
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__23793\,
            I => data_in_6_7
        );

    \I__4910\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23784\
        );

    \I__4909\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23781\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23778\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__23781\,
            I => \N__23775\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__23778\,
            I => \N__23768\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__23775\,
            I => \N__23768\
        );

    \I__4904\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23763\
        );

    \I__4903\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23763\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__23768\,
            I => data_in_3_1
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__23763\,
            I => data_in_3_1
        );

    \I__4900\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23754\
        );

    \I__4899\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23751\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__23754\,
            I => \N__23747\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__23751\,
            I => \N__23744\
        );

    \I__4896\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23741\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__23747\,
            I => \N__23736\
        );

    \I__4894\ : Span4Mux_h
    port map (
            O => \N__23744\,
            I => \N__23731\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__23741\,
            I => \N__23731\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__23740\,
            I => \N__23728\
        );

    \I__4891\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23725\
        );

    \I__4890\ : Span4Mux_h
    port map (
            O => \N__23736\,
            I => \N__23722\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__23731\,
            I => \N__23719\
        );

    \I__4888\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23716\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__23725\,
            I => \c0.data_in_field_21\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__23722\,
            I => \c0.data_in_field_21\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__23719\,
            I => \c0.data_in_field_21\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__23716\,
            I => \c0.data_in_field_21\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__23707\,
            I => \N__23704\
        );

    \I__4882\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23701\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__23701\,
            I => \N__23698\
        );

    \I__4880\ : Span12Mux_s8_h
    port map (
            O => \N__23698\,
            I => \N__23695\
        );

    \I__4879\ : Odrv12
    port map (
            O => \N__23695\,
            I => \c0.n5881\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23688\
        );

    \I__4877\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23685\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__23688\,
            I => \N__23682\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23679\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__23682\,
            I => \N__23676\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__23679\,
            I => \N__23673\
        );

    \I__4872\ : Span4Mux_s2_v
    port map (
            O => \N__23676\,
            I => \N__23669\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__23673\,
            I => \N__23666\
        );

    \I__4870\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23663\
        );

    \I__4869\ : Odrv4
    port map (
            O => \N__23669\,
            I => data_in_15_6
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__23666\,
            I => data_in_15_6
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__23663\,
            I => data_in_15_6
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__23656\,
            I => \N__23653\
        );

    \I__4865\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23648\
        );

    \I__4864\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23643\
        );

    \I__4863\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23643\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__23648\,
            I => \c0.data_in_field_29\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__23643\,
            I => \c0.data_in_field_29\
        );

    \I__4860\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__23635\,
            I => \N__23632\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__23632\,
            I => \N__23629\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__23626\,
            I => \c0.n2046\
        );

    \I__4855\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23620\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__23620\,
            I => \N__23615\
        );

    \I__4853\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23612\
        );

    \I__4852\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23609\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__23615\,
            I => \N__23604\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23604\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23601\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__23604\,
            I => \N__23597\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__23601\,
            I => \N__23594\
        );

    \I__4846\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23591\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__23597\,
            I => \N__23588\
        );

    \I__4844\ : Span4Mux_h
    port map (
            O => \N__23594\,
            I => \N__23585\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__23591\,
            I => \c0.data_in_field_85\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__23588\,
            I => \c0.data_in_field_85\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__23585\,
            I => \c0.data_in_field_85\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__23578\,
            I => \c0.n2046_cascade_\
        );

    \I__4839\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23572\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__23572\,
            I => \N__23568\
        );

    \I__4837\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23565\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__23568\,
            I => \N__23562\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23559\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__23562\,
            I => \c0.n5108\
        );

    \I__4833\ : Odrv12
    port map (
            O => \N__23559\,
            I => \c0.n5108\
        );

    \I__4832\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23550\
        );

    \I__4831\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23547\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23543\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23540\
        );

    \I__4828\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23536\
        );

    \I__4827\ : Span4Mux_h
    port map (
            O => \N__23543\,
            I => \N__23532\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__23540\,
            I => \N__23529\
        );

    \I__4825\ : InMux
    port map (
            O => \N__23539\,
            I => \N__23526\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__23536\,
            I => \N__23523\
        );

    \I__4823\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23520\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__23532\,
            I => \N__23517\
        );

    \I__4821\ : Span4Mux_h
    port map (
            O => \N__23529\,
            I => \N__23512\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__23526\,
            I => \N__23512\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__23523\,
            I => \N__23509\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__23520\,
            I => \c0.data_in_field_89\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__23517\,
            I => \c0.data_in_field_89\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__23512\,
            I => \c0.data_in_field_89\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__23509\,
            I => \c0.data_in_field_89\
        );

    \I__4814\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23496\
        );

    \I__4813\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23493\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__23496\,
            I => \N__23488\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__23493\,
            I => \N__23485\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23482\
        );

    \I__4809\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23479\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__23488\,
            I => \N__23472\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__23485\,
            I => \N__23472\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23472\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23469\
        );

    \I__4804\ : Span4Mux_h
    port map (
            O => \N__23472\,
            I => \N__23464\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__23469\,
            I => \N__23461\
        );

    \I__4802\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23456\
        );

    \I__4801\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23456\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__23464\,
            I => \c0.data_in_field_120\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__23461\,
            I => \c0.data_in_field_120\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__23456\,
            I => \c0.data_in_field_120\
        );

    \I__4797\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23446\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__23446\,
            I => \N__23443\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__23443\,
            I => \N__23440\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__23440\,
            I => \c0.n23_adj_1925\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__23437\,
            I => \N__23433\
        );

    \I__4792\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23429\
        );

    \I__4791\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23426\
        );

    \I__4790\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23423\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__23429\,
            I => \N__23419\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__23426\,
            I => \N__23416\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23413\
        );

    \I__4786\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23410\
        );

    \I__4785\ : Span12Mux_h
    port map (
            O => \N__23419\,
            I => \N__23407\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__23416\,
            I => \N__23404\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__23413\,
            I => \N__23401\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__23410\,
            I => \c0.data_in_field_83\
        );

    \I__4781\ : Odrv12
    port map (
            O => \N__23407\,
            I => \c0.data_in_field_83\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__23404\,
            I => \c0.data_in_field_83\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__23401\,
            I => \c0.data_in_field_83\
        );

    \I__4778\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23389\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__23389\,
            I => \N__23386\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__23383\,
            I => \c0.n5797\
        );

    \I__4774\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23376\
        );

    \I__4773\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23373\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__23376\,
            I => \N__23369\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__23373\,
            I => \N__23366\
        );

    \I__4770\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23363\
        );

    \I__4769\ : Span4Mux_v
    port map (
            O => \N__23369\,
            I => \N__23358\
        );

    \I__4768\ : Span4Mux_h
    port map (
            O => \N__23366\,
            I => \N__23358\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__23363\,
            I => \N__23355\
        );

    \I__4766\ : Span4Mux_h
    port map (
            O => \N__23358\,
            I => \N__23350\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__23355\,
            I => \N__23347\
        );

    \I__4764\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23342\
        );

    \I__4763\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23342\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__23350\,
            I => \c0.data_in_field_19\
        );

    \I__4761\ : Odrv4
    port map (
            O => \N__23347\,
            I => \c0.data_in_field_19\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__23342\,
            I => \c0.data_in_field_19\
        );

    \I__4759\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23332\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__23332\,
            I => \N__23329\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__23329\,
            I => \N__23326\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__23326\,
            I => \c0.n23\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__23323\,
            I => \N__23320\
        );

    \I__4754\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23316\
        );

    \I__4753\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23313\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__23316\,
            I => \N__23309\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23306\
        );

    \I__4750\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23302\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__23309\,
            I => \N__23299\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__23306\,
            I => \N__23296\
        );

    \I__4747\ : InMux
    port map (
            O => \N__23305\,
            I => \N__23293\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__23302\,
            I => \N__23290\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__23299\,
            I => \N__23287\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__23296\,
            I => \N__23284\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__23293\,
            I => data_in_3_3
        );

    \I__4742\ : Odrv12
    port map (
            O => \N__23290\,
            I => data_in_3_3
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__23287\,
            I => data_in_3_3
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__23284\,
            I => data_in_3_3
        );

    \I__4739\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23272\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__23272\,
            I => \N__23269\
        );

    \I__4737\ : Span4Mux_s2_v
    port map (
            O => \N__23269\,
            I => \N__23266\
        );

    \I__4736\ : Span4Mux_h
    port map (
            O => \N__23266\,
            I => \N__23263\
        );

    \I__4735\ : Odrv4
    port map (
            O => \N__23263\,
            I => \c0.n25_adj_1960\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__23260\,
            I => \N__23257\
        );

    \I__4733\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23252\
        );

    \I__4732\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23249\
        );

    \I__4731\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23245\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__23252\,
            I => \N__23240\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__23249\,
            I => \N__23240\
        );

    \I__4728\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23236\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23233\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__23240\,
            I => \N__23230\
        );

    \I__4725\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23227\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23222\
        );

    \I__4723\ : Span4Mux_h
    port map (
            O => \N__23233\,
            I => \N__23222\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__23230\,
            I => \c0.data_in_field_67\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__23227\,
            I => \c0.data_in_field_67\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__23222\,
            I => \c0.data_in_field_67\
        );

    \I__4719\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23208\
        );

    \I__4717\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23205\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__23208\,
            I => \N__23202\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__23205\,
            I => \N__23199\
        );

    \I__4714\ : Span4Mux_v
    port map (
            O => \N__23202\,
            I => \N__23194\
        );

    \I__4713\ : Span4Mux_v
    port map (
            O => \N__23199\,
            I => \N__23194\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__23194\,
            I => \c0.n5093\
        );

    \I__4711\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23188\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__4709\ : Span4Mux_h
    port map (
            O => \N__23185\,
            I => \N__23182\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__23182\,
            I => \c0.n5162\
        );

    \I__4707\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23172\
        );

    \I__4705\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23169\
        );

    \I__4704\ : Odrv12
    port map (
            O => \N__23172\,
            I => \c0.n5213\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__23169\,
            I => \c0.n5213\
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__23164\,
            I => \c0.n5099_cascade_\
        );

    \I__4701\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23158\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__23158\,
            I => \N__23155\
        );

    \I__4699\ : Span4Mux_h
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__23152\,
            I => \c0.n19\
        );

    \I__4697\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23145\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__23148\,
            I => \N__23142\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23139\
        );

    \I__4694\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23135\
        );

    \I__4693\ : Span4Mux_h
    port map (
            O => \N__23139\,
            I => \N__23132\
        );

    \I__4692\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23129\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__23135\,
            I => \c0.data_in_field_104\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__23132\,
            I => \c0.data_in_field_104\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__23129\,
            I => \c0.data_in_field_104\
        );

    \I__4688\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__23116\,
            I => \N__23113\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__23113\,
            I => \N__23108\
        );

    \I__4684\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23103\
        );

    \I__4683\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23103\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__23108\,
            I => data_in_0_6
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__23103\,
            I => data_in_0_6
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__4679\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23090\
        );

    \I__4678\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23085\
        );

    \I__4677\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23085\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__23090\,
            I => data_in_12_0
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__23085\,
            I => data_in_12_0
        );

    \I__4674\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__23071\,
            I => \c0.n13\
        );

    \I__4670\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23064\
        );

    \I__4669\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23061\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23058\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__23061\,
            I => \N__23055\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__23058\,
            I => \N__23051\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__23055\,
            I => \N__23048\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23044\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__23051\,
            I => \N__23041\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__23048\,
            I => \N__23038\
        );

    \I__4661\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23033\
        );

    \I__4660\ : InMux
    port map (
            O => \N__23044\,
            I => \N__23033\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__23041\,
            I => \c0.data_in_field_117\
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__23038\,
            I => \c0.data_in_field_117\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__23033\,
            I => \c0.data_in_field_117\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__23026\,
            I => \c0.n2074_cascade_\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__23023\,
            I => \N__23020\
        );

    \I__4654\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23017\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__23014\,
            I => \N__23011\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__23011\,
            I => \c0.n10_adj_1888\
        );

    \I__4650\ : InMux
    port map (
            O => \N__23008\,
            I => \N__23004\
        );

    \I__4649\ : InMux
    port map (
            O => \N__23007\,
            I => \N__23001\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__23004\,
            I => \N__22998\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22992\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__22998\,
            I => \N__22989\
        );

    \I__4645\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22982\
        );

    \I__4644\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22982\
        );

    \I__4643\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22982\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__22992\,
            I => \c0.data_in_field_95\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__22989\,
            I => \c0.data_in_field_95\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__22982\,
            I => \c0.data_in_field_95\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__22972\,
            I => \N__22968\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__22971\,
            I => \N__22965\
        );

    \I__4636\ : Span4Mux_h
    port map (
            O => \N__22968\,
            I => \N__22962\
        );

    \I__4635\ : InMux
    port map (
            O => \N__22965\,
            I => \N__22959\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__22962\,
            I => \c0.n1851\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__22959\,
            I => \c0.n1851\
        );

    \I__4632\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__22951\,
            I => \N__22947\
        );

    \I__4630\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22943\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__22947\,
            I => \N__22940\
        );

    \I__4628\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22937\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__22943\,
            I => \N__22933\
        );

    \I__4626\ : Sp12to4
    port map (
            O => \N__22940\,
            I => \N__22928\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__22937\,
            I => \N__22928\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__22936\,
            I => \N__22922\
        );

    \I__4623\ : Span4Mux_v
    port map (
            O => \N__22933\,
            I => \N__22919\
        );

    \I__4622\ : Span12Mux_s7_v
    port map (
            O => \N__22928\,
            I => \N__22916\
        );

    \I__4621\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22911\
        );

    \I__4620\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22911\
        );

    \I__4619\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22906\
        );

    \I__4618\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22906\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__22919\,
            I => \c0.data_in_field_96\
        );

    \I__4616\ : Odrv12
    port map (
            O => \N__22916\,
            I => \c0.data_in_field_96\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__22911\,
            I => \c0.data_in_field_96\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__22906\,
            I => \c0.data_in_field_96\
        );

    \I__4613\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__4611\ : Odrv12
    port map (
            O => \N__22891\,
            I => \c0.n5099\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__22888\,
            I => \c0.n5447_cascade_\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__22885\,
            I => \c0.n5755_cascade_\
        );

    \I__4608\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__4606\ : Span12Mux_s9_v
    port map (
            O => \N__22876\,
            I => \N__22873\
        );

    \I__4605\ : Odrv12
    port map (
            O => \N__22873\,
            I => \c0.n5758\
        );

    \I__4604\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22866\
        );

    \I__4603\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22861\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22858\
        );

    \I__4601\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22855\
        );

    \I__4600\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22852\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__22861\,
            I => \N__22849\
        );

    \I__4598\ : Span12Mux_s5_h
    port map (
            O => \N__22858\,
            I => \N__22846\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22843\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__22852\,
            I => \c0.data_in_field_54\
        );

    \I__4595\ : Odrv12
    port map (
            O => \N__22849\,
            I => \c0.data_in_field_54\
        );

    \I__4594\ : Odrv12
    port map (
            O => \N__22846\,
            I => \c0.data_in_field_54\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__22843\,
            I => \c0.data_in_field_54\
        );

    \I__4592\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22831\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__22831\,
            I => \N__22827\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22824\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__22827\,
            I => \N__22818\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22815\
        );

    \I__4587\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22812\
        );

    \I__4586\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22807\
        );

    \I__4585\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22807\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__22818\,
            I => \N__22800\
        );

    \I__4583\ : Span4Mux_v
    port map (
            O => \N__22815\,
            I => \N__22800\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22800\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__22807\,
            I => \c0.data_in_field_10\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__22800\,
            I => \c0.data_in_field_10\
        );

    \I__4579\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__22792\,
            I => \c0.n5438\
        );

    \I__4577\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22786\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__22786\,
            I => \N__22782\
        );

    \I__4575\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22779\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__22782\,
            I => \N__22773\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__22779\,
            I => \N__22773\
        );

    \I__4572\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22770\
        );

    \I__4571\ : Span4Mux_v
    port map (
            O => \N__22773\,
            I => \N__22763\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__22770\,
            I => \N__22763\
        );

    \I__4569\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22758\
        );

    \I__4568\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22758\
        );

    \I__4567\ : Span4Mux_h
    port map (
            O => \N__22763\,
            I => \N__22755\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__22758\,
            I => \c0.data_in_field_82\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__22755\,
            I => \c0.data_in_field_82\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__22750\,
            I => \c0.n5767_cascade_\
        );

    \I__4563\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__22744\,
            I => \c0.n5444\
        );

    \I__4561\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22738\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__22738\,
            I => \c0.n5761\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__22735\,
            I => \N__22731\
        );

    \I__4558\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22728\
        );

    \I__4557\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22725\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22722\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__22725\,
            I => \N__22718\
        );

    \I__4554\ : Span4Mux_h
    port map (
            O => \N__22722\,
            I => \N__22715\
        );

    \I__4553\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22712\
        );

    \I__4552\ : Odrv12
    port map (
            O => \N__22718\,
            I => data_in_11_7
        );

    \I__4551\ : Odrv4
    port map (
            O => \N__22715\,
            I => data_in_11_7
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__22712\,
            I => data_in_11_7
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__22705\,
            I => \N__22702\
        );

    \I__4548\ : InMux
    port map (
            O => \N__22702\,
            I => \N__22699\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__22699\,
            I => \N__22696\
        );

    \I__4546\ : Span4Mux_h
    port map (
            O => \N__22696\,
            I => \N__22691\
        );

    \I__4545\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22688\
        );

    \I__4544\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22685\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__22691\,
            I => data_in_10_7
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__22688\,
            I => data_in_10_7
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__22685\,
            I => data_in_10_7
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__22678\,
            I => \N__22675\
        );

    \I__4539\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22672\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__22672\,
            I => \N__22667\
        );

    \I__4537\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22664\
        );

    \I__4536\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22660\
        );

    \I__4535\ : Span4Mux_v
    port map (
            O => \N__22667\,
            I => \N__22655\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__22664\,
            I => \N__22655\
        );

    \I__4533\ : InMux
    port map (
            O => \N__22663\,
            I => \N__22652\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__22660\,
            I => data_in_2_7
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__22655\,
            I => data_in_2_7
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__22652\,
            I => data_in_2_7
        );

    \I__4529\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22642\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__22642\,
            I => \c0.n27_adj_1956\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__4526\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22633\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__22633\,
            I => \N__22630\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__22630\,
            I => \c0.n26_adj_1958\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22624\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22619\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__22623\,
            I => \N__22616\
        );

    \I__4520\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22613\
        );

    \I__4519\ : Span4Mux_s1_h
    port map (
            O => \N__22619\,
            I => \N__22610\
        );

    \I__4518\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22607\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22604\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__22610\,
            I => \N__22598\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__22607\,
            I => \N__22598\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__22604\,
            I => \N__22594\
        );

    \I__4513\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22591\
        );

    \I__4512\ : Sp12to4
    port map (
            O => \N__22598\,
            I => \N__22588\
        );

    \I__4511\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22585\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__22594\,
            I => \N__22582\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__22591\,
            I => \c0.data_in_field_135\
        );

    \I__4508\ : Odrv12
    port map (
            O => \N__22588\,
            I => \c0.data_in_field_135\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__22585\,
            I => \c0.data_in_field_135\
        );

    \I__4506\ : Odrv4
    port map (
            O => \N__22582\,
            I => \c0.data_in_field_135\
        );

    \I__4505\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22568\
        );

    \I__4504\ : CascadeMux
    port map (
            O => \N__22572\,
            I => \N__22564\
        );

    \I__4503\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22561\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__22568\,
            I => \N__22558\
        );

    \I__4501\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22555\
        );

    \I__4500\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22552\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__22561\,
            I => \N__22549\
        );

    \I__4498\ : Span4Mux_v
    port map (
            O => \N__22558\,
            I => \N__22546\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__22555\,
            I => \N__22541\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__22552\,
            I => \N__22541\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__22549\,
            I => \c0.data_in_field_113\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__22546\,
            I => \c0.data_in_field_113\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__22541\,
            I => \c0.data_in_field_113\
        );

    \I__4492\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22530\
        );

    \I__4491\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22527\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__22530\,
            I => \c0.n1772\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__22527\,
            I => \c0.n1772\
        );

    \I__4488\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__4486\ : Span4Mux_v
    port map (
            O => \N__22516\,
            I => \N__22513\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__22513\,
            I => \N__22510\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__22510\,
            I => \c0.n5144\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__22507\,
            I => \c0.n5144_cascade_\
        );

    \I__4482\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__22501\,
            I => \c0.n31\
        );

    \I__4480\ : CascadeMux
    port map (
            O => \N__22498\,
            I => \N__22494\
        );

    \I__4479\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22491\
        );

    \I__4478\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22488\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22485\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22481\
        );

    \I__4475\ : Span4Mux_h
    port map (
            O => \N__22485\,
            I => \N__22478\
        );

    \I__4474\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22475\
        );

    \I__4473\ : Odrv12
    port map (
            O => \N__22481\,
            I => data_in_8_5
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__22478\,
            I => data_in_8_5
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__22475\,
            I => data_in_8_5
        );

    \I__4470\ : InMux
    port map (
            O => \N__22468\,
            I => \N__22465\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__22465\,
            I => \N__22461\
        );

    \I__4468\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22458\
        );

    \I__4467\ : Span4Mux_v
    port map (
            O => \N__22461\,
            I => \N__22454\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22451\
        );

    \I__4465\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22448\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__22454\,
            I => data_in_8_7
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__22451\,
            I => data_in_8_7
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__22448\,
            I => data_in_8_7
        );

    \I__4461\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22434\
        );

    \I__4459\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22431\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__22434\,
            I => \N__22426\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22426\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__22426\,
            I => \c0.n5249\
        );

    \I__4455\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22417\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__22417\,
            I => \N__22413\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__22416\,
            I => \N__22410\
        );

    \I__4451\ : Span4Mux_s0_v
    port map (
            O => \N__22413\,
            I => \N__22407\
        );

    \I__4450\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22404\
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__22407\,
            I => rx_data_2
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__22404\,
            I => rx_data_2
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__4446\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22393\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__22390\,
            I => \N__22386\
        );

    \I__4443\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22383\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__22386\,
            I => \N__22380\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__22383\,
            I => \c0.n5255\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__22380\,
            I => \c0.n5255\
        );

    \I__4439\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22372\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22368\
        );

    \I__4437\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22365\
        );

    \I__4436\ : Span4Mux_s3_h
    port map (
            O => \N__22368\,
            I => \N__22358\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22358\
        );

    \I__4434\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22355\
        );

    \I__4433\ : InMux
    port map (
            O => \N__22363\,
            I => \N__22352\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__22358\,
            I => \N__22347\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__22355\,
            I => \N__22347\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__22352\,
            I => data_in_1_3
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__22347\,
            I => data_in_1_3
        );

    \I__4428\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__22336\,
            I => \c0.n28_adj_1954\
        );

    \I__4425\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22330\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__4423\ : Odrv12
    port map (
            O => \N__22327\,
            I => \c0.n26_adj_1955\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__22324\,
            I => \c0.n25_adj_1957_cascade_\
        );

    \I__4421\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__22318\,
            I => \c0.n4465\
        );

    \I__4419\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22312\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__22312\,
            I => \N__22309\
        );

    \I__4417\ : Span4Mux_h
    port map (
            O => \N__22309\,
            I => \N__22304\
        );

    \I__4416\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22300\
        );

    \I__4415\ : InMux
    port map (
            O => \N__22307\,
            I => \N__22297\
        );

    \I__4414\ : Span4Mux_v
    port map (
            O => \N__22304\,
            I => \N__22294\
        );

    \I__4413\ : InMux
    port map (
            O => \N__22303\,
            I => \N__22291\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__22300\,
            I => \c0.data_in_field_17\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__22297\,
            I => \c0.data_in_field_17\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__22294\,
            I => \c0.data_in_field_17\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__22291\,
            I => \c0.data_in_field_17\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22278\
        );

    \I__4407\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22273\
        );

    \I__4406\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22273\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22269\
        );

    \I__4404\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22266\
        );

    \I__4403\ : Span4Mux_h
    port map (
            O => \N__22269\,
            I => \N__22262\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22259\
        );

    \I__4401\ : InMux
    port map (
            O => \N__22265\,
            I => \N__22256\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__22262\,
            I => \N__22253\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__22259\,
            I => data_in_1_4
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__22256\,
            I => data_in_1_4
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__22253\,
            I => data_in_1_4
        );

    \I__4396\ : InMux
    port map (
            O => \N__22246\,
            I => \N__22242\
        );

    \I__4395\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22239\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__22242\,
            I => \N__22235\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__22239\,
            I => \N__22232\
        );

    \I__4392\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22228\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__22235\,
            I => \N__22225\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__22232\,
            I => \N__22222\
        );

    \I__4389\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22219\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__22228\,
            I => \c0.data_in_field_22\
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__22225\,
            I => \c0.data_in_field_22\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__22222\,
            I => \c0.data_in_field_22\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__22219\,
            I => \c0.data_in_field_22\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__22210\,
            I => \c0.n2005_cascade_\
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__22207\,
            I => \c0.n10_adj_1873_cascade_\
        );

    \I__4382\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22201\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__22201\,
            I => \c0.n1825\
        );

    \I__4380\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22195\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__22195\,
            I => \N__22190\
        );

    \I__4378\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22184\
        );

    \I__4377\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22184\
        );

    \I__4376\ : Span4Mux_v
    port map (
            O => \N__22190\,
            I => \N__22181\
        );

    \I__4375\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22178\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__22184\,
            I => \c0.data_in_field_55\
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__22181\,
            I => \c0.data_in_field_55\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__22178\,
            I => \c0.data_in_field_55\
        );

    \I__4371\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__22168\,
            I => \c0.n13_adj_1951\
        );

    \I__4369\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__22162\,
            I => \N__22157\
        );

    \I__4367\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22154\
        );

    \I__4366\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22151\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__22157\,
            I => \N__22146\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__22154\,
            I => \N__22146\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22142\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__22146\,
            I => \N__22138\
        );

    \I__4361\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22135\
        );

    \I__4360\ : Span4Mux_v
    port map (
            O => \N__22142\,
            I => \N__22132\
        );

    \I__4359\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22129\
        );

    \I__4358\ : Span4Mux_s2_v
    port map (
            O => \N__22138\,
            I => \N__22126\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__22135\,
            I => \c0.data_in_field_23\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__22132\,
            I => \c0.data_in_field_23\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__22129\,
            I => \c0.data_in_field_23\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__22126\,
            I => \c0.data_in_field_23\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__22117\,
            I => \N__22114\
        );

    \I__4352\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22108\
        );

    \I__4350\ : Span4Mux_v
    port map (
            O => \N__22108\,
            I => \N__22105\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__22105\,
            I => \c0.n6107\
        );

    \I__4348\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__4346\ : Span4Mux_v
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__22093\,
            I => \c0.n18_adj_1891\
        );

    \I__4344\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22086\
        );

    \I__4343\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22083\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__22086\,
            I => \c0.n1978\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__22083\,
            I => \c0.n1978\
        );

    \I__4340\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22074\
        );

    \I__4339\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22071\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__22068\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__22071\,
            I => \c0.n5261\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__22068\,
            I => \c0.n5261\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__22063\,
            I => \c0.n5689_cascade_\
        );

    \I__4334\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__4332\ : Sp12to4
    port map (
            O => \N__22054\,
            I => \N__22051\
        );

    \I__4331\ : Span12Mux_v
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__4330\ : Odrv12
    port map (
            O => \N__22048\,
            I => \c0.n5366\
        );

    \I__4329\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22042\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__22042\,
            I => \N__22039\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__22036\,
            I => \c0.n14_adj_1967\
        );

    \I__4325\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22030\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__22030\,
            I => \c0.n5276\
        );

    \I__4323\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22024\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__22024\,
            I => \N__22020\
        );

    \I__4321\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22017\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__22020\,
            I => \c0.n5201\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__22017\,
            I => \c0.n5201\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__22012\,
            I => \c0.n5276_cascade_\
        );

    \I__4317\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__22003\,
            I => \N__22000\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__22000\,
            I => \c0.n37\
        );

    \I__4313\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21994\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21989\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21986\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__21992\,
            I => \N__21983\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__21989\,
            I => \N__21980\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21977\
        );

    \I__4307\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21973\
        );

    \I__4306\ : Span4Mux_h
    port map (
            O => \N__21980\,
            I => \N__21970\
        );

    \I__4305\ : Span4Mux_h
    port map (
            O => \N__21977\,
            I => \N__21967\
        );

    \I__4304\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21964\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__21973\,
            I => \c0.data_in_field_36\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__21970\,
            I => \c0.data_in_field_36\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__21967\,
            I => \c0.data_in_field_36\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__21964\,
            I => \c0.data_in_field_36\
        );

    \I__4299\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21951\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__21954\,
            I => \N__21948\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21943\
        );

    \I__4296\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21940\
        );

    \I__4295\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21935\
        );

    \I__4294\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21935\
        );

    \I__4293\ : Span4Mux_h
    port map (
            O => \N__21943\,
            I => \N__21932\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__21940\,
            I => \c0.data_in_field_105\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__21935\,
            I => \c0.data_in_field_105\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__21932\,
            I => \c0.data_in_field_105\
        );

    \I__4289\ : CascadeMux
    port map (
            O => \N__21925\,
            I => \c0.n2095_cascade_\
        );

    \I__4288\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21915\
        );

    \I__4286\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21912\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__21915\,
            I => \N__21909\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__21912\,
            I => \N__21906\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__21909\,
            I => \c0.n1821\
        );

    \I__4282\ : Odrv12
    port map (
            O => \N__21906\,
            I => \c0.n1821\
        );

    \I__4281\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21898\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__21898\,
            I => \c0.n34_adj_1896\
        );

    \I__4279\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21891\
        );

    \I__4278\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21888\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__21891\,
            I => \N__21883\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__21888\,
            I => \N__21883\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__21883\,
            I => \N__21879\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21876\
        );

    \I__4273\ : Span4Mux_h
    port map (
            O => \N__21879\,
            I => \N__21871\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21868\
        );

    \I__4271\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21863\
        );

    \I__4270\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21863\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__21871\,
            I => \c0.data_in_field_11\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__21868\,
            I => \c0.data_in_field_11\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__21863\,
            I => \c0.data_in_field_11\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__21856\,
            I => \c0.n5821_cascade_\
        );

    \I__4265\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21850\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21847\
        );

    \I__4263\ : Span4Mux_s3_h
    port map (
            O => \N__21847\,
            I => \N__21844\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__21844\,
            I => \N__21841\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__21841\,
            I => \c0.n5423\
        );

    \I__4260\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21829\
        );

    \I__4259\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21829\
        );

    \I__4258\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21829\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__21829\,
            I => \c0.data_in_field_27\
        );

    \I__4256\ : InMux
    port map (
            O => \N__21826\,
            I => \N__21823\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__4254\ : Span4Mux_h
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__21817\,
            I => \c0.n2080\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__21814\,
            I => \c0.n2080_cascade_\
        );

    \I__4251\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21805\
        );

    \I__4250\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21805\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__21805\,
            I => \c0.n5243\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__4247\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__4245\ : Span4Mux_v
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__4244\ : Span4Mux_h
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__4243\ : Span4Mux_s2_h
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__21784\,
            I => \c0.n16_adj_1922\
        );

    \I__4241\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21778\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__21778\,
            I => \c0.n25_adj_1926\
        );

    \I__4239\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21772\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__4237\ : Span4Mux_s3_h
    port map (
            O => \N__21769\,
            I => \N__21766\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__21766\,
            I => \c0.n5429\
        );

    \I__4235\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21760\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__21760\,
            I => \N__21757\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__21757\,
            I => \N__21754\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__21754\,
            I => \c0.n5791\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21748\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__21748\,
            I => \N__21745\
        );

    \I__4229\ : Odrv12
    port map (
            O => \N__21745\,
            I => \c0.n5432\
        );

    \I__4228\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21739\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__21739\,
            I => \N__21736\
        );

    \I__4226\ : Span4Mux_h
    port map (
            O => \N__21736\,
            I => \N__21730\
        );

    \I__4225\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21727\
        );

    \I__4224\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21722\
        );

    \I__4223\ : InMux
    port map (
            O => \N__21733\,
            I => \N__21722\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__21730\,
            I => \c0.data_in_field_30\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__21727\,
            I => \c0.data_in_field_30\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__21722\,
            I => \c0.data_in_field_30\
        );

    \I__4219\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21708\
        );

    \I__4217\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21704\
        );

    \I__4216\ : Span4Mux_v
    port map (
            O => \N__21708\,
            I => \N__21701\
        );

    \I__4215\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21698\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__21704\,
            I => \N__21695\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__21701\,
            I => \N__21692\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21687\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__21695\,
            I => \N__21687\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__21692\,
            I => \c0.data_in_field_13\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__21687\,
            I => \c0.data_in_field_13\
        );

    \I__4208\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__4206\ : Span4Mux_s3_h
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__21673\,
            I => \N__21670\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__21670\,
            I => \c0.n5393\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__21667\,
            I => \N__21664\
        );

    \I__4202\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21660\
        );

    \I__4201\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21657\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__21660\,
            I => \N__21652\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__21657\,
            I => \N__21652\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__4197\ : Span4Mux_h
    port map (
            O => \N__21649\,
            I => \N__21645\
        );

    \I__4196\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21642\
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__21645\,
            I => data_in_14_7
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__21642\,
            I => data_in_14_7
        );

    \I__4193\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__21634\,
            I => \c0.n10_adj_1898\
        );

    \I__4191\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__21628\,
            I => \N__21625\
        );

    \I__4189\ : Span4Mux_s2_h
    port map (
            O => \N__21625\,
            I => \N__21621\
        );

    \I__4188\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21618\
        );

    \I__4187\ : Span4Mux_h
    port map (
            O => \N__21621\,
            I => \N__21613\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__21618\,
            I => \N__21610\
        );

    \I__4185\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21605\
        );

    \I__4184\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21605\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__21613\,
            I => \c0.data_in_field_69\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__21610\,
            I => \c0.data_in_field_69\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__21605\,
            I => \c0.data_in_field_69\
        );

    \I__4180\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__21595\,
            I => \c0.n5159\
        );

    \I__4178\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__21589\,
            I => \N__21585\
        );

    \I__4176\ : InMux
    port map (
            O => \N__21588\,
            I => \N__21582\
        );

    \I__4175\ : Span4Mux_v
    port map (
            O => \N__21585\,
            I => \N__21574\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__21582\,
            I => \N__21574\
        );

    \I__4173\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21569\
        );

    \I__4172\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21569\
        );

    \I__4171\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21566\
        );

    \I__4170\ : Span4Mux_h
    port map (
            O => \N__21574\,
            I => \N__21563\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__21569\,
            I => \c0.data_in_field_99\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__21566\,
            I => \c0.data_in_field_99\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__21563\,
            I => \c0.data_in_field_99\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__21556\,
            I => \c0.n5159_cascade_\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__21553\,
            I => \c0.n5683_cascade_\
        );

    \I__4164\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21547\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__21547\,
            I => \c0.n5695\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__21544\,
            I => \c0.n5480_cascade_\
        );

    \I__4161\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__21538\,
            I => \c0.n5483\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__21535\,
            I => \c0.n5677_cascade_\
        );

    \I__4158\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21526\
        );

    \I__4156\ : Odrv12
    port map (
            O => \N__21526\,
            I => \c0.n5680\
        );

    \I__4155\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21518\
        );

    \I__4154\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21514\
        );

    \I__4153\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21511\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21508\
        );

    \I__4151\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21505\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__21514\,
            I => data_in_18_5
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__21511\,
            I => data_in_18_5
        );

    \I__4148\ : Odrv12
    port map (
            O => \N__21508\,
            I => data_in_18_5
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__21505\,
            I => data_in_18_5
        );

    \I__4146\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__21493\,
            I => \c0.n24_adj_1895\
        );

    \I__4144\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21487\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__21487\,
            I => \N__21484\
        );

    \I__4142\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21481\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__21481\,
            I => \N__21477\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__21480\,
            I => \N__21474\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__21477\,
            I => \N__21471\
        );

    \I__4138\ : InMux
    port map (
            O => \N__21474\,
            I => \N__21468\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__21471\,
            I => rx_data_0
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__21468\,
            I => rx_data_0
        );

    \I__4135\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21459\
        );

    \I__4134\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21456\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21453\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21450\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__21453\,
            I => \N__21447\
        );

    \I__4130\ : Span12Mux_s7_v
    port map (
            O => \N__21450\,
            I => \N__21442\
        );

    \I__4129\ : Span4Mux_v
    port map (
            O => \N__21447\,
            I => \N__21439\
        );

    \I__4128\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21434\
        );

    \I__4127\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21434\
        );

    \I__4126\ : Odrv12
    port map (
            O => \N__21442\,
            I => data_in_19_0
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__21439\,
            I => data_in_19_0
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__21434\,
            I => data_in_19_0
        );

    \I__4123\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21421\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__21421\,
            I => \c0.n3567\
        );

    \I__4120\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21409\
        );

    \I__4119\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21404\
        );

    \I__4118\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21401\
        );

    \I__4117\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21398\
        );

    \I__4116\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21395\
        );

    \I__4115\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21392\
        );

    \I__4114\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21389\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__21409\,
            I => \N__21386\
        );

    \I__4112\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21381\
        );

    \I__4111\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21381\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__21404\,
            I => \N__21376\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__21401\,
            I => \N__21367\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__21398\,
            I => \N__21367\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__21395\,
            I => \N__21367\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21367\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__21389\,
            I => \N__21364\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__21386\,
            I => \N__21361\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21358\
        );

    \I__4102\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21353\
        );

    \I__4101\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21353\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__21376\,
            I => \N__21346\
        );

    \I__4099\ : Span4Mux_v
    port map (
            O => \N__21367\,
            I => \N__21346\
        );

    \I__4098\ : Span4Mux_h
    port map (
            O => \N__21364\,
            I => \N__21346\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__21361\,
            I => \N__21340\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__21358\,
            I => \N__21340\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21335\
        );

    \I__4094\ : Span4Mux_h
    port map (
            O => \N__21346\,
            I => \N__21335\
        );

    \I__4093\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21332\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__21340\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__21335\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__21332\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__21325\,
            I => \c0.n5523_cascade_\
        );

    \I__4088\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21315\
        );

    \I__4087\ : InMux
    port map (
            O => \N__21321\,
            I => \N__21309\
        );

    \I__4086\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21306\
        );

    \I__4085\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21303\
        );

    \I__4084\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21300\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__21315\,
            I => \N__21297\
        );

    \I__4082\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21294\
        );

    \I__4081\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21289\
        );

    \I__4080\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21289\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21283\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__21306\,
            I => \N__21283\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21280\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__21300\,
            I => \N__21275\
        );

    \I__4075\ : Span4Mux_v
    port map (
            O => \N__21297\,
            I => \N__21275\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21270\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__21289\,
            I => \N__21270\
        );

    \I__4072\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21267\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__21283\,
            I => \N__21262\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__21280\,
            I => \N__21262\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__21275\,
            I => \N__21258\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__21270\,
            I => \N__21255\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21250\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__21262\,
            I => \N__21250\
        );

    \I__4065\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21247\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__21258\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__21255\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__21250\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__21247\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__21238\,
            I => \N__21235\
        );

    \I__4059\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21227\
        );

    \I__4057\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21224\
        );

    \I__4056\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21221\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__21227\,
            I => \N__21218\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21215\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21212\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__21218\,
            I => \c0.n1236\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__21215\,
            I => \c0.n1236\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__21212\,
            I => \c0.n1236\
        );

    \I__4049\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21202\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__21202\,
            I => \c0.n5515\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__21199\,
            I => \c0.n5513_cascade_\
        );

    \I__4046\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21192\
        );

    \I__4045\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21183\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21180\
        );

    \I__4043\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21177\
        );

    \I__4042\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21174\
        );

    \I__4041\ : InMux
    port map (
            O => \N__21189\,
            I => \N__21169\
        );

    \I__4040\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21169\
        );

    \I__4039\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21166\
        );

    \I__4038\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21163\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21160\
        );

    \I__4036\ : Span4Mux_h
    port map (
            O => \N__21180\,
            I => \N__21149\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21149\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21149\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__21169\,
            I => \N__21149\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N__21149\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N__21143\
        );

    \I__4030\ : Span4Mux_h
    port map (
            O => \N__21160\,
            I => \N__21143\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__21149\,
            I => \N__21140\
        );

    \I__4028\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21137\
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__21143\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__21140\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__21137\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__4024\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21127\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__21127\,
            I => \tx_data_6_N_keep\
        );

    \I__4022\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21120\
        );

    \I__4021\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21116\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21113\
        );

    \I__4019\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21110\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21105\
        );

    \I__4017\ : Span4Mux_v
    port map (
            O => \N__21113\,
            I => \N__21100\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__21110\,
            I => \N__21100\
        );

    \I__4015\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21097\
        );

    \I__4014\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21094\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__21105\,
            I => \N__21091\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__21100\,
            I => \N__21088\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__21097\,
            I => data_out_10_5
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__21094\,
            I => data_out_10_5
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__21091\,
            I => data_out_10_5
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__21088\,
            I => data_out_10_5
        );

    \I__4007\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21072\
        );

    \I__4006\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21069\
        );

    \I__4005\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21066\
        );

    \I__4004\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21063\
        );

    \I__4003\ : InMux
    port map (
            O => \N__21075\,
            I => \N__21060\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__21056\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21053\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21050\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__21063\,
            I => \N__21045\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__21060\,
            I => \N__21045\
        );

    \I__3997\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21041\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__21056\,
            I => \N__21038\
        );

    \I__3995\ : Span4Mux_h
    port map (
            O => \N__21053\,
            I => \N__21035\
        );

    \I__3994\ : Span4Mux_v
    port map (
            O => \N__21050\,
            I => \N__21030\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__21045\,
            I => \N__21030\
        );

    \I__3992\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21027\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__21041\,
            I => data_out_10_1
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__21038\,
            I => data_out_10_1
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__21035\,
            I => data_out_10_1
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__21030\,
            I => data_out_10_1
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__21027\,
            I => data_out_10_1
        );

    \I__3986\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21013\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__21013\,
            I => \N__21009\
        );

    \I__3984\ : InMux
    port map (
            O => \N__21012\,
            I => \N__21003\
        );

    \I__3983\ : Span4Mux_v
    port map (
            O => \N__21009\,
            I => \N__21000\
        );

    \I__3982\ : InMux
    port map (
            O => \N__21008\,
            I => \N__20995\
        );

    \I__3981\ : InMux
    port map (
            O => \N__21007\,
            I => \N__20995\
        );

    \I__3980\ : InMux
    port map (
            O => \N__21006\,
            I => \N__20992\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__21003\,
            I => data_out_10_3
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__21000\,
            I => data_out_10_3
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__20995\,
            I => data_out_10_3
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__20992\,
            I => data_out_10_3
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__20983\,
            I => \N__20980\
        );

    \I__3974\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20976\
        );

    \I__3973\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20973\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__20976\,
            I => \N__20970\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__20973\,
            I => \N__20967\
        );

    \I__3970\ : Span4Mux_v
    port map (
            O => \N__20970\,
            I => \N__20962\
        );

    \I__3969\ : Span4Mux_s3_h
    port map (
            O => \N__20967\,
            I => \N__20962\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__20962\,
            I => \N__20959\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__20959\,
            I => n5132
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__20956\,
            I => \c0.n5839_cascade_\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__20953\,
            I => \c0.n5833_cascade_\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__20950\,
            I => \c0.n5417_cascade_\
        );

    \I__3963\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20944\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__20944\,
            I => \c0.n5414\
        );

    \I__3961\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20938\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__20938\,
            I => \c0.n5827\
        );

    \I__3959\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20927\
        );

    \I__3958\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20922\
        );

    \I__3957\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20922\
        );

    \I__3956\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20917\
        );

    \I__3955\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20917\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__20930\,
            I => \N__20912\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20908\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20903\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20903\
        );

    \I__3950\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20900\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__20915\,
            I => \N__20895\
        );

    \I__3948\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20892\
        );

    \I__3947\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20889\
        );

    \I__3946\ : Sp12to4
    port map (
            O => \N__20908\,
            I => \N__20882\
        );

    \I__3945\ : Sp12to4
    port map (
            O => \N__20903\,
            I => \N__20882\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__20900\,
            I => \N__20882\
        );

    \I__3943\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20877\
        );

    \I__3942\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20877\
        );

    \I__3941\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20874\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__20892\,
            I => \r_Rx_Data\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__20889\,
            I => \r_Rx_Data\
        );

    \I__3938\ : Odrv12
    port map (
            O => \N__20882\,
            I => \r_Rx_Data\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__20877\,
            I => \r_Rx_Data\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__20874\,
            I => \r_Rx_Data\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__20863\,
            I => \N__20860\
        );

    \I__3934\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20854\
        );

    \I__3933\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20854\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__20854\,
            I => \N__20851\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__20851\,
            I => \N__20847\
        );

    \I__3930\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20844\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__20847\,
            I => n1714
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__20844\,
            I => n1714
        );

    \I__3927\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20836\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__20836\,
            I => \N__20832\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20835\,
            I => \N__20829\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__20832\,
            I => n3342
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__20829\,
            I => n3342
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__3921\ : InMux
    port map (
            O => \N__20821\,
            I => \N__20815\
        );

    \I__3920\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20815\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__20815\,
            I => rx_data_7
        );

    \I__3918\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20808\
        );

    \I__3917\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20805\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__20808\,
            I => \N__20802\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20799\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__20802\,
            I => \N__20793\
        );

    \I__3913\ : Span4Mux_s1_v
    port map (
            O => \N__20799\,
            I => \N__20793\
        );

    \I__3912\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20790\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__20793\,
            I => data_in_17_1
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__20790\,
            I => data_in_17_1
        );

    \I__3909\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20781\
        );

    \I__3908\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20778\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20775\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__20778\,
            I => data_out_19_6
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__20775\,
            I => data_out_19_6
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__20770\,
            I => \N__20767\
        );

    \I__3903\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20764\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20760\
        );

    \I__3901\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20757\
        );

    \I__3900\ : Span4Mux_h
    port map (
            O => \N__20760\,
            I => \N__20754\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__20757\,
            I => data_out_18_6
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__20754\,
            I => data_out_18_6
        );

    \I__3897\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20745\
        );

    \I__3896\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20740\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__20745\,
            I => \N__20736\
        );

    \I__3894\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20731\
        );

    \I__3893\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20731\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__20740\,
            I => \N__20727\
        );

    \I__3891\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20724\
        );

    \I__3890\ : Span4Mux_v
    port map (
            O => \N__20736\,
            I => \N__20719\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20719\
        );

    \I__3888\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20715\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__20727\,
            I => \N__20712\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__20724\,
            I => \N__20709\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__20719\,
            I => \N__20706\
        );

    \I__3884\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20703\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__20715\,
            I => data_out_11_5
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__20712\,
            I => data_out_11_5
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__20709\,
            I => data_out_11_5
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__20706\,
            I => data_out_11_5
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__20703\,
            I => data_out_11_5
        );

    \I__3878\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20689\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__20689\,
            I => \N__20686\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__20686\,
            I => n5176
        );

    \I__3875\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20674\
        );

    \I__3873\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20671\
        );

    \I__3872\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20668\
        );

    \I__3871\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20665\
        );

    \I__3870\ : Span4Mux_v
    port map (
            O => \N__20674\,
            I => \N__20658\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__20671\,
            I => \N__20658\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20658\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__20665\,
            I => \N__20655\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__20658\,
            I => \N__20652\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__20655\,
            I => \c0.n1590\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__20652\,
            I => \c0.n1590\
        );

    \I__3863\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20635\
        );

    \I__3861\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20632\
        );

    \I__3860\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20627\
        );

    \I__3859\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20627\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__20640\,
            I => \N__20624\
        );

    \I__3857\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20621\
        );

    \I__3856\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20618\
        );

    \I__3855\ : Span4Mux_v
    port map (
            O => \N__20635\,
            I => \N__20611\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20611\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20611\
        );

    \I__3852\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20607\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__20621\,
            I => \N__20604\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__20618\,
            I => \N__20599\
        );

    \I__3849\ : Span4Mux_h
    port map (
            O => \N__20611\,
            I => \N__20599\
        );

    \I__3848\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20596\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20607\,
            I => data_out_11_6
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__20604\,
            I => data_out_11_6
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__20599\,
            I => data_out_11_6
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__20596\,
            I => data_out_11_6
        );

    \I__3843\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20576\
        );

    \I__3842\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20573\
        );

    \I__3841\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20568\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20565\
        );

    \I__3839\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20562\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20557\
        );

    \I__3837\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20557\
        );

    \I__3836\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20554\
        );

    \I__3835\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20551\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__20576\,
            I => \N__20548\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20545\
        );

    \I__3832\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20540\
        );

    \I__3831\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20540\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__20568\,
            I => \N__20531\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__20565\,
            I => \N__20531\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20531\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__20557\,
            I => \N__20531\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__20554\,
            I => \N__20525\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20525\
        );

    \I__3824\ : Span4Mux_v
    port map (
            O => \N__20548\,
            I => \N__20518\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__20545\,
            I => \N__20518\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__20540\,
            I => \N__20518\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__20531\,
            I => \N__20515\
        );

    \I__3820\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20512\
        );

    \I__3819\ : Span4Mux_v
    port map (
            O => \N__20525\,
            I => \N__20505\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__20518\,
            I => \N__20502\
        );

    \I__3817\ : Sp12to4
    port map (
            O => \N__20515\,
            I => \N__20497\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__20512\,
            I => \N__20497\
        );

    \I__3815\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20490\
        );

    \I__3814\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20490\
        );

    \I__3813\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20490\
        );

    \I__3812\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20487\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__20505\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__20502\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__3809\ : Odrv12
    port map (
            O => \N__20497\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__20490\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__20487\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__20476\,
            I => \N__20472\
        );

    \I__3805\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20463\
        );

    \I__3804\ : InMux
    port map (
            O => \N__20472\,
            I => \N__20463\
        );

    \I__3803\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20460\
        );

    \I__3802\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20456\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__20469\,
            I => \N__20453\
        );

    \I__3800\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20450\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__20463\,
            I => \N__20447\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__20460\,
            I => \N__20444\
        );

    \I__3797\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20441\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__20456\,
            I => \N__20438\
        );

    \I__3795\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20435\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20432\
        );

    \I__3793\ : Span4Mux_h
    port map (
            O => \N__20447\,
            I => \N__20427\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__20444\,
            I => \N__20427\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__20441\,
            I => data_out_10_6
        );

    \I__3790\ : Odrv12
    port map (
            O => \N__20438\,
            I => data_out_10_6
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__20435\,
            I => data_out_10_6
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__20432\,
            I => data_out_10_6
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__20427\,
            I => data_out_10_6
        );

    \I__3786\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20400\
        );

    \I__3785\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20397\
        );

    \I__3784\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20394\
        );

    \I__3783\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20388\
        );

    \I__3782\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20385\
        );

    \I__3781\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20380\
        );

    \I__3780\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20380\
        );

    \I__3779\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20373\
        );

    \I__3778\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20373\
        );

    \I__3777\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20373\
        );

    \I__3776\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20368\
        );

    \I__3775\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20368\
        );

    \I__3774\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20363\
        );

    \I__3773\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20363\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__20400\,
            I => \N__20356\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__20397\,
            I => \N__20356\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__20394\,
            I => \N__20356\
        );

    \I__3769\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20351\
        );

    \I__3768\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20348\
        );

    \I__3767\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20345\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__20388\,
            I => \N__20334\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20334\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__20380\,
            I => \N__20334\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__20373\,
            I => \N__20334\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__20368\,
            I => \N__20334\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20329\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__20356\,
            I => \N__20329\
        );

    \I__3759\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20326\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__20354\,
            I => \N__20321\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20318\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__20348\,
            I => \N__20315\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20310\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__20334\,
            I => \N__20310\
        );

    \I__3753\ : Sp12to4
    port map (
            O => \N__20329\,
            I => \N__20305\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20305\
        );

    \I__3751\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20300\
        );

    \I__3750\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20300\
        );

    \I__3749\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20297\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__20318\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__20315\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__20310\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__3745\ : Odrv12
    port map (
            O => \N__20305\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__20300\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__20297\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__3742\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20281\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20278\
        );

    \I__3740\ : Span4Mux_v
    port map (
            O => \N__20278\,
            I => \N__20275\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__20275\,
            I => \c0.n6_adj_1877\
        );

    \I__3738\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20269\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20266\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__20266\,
            I => \N__20260\
        );

    \I__3735\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20253\
        );

    \I__3734\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20253\
        );

    \I__3733\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20253\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__20260\,
            I => \c0.data_in_field_31\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__20253\,
            I => \c0.data_in_field_31\
        );

    \I__3730\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20245\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__20245\,
            I => \c0.n28_adj_1886\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__3727\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20236\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__20236\,
            I => \N__20233\
        );

    \I__3725\ : Span4Mux_h
    port map (
            O => \N__20233\,
            I => \N__20230\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__20230\,
            I => \c0.n5222\
        );

    \I__3723\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__20221\,
            I => \c0.n34\
        );

    \I__3720\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20214\
        );

    \I__3719\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20211\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20208\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20204\
        );

    \I__3716\ : Sp12to4
    port map (
            O => \N__20208\,
            I => \N__20201\
        );

    \I__3715\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20198\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__20204\,
            I => data_in_15_5
        );

    \I__3713\ : Odrv12
    port map (
            O => \N__20201\,
            I => data_in_15_5
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__20198\,
            I => data_in_15_5
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__20191\,
            I => \c0.n1686_cascade_\
        );

    \I__3710\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20182\
        );

    \I__3709\ : InMux
    port map (
            O => \N__20187\,
            I => \N__20179\
        );

    \I__3708\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20176\
        );

    \I__3707\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20173\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__20182\,
            I => \c0.data_in_field_25\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__20179\,
            I => \c0.data_in_field_25\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__20176\,
            I => \c0.data_in_field_25\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__20173\,
            I => \c0.data_in_field_25\
        );

    \I__3702\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20160\
        );

    \I__3701\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20156\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20153\
        );

    \I__3699\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20150\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20146\
        );

    \I__3697\ : Span4Mux_v
    port map (
            O => \N__20153\,
            I => \N__20143\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20140\
        );

    \I__3695\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20137\
        );

    \I__3694\ : Span4Mux_h
    port map (
            O => \N__20146\,
            I => \N__20134\
        );

    \I__3693\ : Span4Mux_h
    port map (
            O => \N__20143\,
            I => \N__20131\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__20140\,
            I => \N__20124\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20124\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__20134\,
            I => \N__20124\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__20131\,
            I => data_in_19_7
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__20124\,
            I => data_in_19_7
        );

    \I__3687\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20116\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__20116\,
            I => \N__20112\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__20115\,
            I => \N__20109\
        );

    \I__3684\ : Span4Mux_h
    port map (
            O => \N__20112\,
            I => \N__20106\
        );

    \I__3683\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20102\
        );

    \I__3682\ : Span4Mux_v
    port map (
            O => \N__20106\,
            I => \N__20099\
        );

    \I__3681\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20096\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__20102\,
            I => \c0.data_in_field_7\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__20099\,
            I => \c0.data_in_field_7\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__20096\,
            I => \c0.data_in_field_7\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__20089\,
            I => \c0.n5162_cascade_\
        );

    \I__3676\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20081\
        );

    \I__3675\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20078\
        );

    \I__3674\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20075\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20072\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20068\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20063\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__20072\,
            I => \N__20063\
        );

    \I__3669\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20060\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__20068\,
            I => data_in_18_1
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__20063\,
            I => data_in_18_1
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__20060\,
            I => data_in_18_1
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__20053\,
            I => \c0.n1825_cascade_\
        );

    \I__3664\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20047\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__20044\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__20044\,
            I => \N__20037\
        );

    \I__3661\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20034\
        );

    \I__3660\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20031\
        );

    \I__3659\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20026\
        );

    \I__3658\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20026\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__20037\,
            I => \c0.data_in_field_133\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__20034\,
            I => \c0.data_in_field_133\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__20031\,
            I => \c0.data_in_field_133\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__20026\,
            I => \c0.data_in_field_133\
        );

    \I__3653\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20009\
        );

    \I__3651\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20006\
        );

    \I__3650\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20002\
        );

    \I__3649\ : Span4Mux_h
    port map (
            O => \N__20009\,
            I => \N__19999\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__20006\,
            I => \N__19996\
        );

    \I__3647\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19993\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__20002\,
            I => \c0.data_in_field_73\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__19999\,
            I => \c0.data_in_field_73\
        );

    \I__3644\ : Odrv12
    port map (
            O => \N__19996\,
            I => \c0.data_in_field_73\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__19993\,
            I => \c0.data_in_field_73\
        );

    \I__3642\ : InMux
    port map (
            O => \N__19984\,
            I => \N__19980\
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__19983\,
            I => \N__19976\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__19980\,
            I => \N__19973\
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__19979\,
            I => \N__19970\
        );

    \I__3638\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19966\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__19973\,
            I => \N__19963\
        );

    \I__3636\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19958\
        );

    \I__3635\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19958\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__19966\,
            I => \c0.data_in_field_35\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__19963\,
            I => \c0.data_in_field_35\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__19958\,
            I => \c0.data_in_field_35\
        );

    \I__3631\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__3629\ : Span4Mux_v
    port map (
            O => \N__19945\,
            I => \N__19942\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__19942\,
            I => \c0.n18\
        );

    \I__3627\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19936\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19932\
        );

    \I__3625\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19929\
        );

    \I__3624\ : Span4Mux_s2_h
    port map (
            O => \N__19932\,
            I => \N__19924\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19924\
        );

    \I__3622\ : Span4Mux_h
    port map (
            O => \N__19924\,
            I => \N__19919\
        );

    \I__3621\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19914\
        );

    \I__3620\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19914\
        );

    \I__3619\ : Odrv4
    port map (
            O => \N__19919\,
            I => \c0.data_in_field_137\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__19914\,
            I => \c0.data_in_field_137\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__19909\,
            I => \N__19906\
        );

    \I__3616\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19900\
        );

    \I__3615\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19900\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19897\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__19894\,
            I => \c0.n2036\
        );

    \I__3611\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__19888\,
            I => \c0.n20_adj_1892\
        );

    \I__3609\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19881\
        );

    \I__3608\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19878\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__19881\,
            I => \c0.n2033\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__19878\,
            I => \c0.n2033\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__19873\,
            I => \c0.n10_adj_1963_cascade_\
        );

    \I__3604\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__19867\,
            I => \c0.n5114\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__19864\,
            I => \c0.n5114_cascade_\
        );

    \I__3601\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19858\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19855\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__19855\,
            I => \c0.n30_adj_1903\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__19852\,
            I => \N__19849\
        );

    \I__3597\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19846\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__19846\,
            I => \N__19843\
        );

    \I__3595\ : Span4Mux_h
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__19840\,
            I => \N__19837\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__19837\,
            I => \c0.n5743\
        );

    \I__3592\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19831\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__19831\,
            I => \N__19827\
        );

    \I__3590\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19821\
        );

    \I__3589\ : Span4Mux_s3_v
    port map (
            O => \N__19827\,
            I => \N__19818\
        );

    \I__3588\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19811\
        );

    \I__3587\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19811\
        );

    \I__3586\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19811\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__19821\,
            I => \c0.data_in_field_87\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__19818\,
            I => \c0.data_in_field_87\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__19811\,
            I => \c0.data_in_field_87\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__19804\,
            I => \N__19801\
        );

    \I__3581\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19797\
        );

    \I__3580\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19794\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__19797\,
            I => \N__19788\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19785\
        );

    \I__3577\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19782\
        );

    \I__3576\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19777\
        );

    \I__3575\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19777\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__19788\,
            I => \N__19772\
        );

    \I__3573\ : Span4Mux_s3_v
    port map (
            O => \N__19785\,
            I => \N__19772\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__19782\,
            I => \N__19769\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__19777\,
            I => \c0.data_in_field_57\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__19772\,
            I => \c0.data_in_field_57\
        );

    \I__3569\ : Odrv12
    port map (
            O => \N__19769\,
            I => \c0.data_in_field_57\
        );

    \I__3568\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__19759\,
            I => \c0.n5198\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__19756\,
            I => \N__19753\
        );

    \I__3565\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19750\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19747\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__19747\,
            I => \N__19743\
        );

    \I__3562\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19740\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__19743\,
            I => \N__19737\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__19740\,
            I => \c0.n1918\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__19737\,
            I => \c0.n1918\
        );

    \I__3558\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__19729\,
            I => \c0.n18_adj_1910\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__19726\,
            I => \c0.n17_adj_1912_cascade_\
        );

    \I__3555\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19720\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__19720\,
            I => \c0.n12_adj_1911\
        );

    \I__3553\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19714\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__19714\,
            I => \c0.n19_adj_1920\
        );

    \I__3551\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__19708\,
            I => \c0.n28_adj_1902\
        );

    \I__3549\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19702\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__19702\,
            I => \c0.n32\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__19699\,
            I => \c0.n29_adj_1905_cascade_\
        );

    \I__3546\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__19693\,
            I => \c0.n31_adj_1904\
        );

    \I__3544\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__19684\,
            I => \c0.n5278\
        );

    \I__3541\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19677\
        );

    \I__3540\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19674\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__19677\,
            I => \N__19671\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__19674\,
            I => \N__19663\
        );

    \I__3537\ : Span4Mux_h
    port map (
            O => \N__19671\,
            I => \N__19663\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19660\
        );

    \I__3535\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19657\
        );

    \I__3534\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19654\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__19663\,
            I => \c0.data_in_field_134\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__19660\,
            I => \c0.data_in_field_134\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__19657\,
            I => \c0.data_in_field_134\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__19654\,
            I => \c0.data_in_field_134\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__19645\,
            I => \c0.n12_cascade_\
        );

    \I__3528\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19638\
        );

    \I__3527\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19635\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__19638\,
            I => \c0.n1880\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__19635\,
            I => \c0.n1880\
        );

    \I__3524\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19626\
        );

    \I__3523\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19623\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__19626\,
            I => \N__19620\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19615\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__19620\,
            I => \N__19615\
        );

    \I__3519\ : Sp12to4
    port map (
            O => \N__19615\,
            I => \N__19611\
        );

    \I__3518\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19608\
        );

    \I__3517\ : Odrv12
    port map (
            O => \N__19611\,
            I => data_in_15_0
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__19608\,
            I => data_in_15_0
        );

    \I__3515\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19597\
        );

    \I__3514\ : InMux
    port map (
            O => \N__19602\,
            I => \N__19597\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19594\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__19594\,
            I => \c0.n5210\
        );

    \I__3511\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19588\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__19588\,
            I => \c0.tx2_transmit_N_1031\
        );

    \I__3509\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19581\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__19584\,
            I => \N__19578\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__19581\,
            I => \N__19575\
        );

    \I__3506\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19572\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__19575\,
            I => \c0.n1785\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__19572\,
            I => \c0.n1785\
        );

    \I__3503\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19564\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__19564\,
            I => \c0.n11\
        );

    \I__3501\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19558\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19555\
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__19555\,
            I => \c0.n24_adj_1924\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__19552\,
            I => \c0.n5259_cascade_\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__19549\,
            I => \N__19546\
        );

    \I__3496\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19543\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__19543\,
            I => \c0.n21_adj_1933\
        );

    \I__3494\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19537\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__19537\,
            I => \N__19534\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__19534\,
            I => \c0.n16\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__19531\,
            I => \N__19528\
        );

    \I__3490\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__19525\,
            I => \N__19522\
        );

    \I__3488\ : Span4Mux_h
    port map (
            O => \N__19522\,
            I => \N__19519\
        );

    \I__3487\ : Span4Mux_s3_h
    port map (
            O => \N__19519\,
            I => \N__19515\
        );

    \I__3486\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19512\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__19515\,
            I => \c0.n1893\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__19512\,
            I => \c0.n1893\
        );

    \I__3483\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19504\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__19504\,
            I => \N__19500\
        );

    \I__3481\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19497\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__19500\,
            I => \N__19494\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19491\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__19494\,
            I => \c0.n2008\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__19491\,
            I => \c0.n2008\
        );

    \I__3476\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__19480\,
            I => \c0.n5225\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__19477\,
            I => \c0.n5198_cascade_\
        );

    \I__3472\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__19471\,
            I => \N__19467\
        );

    \I__3470\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19464\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__19467\,
            I => \N__19461\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__19464\,
            I => \N__19458\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__19461\,
            I => \c0.n6103\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__19458\,
            I => \c0.n6103\
        );

    \I__3465\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19450\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__19450\,
            I => \c0.n28\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__19447\,
            I => \N__19444\
        );

    \I__3462\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19441\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__19441\,
            I => \N__19437\
        );

    \I__3460\ : InMux
    port map (
            O => \N__19440\,
            I => \N__19434\
        );

    \I__3459\ : Span4Mux_v
    port map (
            O => \N__19437\,
            I => \N__19430\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19427\
        );

    \I__3457\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19424\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__19430\,
            I => data_in_14_5
        );

    \I__3455\ : Odrv12
    port map (
            O => \N__19427\,
            I => data_in_14_5
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__19424\,
            I => data_in_14_5
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__19417\,
            I => \N__19414\
        );

    \I__3452\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__19411\,
            I => \N__19408\
        );

    \I__3450\ : Span4Mux_h
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__19405\,
            I => \c0.n5809\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__3447\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19396\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__19393\,
            I => \c0.n5241\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__19390\,
            I => \c0.tx2_transmit_N_1031_cascade_\
        );

    \I__3443\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19384\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__19384\,
            I => \N__19381\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__19381\,
            I => \c0.n38_adj_1934\
        );

    \I__3440\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__19375\,
            I => \c0.n14_adj_1900\
        );

    \I__3438\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19363\
        );

    \I__3437\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19363\
        );

    \I__3436\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19360\
        );

    \I__3435\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19357\
        );

    \I__3434\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19354\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__19363\,
            I => \N__19351\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__19360\,
            I => \N__19346\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__19357\,
            I => \N__19346\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__19354\,
            I => \N__19343\
        );

    \I__3429\ : Span4Mux_v
    port map (
            O => \N__19351\,
            I => \N__19337\
        );

    \I__3428\ : Span4Mux_v
    port map (
            O => \N__19346\,
            I => \N__19332\
        );

    \I__3427\ : Span4Mux_v
    port map (
            O => \N__19343\,
            I => \N__19332\
        );

    \I__3426\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19329\
        );

    \I__3425\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19326\
        );

    \I__3424\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19323\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__19337\,
            I => n1442
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__19332\,
            I => n1442
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__19329\,
            I => n1442
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__19326\,
            I => n1442
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__19323\,
            I => n1442
        );

    \I__3418\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19308\
        );

    \I__3417\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19305\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__19308\,
            I => \r_Tx_Data_6\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__19305\,
            I => \r_Tx_Data_6\
        );

    \I__3414\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19293\
        );

    \I__3413\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19287\
        );

    \I__3412\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19287\
        );

    \I__3411\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19284\
        );

    \I__3410\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19279\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__19293\,
            I => \N__19276\
        );

    \I__3408\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19273\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__19287\,
            I => \N__19268\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__19284\,
            I => \N__19268\
        );

    \I__3405\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19265\
        );

    \I__3404\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19262\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__19279\,
            I => \N__19257\
        );

    \I__3402\ : Span4Mux_v
    port map (
            O => \N__19276\,
            I => \N__19257\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__19273\,
            I => \N__19252\
        );

    \I__3400\ : Span4Mux_h
    port map (
            O => \N__19268\,
            I => \N__19252\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19249\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__19262\,
            I => data_out_10_0
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__19257\,
            I => data_out_10_0
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__19252\,
            I => data_out_10_0
        );

    \I__3395\ : Odrv12
    port map (
            O => \N__19249\,
            I => data_out_10_0
        );

    \I__3394\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19237\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__19237\,
            I => \N__19234\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__19234\,
            I => \N__19231\
        );

    \I__3391\ : Span4Mux_s3_h
    port map (
            O => \N__19231\,
            I => \N__19228\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__19228\,
            I => n1748
        );

    \I__3389\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19217\
        );

    \I__3388\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19214\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19210\
        );

    \I__3386\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19202\
        );

    \I__3385\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19202\
        );

    \I__3384\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19199\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19196\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__19214\,
            I => \N__19193\
        );

    \I__3381\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19188\
        );

    \I__3380\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19188\
        );

    \I__3379\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19185\
        );

    \I__3378\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19182\
        );

    \I__3377\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19171\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19168\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__19199\,
            I => \N__19160\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__19196\,
            I => \N__19160\
        );

    \I__3373\ : Span4Mux_h
    port map (
            O => \N__19193\,
            I => \N__19160\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__19188\,
            I => \N__19153\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19153\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__19182\,
            I => \N__19153\
        );

    \I__3369\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19142\
        );

    \I__3368\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19142\
        );

    \I__3367\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19142\
        );

    \I__3366\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19142\
        );

    \I__3365\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19142\
        );

    \I__3364\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19135\
        );

    \I__3363\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19135\
        );

    \I__3362\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19135\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__19171\,
            I => \N__19132\
        );

    \I__3360\ : Span4Mux_h
    port map (
            O => \N__19168\,
            I => \N__19129\
        );

    \I__3359\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19126\
        );

    \I__3358\ : Span4Mux_v
    port map (
            O => \N__19160\,
            I => \N__19123\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__19153\,
            I => \N__19118\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19118\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__19135\,
            I => n21_adj_1999
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__19132\,
            I => n21_adj_1999
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__19129\,
            I => n21_adj_1999
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__19126\,
            I => n21_adj_1999
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__19123\,
            I => n21_adj_1999
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__19118\,
            I => n21_adj_1999
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__3348\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19099\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__19095\
        );

    \I__3346\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19092\
        );

    \I__3345\ : Odrv12
    port map (
            O => \N__19095\,
            I => data_10
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__19092\,
            I => data_10
        );

    \I__3343\ : InMux
    port map (
            O => \N__19087\,
            I => \N__19084\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__19084\,
            I => \N__19075\
        );

    \I__3341\ : InMux
    port map (
            O => \N__19083\,
            I => \N__19072\
        );

    \I__3340\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19065\
        );

    \I__3339\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19065\
        );

    \I__3338\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19065\
        );

    \I__3337\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19062\
        );

    \I__3336\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19059\
        );

    \I__3335\ : Span4Mux_h
    port map (
            O => \N__19075\,
            I => \N__19051\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__19072\,
            I => \N__19051\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__19065\,
            I => \N__19046\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__19062\,
            I => \N__19046\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__19059\,
            I => \N__19043\
        );

    \I__3330\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19040\
        );

    \I__3329\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19035\
        );

    \I__3328\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19035\
        );

    \I__3327\ : Span4Mux_v
    port map (
            O => \N__19051\,
            I => \N__19024\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__19046\,
            I => \N__19021\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__19043\,
            I => \N__19016\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19016\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__19013\
        );

    \I__3322\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19008\
        );

    \I__3321\ : InMux
    port map (
            O => \N__19033\,
            I => \N__19008\
        );

    \I__3320\ : InMux
    port map (
            O => \N__19032\,
            I => \N__18997\
        );

    \I__3319\ : InMux
    port map (
            O => \N__19031\,
            I => \N__18997\
        );

    \I__3318\ : InMux
    port map (
            O => \N__19030\,
            I => \N__18997\
        );

    \I__3317\ : InMux
    port map (
            O => \N__19029\,
            I => \N__18997\
        );

    \I__3316\ : InMux
    port map (
            O => \N__19028\,
            I => \N__18997\
        );

    \I__3315\ : InMux
    port map (
            O => \N__19027\,
            I => \N__18994\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__19024\,
            I => n4315
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__19021\,
            I => n4315
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__19016\,
            I => n4315
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__19013\,
            I => n4315
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__19008\,
            I => n4315
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__18997\,
            I => n4315
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__18994\,
            I => n4315
        );

    \I__3307\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18973\
        );

    \I__3306\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18968\
        );

    \I__3305\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18968\
        );

    \I__3304\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18964\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__18973\,
            I => \N__18959\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__18968\,
            I => \N__18959\
        );

    \I__3301\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18956\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18951\
        );

    \I__3299\ : Span4Mux_v
    port map (
            O => \N__18959\,
            I => \N__18946\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__18956\,
            I => \N__18946\
        );

    \I__3297\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18943\
        );

    \I__3296\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18940\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__18951\,
            I => \N__18935\
        );

    \I__3294\ : Span4Mux_h
    port map (
            O => \N__18946\,
            I => \N__18935\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__18943\,
            I => data_out_10_2
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__18940\,
            I => data_out_10_2
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__18935\,
            I => data_out_10_2
        );

    \I__3290\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18925\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__18925\,
            I => \N__18922\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__18922\,
            I => \N__18919\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__18919\,
            I => \c0.n5411\
        );

    \I__3286\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18913\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__18913\,
            I => \N__18910\
        );

    \I__3284\ : Span4Mux_h
    port map (
            O => \N__18910\,
            I => \N__18907\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__18907\,
            I => \c0.n5830\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__18904\,
            I => \N__18901\
        );

    \I__3281\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18898\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18895\
        );

    \I__3279\ : Span4Mux_h
    port map (
            O => \N__18895\,
            I => \N__18892\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__18892\,
            I => \c0.n5941\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__18889\,
            I => \N__18885\
        );

    \I__3276\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18882\
        );

    \I__3275\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18879\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__18882\,
            I => \c0.data_in_frame_19_2\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__18879\,
            I => \c0.data_in_frame_19_2\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__18874\,
            I => \N__18871\
        );

    \I__3271\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18865\
        );

    \I__3270\ : InMux
    port map (
            O => \N__18870\,
            I => \N__18865\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__18865\,
            I => \c0.data_in_frame_18_5\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__18862\,
            I => \N__18858\
        );

    \I__3267\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18853\
        );

    \I__3266\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18853\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__18853\,
            I => \c0.data_in_frame_19_5\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__18850\,
            I => \N__18847\
        );

    \I__3263\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18840\
        );

    \I__3261\ : InMux
    port map (
            O => \N__18843\,
            I => \N__18837\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__18840\,
            I => data_4
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__18837\,
            I => data_4
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__18832\,
            I => \N__18829\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18825\
        );

    \I__3256\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18822\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__18825\,
            I => data_14
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18822\,
            I => data_14
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__18817\,
            I => \N__18814\
        );

    \I__3252\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18810\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__18813\,
            I => \N__18807\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__18810\,
            I => \N__18802\
        );

    \I__3249\ : InMux
    port map (
            O => \N__18807\,
            I => \N__18799\
        );

    \I__3248\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18796\
        );

    \I__3247\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18793\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__18802\,
            I => \N__18785\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__18799\,
            I => \N__18785\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__18796\,
            I => \N__18785\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__18793\,
            I => \N__18782\
        );

    \I__3242\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18776\
        );

    \I__3241\ : Span4Mux_v
    port map (
            O => \N__18785\,
            I => \N__18771\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__18782\,
            I => \N__18771\
        );

    \I__3239\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18768\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18763\
        );

    \I__3237\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18763\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__18776\,
            I => data_out_11_4
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__18771\,
            I => data_out_11_4
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__18768\,
            I => data_out_11_4
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__18763\,
            I => data_out_11_4
        );

    \I__3232\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18751\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__18751\,
            I => \N__18745\
        );

    \I__3230\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18742\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__18749\,
            I => \N__18739\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18736\
        );

    \I__3227\ : Span4Mux_s3_h
    port map (
            O => \N__18745\,
            I => \N__18730\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__18742\,
            I => \N__18730\
        );

    \I__3225\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18727\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__18736\,
            I => \N__18724\
        );

    \I__3223\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18721\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__18730\,
            I => \N__18718\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__18727\,
            I => data_out_10_4
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__18724\,
            I => data_out_10_4
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__18721\,
            I => data_out_10_4
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__18718\,
            I => data_out_10_4
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__18709\,
            I => \c0.n9_adj_1887_cascade_\
        );

    \I__3216\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__18703\,
            I => \N__18700\
        );

    \I__3214\ : Odrv12
    port map (
            O => \N__18700\,
            I => \c0.n15_adj_1889\
        );

    \I__3213\ : InMux
    port map (
            O => \N__18697\,
            I => \N__18693\
        );

    \I__3212\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18690\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__18693\,
            I => data_8
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__18690\,
            I => data_8
        );

    \I__3209\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__18679\,
            I => \N__18676\
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__18676\,
            I => \c0.n17_adj_1961\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__18673\,
            I => \c0.n1236_cascade_\
        );

    \I__3204\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18667\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__18667\,
            I => \c0.n2247\
        );

    \I__3202\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18661\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18661\,
            I => \N__18658\
        );

    \I__3200\ : Span4Mux_v
    port map (
            O => \N__18658\,
            I => \N__18654\
        );

    \I__3199\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18651\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__18654\,
            I => \c0.n1227\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__18651\,
            I => \c0.n1227\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__18646\,
            I => \c0.n5511_cascade_\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__18643\,
            I => \tx_data_7_N_keep_cascade_\
        );

    \I__3194\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18636\
        );

    \I__3193\ : InMux
    port map (
            O => \N__18639\,
            I => \N__18633\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__18636\,
            I => \r_Tx_Data_7\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__18633\,
            I => \r_Tx_Data_7\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__18628\,
            I => \N__18625\
        );

    \I__3189\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18622\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__18622\,
            I => \N__18619\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__18619\,
            I => \N__18615\
        );

    \I__3186\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18612\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__18615\,
            I => data_7
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__18612\,
            I => data_7
        );

    \I__3183\ : InMux
    port map (
            O => \N__18607\,
            I => \c0.n4391\
        );

    \I__3182\ : InMux
    port map (
            O => \N__18604\,
            I => \bfn_6_18_0_\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__3180\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18595\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__18595\,
            I => \N__18592\
        );

    \I__3178\ : Span4Mux_v
    port map (
            O => \N__18592\,
            I => \N__18588\
        );

    \I__3177\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18585\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__18588\,
            I => data_9
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__18585\,
            I => data_9
        );

    \I__3174\ : InMux
    port map (
            O => \N__18580\,
            I => \c0.n4393\
        );

    \I__3173\ : InMux
    port map (
            O => \N__18577\,
            I => \c0.n4394\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__18574\,
            I => \N__18571\
        );

    \I__3171\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18568\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__18568\,
            I => \N__18564\
        );

    \I__3169\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18561\
        );

    \I__3168\ : Odrv12
    port map (
            O => \N__18564\,
            I => data_11
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__18561\,
            I => data_11
        );

    \I__3166\ : InMux
    port map (
            O => \N__18556\,
            I => \c0.n4395\
        );

    \I__3165\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18550\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18546\
        );

    \I__3163\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18543\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__18546\,
            I => data_12
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__18543\,
            I => data_12
        );

    \I__3160\ : InMux
    port map (
            O => \N__18538\,
            I => \c0.n4396\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__18535\,
            I => \N__18532\
        );

    \I__3158\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18529\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__18529\,
            I => \N__18525\
        );

    \I__3156\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18522\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__18525\,
            I => data_13
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__18522\,
            I => data_13
        );

    \I__3153\ : InMux
    port map (
            O => \N__18517\,
            I => \c0.n4397\
        );

    \I__3152\ : InMux
    port map (
            O => \N__18514\,
            I => \c0.n4398\
        );

    \I__3151\ : InMux
    port map (
            O => \N__18511\,
            I => \c0.n4399\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__18508\,
            I => \N__18505\
        );

    \I__3149\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18501\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18498\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__18501\,
            I => \N__18495\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__18498\,
            I => data_15
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__18495\,
            I => data_15
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__18490\,
            I => \N__18487\
        );

    \I__3143\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18483\
        );

    \I__3142\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18480\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__18483\,
            I => data_0
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__18480\,
            I => data_0
        );

    \I__3139\ : InMux
    port map (
            O => \N__18475\,
            I => \bfn_6_17_0_\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__3137\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__3135\ : Span4Mux_h
    port map (
            O => \N__18463\,
            I => \N__18459\
        );

    \I__3134\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18456\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__18459\,
            I => data_1
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__18456\,
            I => data_1
        );

    \I__3131\ : InMux
    port map (
            O => \N__18451\,
            I => \c0.n4385\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__18448\,
            I => \N__18445\
        );

    \I__3129\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18442\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__18442\,
            I => \N__18438\
        );

    \I__3127\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18435\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__18438\,
            I => data_2
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__18435\,
            I => data_2
        );

    \I__3124\ : InMux
    port map (
            O => \N__18430\,
            I => \c0.n4386\
        );

    \I__3123\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18424\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18420\
        );

    \I__3121\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18417\
        );

    \I__3120\ : Odrv12
    port map (
            O => \N__18420\,
            I => data_3
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__18417\,
            I => data_3
        );

    \I__3118\ : InMux
    port map (
            O => \N__18412\,
            I => \c0.n4387\
        );

    \I__3117\ : InMux
    port map (
            O => \N__18409\,
            I => \c0.n4388\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__18406\,
            I => \N__18403\
        );

    \I__3115\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18400\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__18400\,
            I => \N__18397\
        );

    \I__3113\ : Span4Mux_s3_h
    port map (
            O => \N__18397\,
            I => \N__18393\
        );

    \I__3112\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18390\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__18393\,
            I => data_5
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__18390\,
            I => data_5
        );

    \I__3109\ : InMux
    port map (
            O => \N__18385\,
            I => \c0.n4389\
        );

    \I__3108\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18379\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__18379\,
            I => \N__18375\
        );

    \I__3106\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18372\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__18375\,
            I => data_6
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__18372\,
            I => data_6
        );

    \I__3103\ : InMux
    port map (
            O => \N__18367\,
            I => \c0.n4390\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__18364\,
            I => \N__18358\
        );

    \I__3101\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18349\
        );

    \I__3100\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18349\
        );

    \I__3099\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18344\
        );

    \I__3098\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18344\
        );

    \I__3097\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18341\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__18356\,
            I => \N__18338\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__18355\,
            I => \N__18334\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__18354\,
            I => \N__18331\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__18349\,
            I => \N__18325\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__18344\,
            I => \N__18322\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__18341\,
            I => \N__18319\
        );

    \I__3090\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18314\
        );

    \I__3089\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18314\
        );

    \I__3088\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18309\
        );

    \I__3087\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18309\
        );

    \I__3086\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18306\
        );

    \I__3085\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18301\
        );

    \I__3084\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18301\
        );

    \I__3083\ : Span4Mux_s1_h
    port map (
            O => \N__18325\,
            I => \N__18292\
        );

    \I__3082\ : Span4Mux_h
    port map (
            O => \N__18322\,
            I => \N__18292\
        );

    \I__3081\ : Span4Mux_h
    port map (
            O => \N__18319\,
            I => \N__18292\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__18314\,
            I => \N__18292\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__18309\,
            I => \r_SM_Main_2_adj_2005\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__18306\,
            I => \r_SM_Main_2_adj_2005\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__18301\,
            I => \r_SM_Main_2_adj_2005\
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__18292\,
            I => \r_SM_Main_2_adj_2005\
        );

    \I__3075\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18273\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__18282\,
            I => \N__18270\
        );

    \I__3073\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18261\
        );

    \I__3072\ : InMux
    port map (
            O => \N__18280\,
            I => \N__18261\
        );

    \I__3071\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18258\
        );

    \I__3070\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18255\
        );

    \I__3069\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18252\
        );

    \I__3068\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18249\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__18273\,
            I => \N__18243\
        );

    \I__3066\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18238\
        );

    \I__3065\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18238\
        );

    \I__3064\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18233\
        );

    \I__3063\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18233\
        );

    \I__3062\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18230\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__18261\,
            I => \N__18227\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__18258\,
            I => \N__18220\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__18255\,
            I => \N__18220\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__18252\,
            I => \N__18220\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__18249\,
            I => \N__18217\
        );

    \I__3056\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18210\
        );

    \I__3055\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18210\
        );

    \I__3054\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18210\
        );

    \I__3053\ : Span4Mux_v
    port map (
            O => \N__18243\,
            I => \N__18205\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__18238\,
            I => \N__18205\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__18233\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__18230\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__18227\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3048\ : Odrv12
    port map (
            O => \N__18220\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__18217\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__18210\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__18205\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__3044\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18187\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__18187\,
            I => \c0.rx.n5058\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__18184\,
            I => \N__18181\
        );

    \I__3041\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18171\
        );

    \I__3040\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18171\
        );

    \I__3039\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18168\
        );

    \I__3038\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18165\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__18177\,
            I => \N__18162\
        );

    \I__3036\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18159\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__18171\,
            I => \N__18152\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__18168\,
            I => \N__18152\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__18165\,
            I => \N__18152\
        );

    \I__3032\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18149\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__18159\,
            I => \N__18144\
        );

    \I__3030\ : Span4Mux_h
    port map (
            O => \N__18152\,
            I => \N__18144\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__18149\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__18144\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__3026\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18125\
        );

    \I__3025\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18125\
        );

    \I__3024\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18120\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18120\
        );

    \I__3022\ : InMux
    port map (
            O => \N__18132\,
            I => \N__18117\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__18131\,
            I => \N__18113\
        );

    \I__3020\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18106\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__18125\,
            I => \N__18103\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__18120\,
            I => \N__18098\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__18117\,
            I => \N__18098\
        );

    \I__3016\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18091\
        );

    \I__3015\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18091\
        );

    \I__3014\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18091\
        );

    \I__3013\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18086\
        );

    \I__3012\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18086\
        );

    \I__3011\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18083\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__18106\,
            I => \r_SM_Main_0_adj_2006\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__18103\,
            I => \r_SM_Main_0_adj_2006\
        );

    \I__3008\ : Odrv12
    port map (
            O => \N__18098\,
            I => \r_SM_Main_0_adj_2006\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__18091\,
            I => \r_SM_Main_0_adj_2006\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__18086\,
            I => \r_SM_Main_0_adj_2006\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__18083\,
            I => \r_SM_Main_0_adj_2006\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__18070\,
            I => \c0.rx.n5058_cascade_\
        );

    \I__3003\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18062\
        );

    \I__3002\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18057\
        );

    \I__3001\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18057\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__18062\,
            I => \N__18050\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__18057\,
            I => \N__18050\
        );

    \I__2998\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18041\
        );

    \I__2997\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18041\
        );

    \I__2996\ : Span4Mux_s1_v
    port map (
            O => \N__18050\,
            I => \N__18038\
        );

    \I__2995\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18035\
        );

    \I__2994\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18030\
        );

    \I__2993\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18030\
        );

    \I__2992\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18027\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__18041\,
            I => \c0.rx.r_SM_Main_2_N_1824_2\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__18038\,
            I => \c0.rx.r_SM_Main_2_N_1824_2\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__18035\,
            I => \c0.rx.r_SM_Main_2_N_1824_2\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__18030\,
            I => \c0.rx.r_SM_Main_2_N_1824_2\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__18027\,
            I => \c0.rx.r_SM_Main_2_N_1824_2\
        );

    \I__2986\ : InMux
    port map (
            O => \N__18016\,
            I => \N__18012\
        );

    \I__2985\ : InMux
    port map (
            O => \N__18015\,
            I => \N__18009\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__18012\,
            I => \N__18004\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__18009\,
            I => \N__18004\
        );

    \I__2982\ : Odrv12
    port map (
            O => \N__18004\,
            I => n4
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__18001\,
            I => \n1714_cascade_\
        );

    \I__2980\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17995\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__17995\,
            I => \N__17991\
        );

    \I__2978\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17988\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__17991\,
            I => rx_data_1
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__17988\,
            I => rx_data_1
        );

    \I__2975\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17978\
        );

    \I__2974\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17973\
        );

    \I__2973\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17973\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__17978\,
            I => data_in_0_7
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__17973\,
            I => data_in_0_7
        );

    \I__2970\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17961\
        );

    \I__2968\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17958\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__17961\,
            I => n4_adj_1986
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__17958\,
            I => n4_adj_1986
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__17953\,
            I => \N__17949\
        );

    \I__2964\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17945\
        );

    \I__2963\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17940\
        );

    \I__2962\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17940\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__17945\,
            I => n1709
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__17940\,
            I => n1709
        );

    \I__2959\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17931\
        );

    \I__2958\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17928\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__17931\,
            I => \N__17925\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__17928\,
            I => \N__17922\
        );

    \I__2955\ : Span4Mux_v
    port map (
            O => \N__17925\,
            I => \N__17918\
        );

    \I__2954\ : Span4Mux_s3_h
    port map (
            O => \N__17922\,
            I => \N__17915\
        );

    \I__2953\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17912\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__17918\,
            I => data_in_16_6
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__17915\,
            I => data_in_16_6
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__17912\,
            I => data_in_16_6
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__17905\,
            I => \N__17902\
        );

    \I__2948\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17899\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__17899\,
            I => \c0.n5731\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__17896\,
            I => \N__17893\
        );

    \I__2945\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17890\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__17890\,
            I => \N__17887\
        );

    \I__2943\ : Span4Mux_h
    port map (
            O => \N__17887\,
            I => \N__17884\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__17884\,
            I => \c0.n5264\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__17881\,
            I => \c0.n5264_cascade_\
        );

    \I__2940\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17874\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__17877\,
            I => \N__17871\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__17874\,
            I => \N__17868\
        );

    \I__2937\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17863\
        );

    \I__2936\ : Span4Mux_h
    port map (
            O => \N__17868\,
            I => \N__17860\
        );

    \I__2935\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17855\
        );

    \I__2934\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17855\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__17863\,
            I => \N__17852\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__17860\,
            I => data_in_19_1
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__17855\,
            I => data_in_19_1
        );

    \I__2930\ : Odrv12
    port map (
            O => \N__17852\,
            I => data_in_19_1
        );

    \I__2929\ : InMux
    port map (
            O => \N__17845\,
            I => \N__17841\
        );

    \I__2928\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17838\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17833\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17830\
        );

    \I__2925\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17827\
        );

    \I__2924\ : InMux
    port map (
            O => \N__17836\,
            I => \N__17824\
        );

    \I__2923\ : Odrv12
    port map (
            O => \N__17833\,
            I => data_in_2_3
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__17830\,
            I => data_in_2_3
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__17827\,
            I => data_in_2_3
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__17824\,
            I => data_in_2_3
        );

    \I__2919\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17812\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__17812\,
            I => \c0.n39\
        );

    \I__2917\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17806\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__17806\,
            I => \c0.n45_adj_1885\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__17803\,
            I => \N__17800\
        );

    \I__2914\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17797\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__17797\,
            I => \N__17794\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__17794\,
            I => \c0.n43\
        );

    \I__2911\ : InMux
    port map (
            O => \N__17791\,
            I => \N__17788\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__17788\,
            I => \N__17785\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__17785\,
            I => \N__17782\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__17782\,
            I => \c0.n30\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__17779\,
            I => \c0.n5275_cascade_\
        );

    \I__2906\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17773\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__17773\,
            I => \N__17770\
        );

    \I__2904\ : Span4Mux_h
    port map (
            O => \N__17770\,
            I => \N__17767\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__17767\,
            I => \c0.n24_adj_1929\
        );

    \I__2902\ : InMux
    port map (
            O => \N__17764\,
            I => \N__17761\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__17761\,
            I => \c0.n5182\
        );

    \I__2900\ : InMux
    port map (
            O => \N__17758\,
            I => \N__17755\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__17755\,
            I => \N__17751\
        );

    \I__2898\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17748\
        );

    \I__2897\ : Odrv12
    port map (
            O => \N__17751\,
            I => \c0.n5147\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__17748\,
            I => \c0.n5147\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__17743\,
            I => \c0.n5182_cascade_\
        );

    \I__2894\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17737\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__17737\,
            I => \c0.n40\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__17734\,
            I => \N__17729\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__17733\,
            I => \N__17726\
        );

    \I__2890\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17722\
        );

    \I__2889\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17717\
        );

    \I__2888\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17717\
        );

    \I__2887\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17714\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__17722\,
            I => \N__17711\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__17717\,
            I => \N__17708\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__17714\,
            I => \c0.data_in_field_119\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__17711\,
            I => \c0.data_in_field_119\
        );

    \I__2882\ : Odrv12
    port map (
            O => \N__17708\,
            I => \c0.data_in_field_119\
        );

    \I__2881\ : InMux
    port map (
            O => \N__17701\,
            I => \N__17698\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__17698\,
            I => \c0.n29\
        );

    \I__2879\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17692\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17689\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__17689\,
            I => \c0.n20_adj_1906\
        );

    \I__2876\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17682\
        );

    \I__2875\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17679\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__17682\,
            I => \N__17676\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__17679\,
            I => \N__17673\
        );

    \I__2872\ : Span4Mux_v
    port map (
            O => \N__17676\,
            I => \N__17670\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__17673\,
            I => \N__17666\
        );

    \I__2870\ : Span4Mux_v
    port map (
            O => \N__17670\,
            I => \N__17663\
        );

    \I__2869\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17660\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__17666\,
            I => data_in_4_3
        );

    \I__2867\ : Odrv4
    port map (
            O => \N__17663\,
            I => data_in_4_3
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__17660\,
            I => data_in_4_3
        );

    \I__2865\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17647\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__17647\,
            I => \N__17644\
        );

    \I__2862\ : Span4Mux_s1_h
    port map (
            O => \N__17644\,
            I => \N__17641\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__17641\,
            I => \c0.n15_adj_1894\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \c0.n16_adj_1893_cascade_\
        );

    \I__2859\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17632\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17629\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__17629\,
            I => \c0.n22_adj_1930\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__17626\,
            I => \N__17623\
        );

    \I__2855\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17620\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__17617\,
            I => \c0.n2058\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__17614\,
            I => \c0.n5096_cascade_\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__17611\,
            I => \c0.n1785_cascade_\
        );

    \I__2850\ : InMux
    port map (
            O => \N__17608\,
            I => \N__17605\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__17605\,
            I => \N__17602\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__17602\,
            I => \c0.n22\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__17599\,
            I => \N__17596\
        );

    \I__2846\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17591\
        );

    \I__2845\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17588\
        );

    \I__2844\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17585\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__17591\,
            I => data_in_13_5
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__17588\,
            I => data_in_13_5
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__17585\,
            I => data_in_13_5
        );

    \I__2840\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17575\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__17575\,
            I => \N__17572\
        );

    \I__2838\ : Sp12to4
    port map (
            O => \N__17572\,
            I => \N__17569\
        );

    \I__2837\ : Odrv12
    port map (
            O => \N__17569\,
            I => \c0.n5150\
        );

    \I__2836\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17563\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__17563\,
            I => \N__17556\
        );

    \I__2834\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17547\
        );

    \I__2833\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17547\
        );

    \I__2832\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17547\
        );

    \I__2831\ : InMux
    port map (
            O => \N__17559\,
            I => \N__17547\
        );

    \I__2830\ : Odrv12
    port map (
            O => \N__17556\,
            I => \c0.data_in_field_109\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__17547\,
            I => \c0.data_in_field_109\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__17542\,
            I => \c0.n26_adj_1915_cascade_\
        );

    \I__2827\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17536\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__17536\,
            I => \N__17531\
        );

    \I__2825\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17528\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__17534\,
            I => \N__17525\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__17531\,
            I => \N__17522\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17519\
        );

    \I__2821\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17516\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__17522\,
            I => data_in_17_3
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__17519\,
            I => data_in_17_3
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__17516\,
            I => data_in_17_3
        );

    \I__2817\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17503\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__17508\,
            I => \N__17500\
        );

    \I__2815\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17496\
        );

    \I__2814\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17493\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__17503\,
            I => \N__17490\
        );

    \I__2812\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17487\
        );

    \I__2811\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17484\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__17496\,
            I => \N__17481\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__17493\,
            I => \N__17478\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__17490\,
            I => \N__17473\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__17487\,
            I => \N__17473\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__17484\,
            I => \c0.data_in_field_71\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__17481\,
            I => \c0.data_in_field_71\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__17478\,
            I => \c0.data_in_field_71\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__17473\,
            I => \c0.data_in_field_71\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__17464\,
            I => \c0.n26_cascade_\
        );

    \I__2801\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17458\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__17458\,
            I => \c0.n27_adj_1919\
        );

    \I__2799\ : InMux
    port map (
            O => \N__17455\,
            I => \N__17452\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__17452\,
            I => \c0.n5250\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__17449\,
            I => \c0.n28_adj_1917_cascade_\
        );

    \I__2796\ : InMux
    port map (
            O => \N__17446\,
            I => \N__17443\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__17443\,
            I => \c0.n26_adj_1939\
        );

    \I__2794\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17437\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17432\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__17436\,
            I => \N__17429\
        );

    \I__2791\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17426\
        );

    \I__2790\ : Span4Mux_v
    port map (
            O => \N__17432\,
            I => \N__17423\
        );

    \I__2789\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17418\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__17426\,
            I => \N__17413\
        );

    \I__2787\ : Span4Mux_h
    port map (
            O => \N__17423\,
            I => \N__17413\
        );

    \I__2786\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17408\
        );

    \I__2785\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17408\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__17418\,
            I => \c0.data_in_field_41\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__17413\,
            I => \c0.data_in_field_41\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__17408\,
            I => \c0.data_in_field_41\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \c0.n14_cascade_\
        );

    \I__2780\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17394\
        );

    \I__2779\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17391\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__17394\,
            I => \c0.data_in_frame_18_2\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__17391\,
            I => \c0.data_in_frame_18_2\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__17386\,
            I => \N__17383\
        );

    \I__2775\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17380\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__17380\,
            I => \N__17377\
        );

    \I__2773\ : Span4Mux_h
    port map (
            O => \N__17377\,
            I => \N__17374\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__17374\,
            I => \c0.n5965\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__17371\,
            I => \N__17367\
        );

    \I__2770\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17364\
        );

    \I__2769\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17361\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__17364\,
            I => \N__17356\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__17361\,
            I => \N__17353\
        );

    \I__2766\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17350\
        );

    \I__2765\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17347\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__17356\,
            I => \N__17344\
        );

    \I__2763\ : Span4Mux_v
    port map (
            O => \N__17353\,
            I => \N__17341\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__17350\,
            I => data_in_19_6
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__17347\,
            I => data_in_19_6
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__17344\,
            I => data_in_19_6
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__17341\,
            I => data_in_19_6
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__17332\,
            I => \c0.n22_adj_1901_cascade_\
        );

    \I__2757\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17326\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__17326\,
            I => \c0.n23_adj_1932\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__17323\,
            I => \c0.n30_adj_1940_cascade_\
        );

    \I__2754\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17310\
        );

    \I__2753\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17310\
        );

    \I__2752\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17310\
        );

    \I__2751\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17307\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__17310\,
            I => \c0.n3563\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__17307\,
            I => \c0.n3563\
        );

    \I__2748\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17299\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__17299\,
            I => \c0.n5280\
        );

    \I__2746\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17293\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__17293\,
            I => \c0.n5277\
        );

    \I__2744\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17287\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__17287\,
            I => \c0.n25_adj_1941\
        );

    \I__2742\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17281\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__17281\,
            I => \N__17278\
        );

    \I__2740\ : Span4Mux_h
    port map (
            O => \N__17278\,
            I => \N__17274\
        );

    \I__2739\ : InMux
    port map (
            O => \N__17277\,
            I => \N__17271\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__17274\,
            I => \c0.n5072\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__17271\,
            I => \c0.n5072\
        );

    \I__2736\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17260\
        );

    \I__2735\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17260\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__17260\,
            I => \r_Tx_Data_3\
        );

    \I__2733\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17253\
        );

    \I__2732\ : InMux
    port map (
            O => \N__17256\,
            I => \N__17250\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__17253\,
            I => \N__17247\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__17250\,
            I => \r_Tx_Data_2\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__17247\,
            I => \r_Tx_Data_2\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__17242\,
            I => \N__17239\
        );

    \I__2727\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17230\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__17238\,
            I => \N__17227\
        );

    \I__2725\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17224\
        );

    \I__2724\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17221\
        );

    \I__2723\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17218\
        );

    \I__2722\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17215\
        );

    \I__2721\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17212\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__17230\,
            I => \N__17209\
        );

    \I__2719\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17206\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__17224\,
            I => \r_Bit_Index_1\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__17221\,
            I => \r_Bit_Index_1\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__17218\,
            I => \r_Bit_Index_1\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__17215\,
            I => \r_Bit_Index_1\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__17212\,
            I => \r_Bit_Index_1\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__17209\,
            I => \r_Bit_Index_1\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__17206\,
            I => \r_Bit_Index_1\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__17191\,
            I => \N__17187\
        );

    \I__2710\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17180\
        );

    \I__2709\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17173\
        );

    \I__2708\ : InMux
    port map (
            O => \N__17186\,
            I => \N__17173\
        );

    \I__2707\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17173\
        );

    \I__2706\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17170\
        );

    \I__2705\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17167\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__17180\,
            I => \r_Bit_Index_0\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__17173\,
            I => \r_Bit_Index_0\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__17170\,
            I => \r_Bit_Index_0\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__17167\,
            I => \r_Bit_Index_0\
        );

    \I__2700\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17155\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__17155\,
            I => \c0.tx.n5719\
        );

    \I__2698\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17147\
        );

    \I__2697\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17144\
        );

    \I__2696\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17141\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__17147\,
            I => \r_Bit_Index_2\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__17144\,
            I => \r_Bit_Index_2\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__17141\,
            I => \r_Bit_Index_2\
        );

    \I__2692\ : InMux
    port map (
            O => \N__17134\,
            I => \N__17131\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__17131\,
            I => \c0.tx.n5716\
        );

    \I__2690\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__17125\,
            I => \c0.tx.n5722\
        );

    \I__2688\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17111\
        );

    \I__2687\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17111\
        );

    \I__2686\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17104\
        );

    \I__2685\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17104\
        );

    \I__2684\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17104\
        );

    \I__2683\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17101\
        );

    \I__2682\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17094\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__17111\,
            I => \N__17091\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__17104\,
            I => \N__17086\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__17101\,
            I => \N__17086\
        );

    \I__2678\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17081\
        );

    \I__2677\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17081\
        );

    \I__2676\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17076\
        );

    \I__2675\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17076\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__17094\,
            I => \r_SM_Main_1\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__17091\,
            I => \r_SM_Main_1\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__17086\,
            I => \r_SM_Main_1\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__17081\,
            I => \r_SM_Main_1\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__17076\,
            I => \r_SM_Main_1\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__17065\,
            I => \c0.tx.o_Tx_Serial_N_1798_cascade_\
        );

    \I__2668\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17055\
        );

    \I__2667\ : InMux
    port map (
            O => \N__17061\,
            I => \N__17052\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17046\
        );

    \I__2665\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17041\
        );

    \I__2664\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17038\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__17055\,
            I => \N__17035\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__17052\,
            I => \N__17032\
        );

    \I__2661\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17029\
        );

    \I__2660\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17026\
        );

    \I__2659\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17017\
        );

    \I__2658\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17017\
        );

    \I__2657\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17017\
        );

    \I__2656\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17017\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__17041\,
            I => \r_SM_Main_0\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__17038\,
            I => \r_SM_Main_0\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__17035\,
            I => \r_SM_Main_0\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__17032\,
            I => \r_SM_Main_0\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__17029\,
            I => \r_SM_Main_0\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__17026\,
            I => \r_SM_Main_0\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__17017\,
            I => \r_SM_Main_0\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__17002\,
            I => \N__16993\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__17001\,
            I => \N__16989\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16986\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__16999\,
            I => \N__16980\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__16998\,
            I => \N__16974\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__16997\,
            I => \N__16969\
        );

    \I__2642\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16962\
        );

    \I__2641\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16962\
        );

    \I__2640\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16959\
        );

    \I__2639\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16950\
        );

    \I__2638\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16950\
        );

    \I__2637\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16950\
        );

    \I__2636\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16950\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__16983\,
            I => \N__16946\
        );

    \I__2634\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16937\
        );

    \I__2633\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16937\
        );

    \I__2632\ : InMux
    port map (
            O => \N__16978\,
            I => \N__16937\
        );

    \I__2631\ : InMux
    port map (
            O => \N__16977\,
            I => \N__16937\
        );

    \I__2630\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16932\
        );

    \I__2629\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16932\
        );

    \I__2628\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16923\
        );

    \I__2627\ : InMux
    port map (
            O => \N__16969\,
            I => \N__16923\
        );

    \I__2626\ : InMux
    port map (
            O => \N__16968\,
            I => \N__16923\
        );

    \I__2625\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16923\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__16962\,
            I => \N__16920\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16959\,
            I => \N__16915\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__16950\,
            I => \N__16915\
        );

    \I__2621\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16912\
        );

    \I__2620\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16909\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__16937\,
            I => \r_SM_Main_2\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__16932\,
            I => \r_SM_Main_2\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__16923\,
            I => \r_SM_Main_2\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__16920\,
            I => \r_SM_Main_2\
        );

    \I__2615\ : Odrv12
    port map (
            O => \N__16915\,
            I => \r_SM_Main_2\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__16912\,
            I => \r_SM_Main_2\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__16909\,
            I => \r_SM_Main_2\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__16894\,
            I => \c0.tx.n3_cascade_\
        );

    \I__2611\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16887\
        );

    \I__2610\ : IoInMux
    port map (
            O => \N__16890\,
            I => \N__16884\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__16887\,
            I => \N__16879\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__16884\,
            I => \N__16879\
        );

    \I__2607\ : Span4Mux_s3_v
    port map (
            O => \N__16879\,
            I => \N__16876\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__16876\,
            I => \N__16873\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__16873\,
            I => \N__16870\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__16870\,
            I => \N__16866\
        );

    \I__2603\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16863\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__16866\,
            I => tx_o
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__16863\,
            I => tx_o
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__16858\,
            I => \N__16855\
        );

    \I__2599\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16852\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__16852\,
            I => \c0.n2018\
        );

    \I__2597\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16846\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__16846\,
            I => \c0.n5519\
        );

    \I__2595\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16840\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__16840\,
            I => \N__16837\
        );

    \I__2593\ : Span4Mux_h
    port map (
            O => \N__16837\,
            I => \N__16834\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__16834\,
            I => \c0.n5980\
        );

    \I__2591\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16828\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__16828\,
            I => \N__16824\
        );

    \I__2589\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16821\
        );

    \I__2588\ : Span4Mux_h
    port map (
            O => \N__16824\,
            I => \N__16818\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__16821\,
            I => \r_Tx_Data_4\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__16818\,
            I => \r_Tx_Data_4\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__16813\,
            I => \c0.tx.n5713_cascade_\
        );

    \I__2584\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16804\
        );

    \I__2583\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16801\
        );

    \I__2582\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16798\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16793\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__16804\,
            I => \N__16790\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__16801\,
            I => \N__16787\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__16798\,
            I => \N__16784\
        );

    \I__2577\ : InMux
    port map (
            O => \N__16797\,
            I => \N__16779\
        );

    \I__2576\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16779\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__16793\,
            I => \N__16770\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__16790\,
            I => \N__16770\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__16787\,
            I => \N__16770\
        );

    \I__2572\ : Span4Mux_v
    port map (
            O => \N__16784\,
            I => \N__16770\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__16779\,
            I => data_out_11_1
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__16770\,
            I => data_out_11_1
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__16765\,
            I => \N__16762\
        );

    \I__2568\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16759\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__16759\,
            I => \c0.n9_adj_1880\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__16756\,
            I => \N__16753\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16750\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__16750\,
            I => \N__16747\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__16747\,
            I => \c0.n9_adj_1890\
        );

    \I__2562\ : InMux
    port map (
            O => \N__16744\,
            I => \N__16741\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__16741\,
            I => \N__16738\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__16738\,
            I => \c0.n5489\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__16735\,
            I => \c0.n991_cascade_\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__16732\,
            I => \tx_data_5_N_keep_cascade_\
        );

    \I__2557\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16723\
        );

    \I__2556\ : InMux
    port map (
            O => \N__16728\,
            I => \N__16723\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__16723\,
            I => \r_Tx_Data_5\
        );

    \I__2554\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16717\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16714\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__16714\,
            I => \tx_data_3_N_keep\
        );

    \I__2551\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16707\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__16710\,
            I => \N__16704\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__16707\,
            I => \N__16700\
        );

    \I__2548\ : InMux
    port map (
            O => \N__16704\,
            I => \N__16695\
        );

    \I__2547\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16695\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__16700\,
            I => n5135
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__16695\,
            I => n5135
        );

    \I__2544\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16687\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__16687\,
            I => n5117
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__16684\,
            I => \n5117_cascade_\
        );

    \I__2541\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16674\
        );

    \I__2540\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16658\
        );

    \I__2539\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16658\
        );

    \I__2538\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16655\
        );

    \I__2537\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16652\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__16674\,
            I => \N__16649\
        );

    \I__2535\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16646\
        );

    \I__2534\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16643\
        );

    \I__2533\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16640\
        );

    \I__2532\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16631\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16631\
        );

    \I__2530\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16631\
        );

    \I__2529\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16631\
        );

    \I__2528\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16626\
        );

    \I__2527\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16626\
        );

    \I__2526\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16621\
        );

    \I__2525\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16621\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__16658\,
            I => n4316
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__16655\,
            I => n4316
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__16652\,
            I => n4316
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__16649\,
            I => n4316
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__16646\,
            I => n4316
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__16643\,
            I => n4316
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__16640\,
            I => n4316
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__16631\,
            I => n4316
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__16626\,
            I => n4316
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__16621\,
            I => n4316
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__16600\,
            I => \N__16596\
        );

    \I__2513\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16591\
        );

    \I__2512\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16591\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16591\,
            I => data_out_19_5
        );

    \I__2510\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16585\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__16585\,
            I => \tx_data_2_N_keep\
        );

    \I__2508\ : InMux
    port map (
            O => \N__16582\,
            I => \N__16576\
        );

    \I__2507\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16571\
        );

    \I__2506\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16571\
        );

    \I__2505\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16567\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__16576\,
            I => \N__16562\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16559\
        );

    \I__2502\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16555\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__16567\,
            I => \N__16552\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__16566\,
            I => \N__16549\
        );

    \I__2499\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16546\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__16562\,
            I => \N__16541\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__16559\,
            I => \N__16541\
        );

    \I__2496\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16538\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__16555\,
            I => \N__16533\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__16552\,
            I => \N__16533\
        );

    \I__2493\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16530\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__16546\,
            I => data_out_11_3
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__16541\,
            I => data_out_11_3
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__16538\,
            I => data_out_11_3
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__16533\,
            I => data_out_11_3
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__16530\,
            I => data_out_11_3
        );

    \I__2487\ : InMux
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__16516\,
            I => \N__16509\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__16515\,
            I => \N__16506\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__16514\,
            I => \N__16503\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__16513\,
            I => \N__16500\
        );

    \I__2482\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16497\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__16509\,
            I => \N__16494\
        );

    \I__2480\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16489\
        );

    \I__2479\ : InMux
    port map (
            O => \N__16503\,
            I => \N__16489\
        );

    \I__2478\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16486\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__16497\,
            I => data_out_11_2
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__16494\,
            I => data_out_11_2
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__16489\,
            I => data_out_11_2
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__16486\,
            I => data_out_11_2
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__16477\,
            I => \c0.n1805_cascade_\
        );

    \I__2472\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16471\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__16471\,
            I => \N__16466\
        );

    \I__2470\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16463\
        );

    \I__2469\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16460\
        );

    \I__2468\ : Span4Mux_h
    port map (
            O => \N__16466\,
            I => \N__16457\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__16463\,
            I => n135
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__16460\,
            I => n135
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__16457\,
            I => n135
        );

    \I__2464\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16447\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__16447\,
            I => \c0.n1805\
        );

    \I__2462\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16441\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__16441\,
            I => \N__16438\
        );

    \I__2460\ : Odrv12
    port map (
            O => \N__16438\,
            I => n5173
        );

    \I__2459\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16427\
        );

    \I__2458\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16420\
        );

    \I__2457\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16420\
        );

    \I__2456\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16420\
        );

    \I__2455\ : InMux
    port map (
            O => \N__16431\,
            I => \N__16417\
        );

    \I__2454\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16412\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__16427\,
            I => \N__16407\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__16420\,
            I => \N__16407\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__16417\,
            I => \N__16404\
        );

    \I__2450\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16401\
        );

    \I__2449\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16398\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__16412\,
            I => \N__16395\
        );

    \I__2447\ : Span4Mux_v
    port map (
            O => \N__16407\,
            I => \N__16392\
        );

    \I__2446\ : Span4Mux_s2_h
    port map (
            O => \N__16404\,
            I => \N__16389\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__16401\,
            I => data_out_11_7
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__16398\,
            I => data_out_11_7
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__16395\,
            I => data_out_11_7
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__16392\,
            I => data_out_11_7
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__16389\,
            I => data_out_11_7
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__16378\,
            I => \N__16375\
        );

    \I__2439\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16372\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16367\
        );

    \I__2437\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16364\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \N__16360\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__16367\,
            I => \N__16355\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__16364\,
            I => \N__16355\
        );

    \I__2433\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16351\
        );

    \I__2432\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16348\
        );

    \I__2431\ : Span4Mux_v
    port map (
            O => \N__16355\,
            I => \N__16345\
        );

    \I__2430\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16341\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__16351\,
            I => \N__16338\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__16348\,
            I => \N__16335\
        );

    \I__2427\ : Span4Mux_s1_h
    port map (
            O => \N__16345\,
            I => \N__16332\
        );

    \I__2426\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16329\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__16341\,
            I => data_out_10_7
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__16338\,
            I => data_out_10_7
        );

    \I__2423\ : Odrv12
    port map (
            O => \N__16335\,
            I => data_out_10_7
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__16332\,
            I => data_out_10_7
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__16329\,
            I => data_out_10_7
        );

    \I__2420\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16315\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__16315\,
            I => \N__16312\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__16312\,
            I => n5079
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16305\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__16308\,
            I => \N__16302\
        );

    \I__2415\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16299\
        );

    \I__2414\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16296\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__16299\,
            I => data_out_19_1
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__16296\,
            I => data_out_19_1
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__16291\,
            I => \N__16288\
        );

    \I__2410\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16285\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__16285\,
            I => \N__16280\
        );

    \I__2408\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16277\
        );

    \I__2407\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16274\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__16280\,
            I => \N__16264\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__16277\,
            I => \N__16264\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__16274\,
            I => \N__16264\
        );

    \I__2403\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16261\
        );

    \I__2402\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16256\
        );

    \I__2401\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16256\
        );

    \I__2400\ : Span4Mux_h
    port map (
            O => \N__16264\,
            I => \N__16253\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__16261\,
            I => data_out_11_0
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__16256\,
            I => data_out_11_0
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__16253\,
            I => data_out_11_0
        );

    \I__2396\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16242\
        );

    \I__2395\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16239\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__16242\,
            I => data_out_18_2
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__16239\,
            I => data_out_18_2
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__16234\,
            I => \N__16231\
        );

    \I__2391\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16228\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__16228\,
            I => \N__16224\
        );

    \I__2389\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16221\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__16224\,
            I => \N__16218\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__16221\,
            I => data_out_19_2
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__16218\,
            I => data_out_19_2
        );

    \I__2385\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__16210\,
            I => \c0.n2249\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__16207\,
            I => \c0.n5522_cascade_\
        );

    \I__2382\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__16201\,
            I => n4_adj_1991
        );

    \I__2380\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16194\
        );

    \I__2379\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__16194\,
            I => data_out_18_5
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__16191\,
            I => data_out_18_5
        );

    \I__2376\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16183\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__16183\,
            I => \N__16180\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__16180\,
            I => n4_adj_1994
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__16177\,
            I => \c0.rx.n2151_cascade_\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__16174\,
            I => \n1709_cascade_\
        );

    \I__2371\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16167\
        );

    \I__2370\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16164\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__16167\,
            I => \N__16161\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__16164\,
            I => n4_adj_1990
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__16161\,
            I => n4_adj_1990
        );

    \I__2366\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16152\
        );

    \I__2365\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16149\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__16152\,
            I => rx_data_4
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__16149\,
            I => rx_data_4
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__16144\,
            I => \N__16141\
        );

    \I__2361\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16138\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__16138\,
            I => \N__16135\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__16135\,
            I => \N__16132\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__16132\,
            I => n4_adj_1992
        );

    \I__2357\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16126\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__16126\,
            I => \N__16122\
        );

    \I__2355\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16119\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__16122\,
            I => \N__16116\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__16119\,
            I => \c0.data_in_frame_18_6\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__16116\,
            I => \c0.data_in_frame_18_6\
        );

    \I__2351\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16108\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__16108\,
            I => \N__16104\
        );

    \I__2349\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16099\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__16104\,
            I => \N__16096\
        );

    \I__2347\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16091\
        );

    \I__2346\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16091\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__16099\,
            I => data_in_2_5
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__16096\,
            I => data_in_2_5
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__16091\,
            I => data_in_2_5
        );

    \I__2342\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16081\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__16081\,
            I => \N__16077\
        );

    \I__2340\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16074\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__16077\,
            I => rx_data_6
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__16074\,
            I => rx_data_6
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__16069\,
            I => \c0.n5222_cascade_\
        );

    \I__2336\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__16063\,
            I => \c0.n42\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__16060\,
            I => \c0.n33_cascade_\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__16057\,
            I => \c0.n2008_cascade_\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \c0.n38_cascade_\
        );

    \I__2331\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16048\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__16048\,
            I => \N__16045\
        );

    \I__2329\ : Span4Mux_s3_h
    port map (
            O => \N__16045\,
            I => \N__16042\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__16042\,
            I => \c0.n5462\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__16039\,
            I => \N__16036\
        );

    \I__2326\ : InMux
    port map (
            O => \N__16036\,
            I => \N__16030\
        );

    \I__2325\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16030\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16026\
        );

    \I__2323\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16023\
        );

    \I__2322\ : Span4Mux_s3_h
    port map (
            O => \N__16026\,
            I => \N__16020\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__16023\,
            I => data_in_12_5
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__16020\,
            I => data_in_12_5
        );

    \I__2319\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16012\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__16012\,
            I => \N__16008\
        );

    \I__2317\ : InMux
    port map (
            O => \N__16011\,
            I => \N__16005\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__16008\,
            I => \N__16002\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__16005\,
            I => \c0.data_in_frame_18_0\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__16002\,
            I => \c0.data_in_frame_18_0\
        );

    \I__2313\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15994\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__15994\,
            I => \N__15990\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15987\
        );

    \I__2310\ : Span4Mux_s3_h
    port map (
            O => \N__15990\,
            I => \N__15984\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__15987\,
            I => \c0.data_in_frame_18_4\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__15984\,
            I => \c0.data_in_frame_18_4\
        );

    \I__2307\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15976\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__15976\,
            I => \c0.n22_adj_1881\
        );

    \I__2305\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__15970\,
            I => \c0.n5266\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__2302\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15960\
        );

    \I__2301\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15955\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__15960\,
            I => \N__15952\
        );

    \I__2299\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15949\
        );

    \I__2298\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15946\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15941\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__15952\,
            I => \N__15941\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15938\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__15946\,
            I => \N__15935\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__15941\,
            I => \c0.data_in_field_101\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__15938\,
            I => \c0.data_in_field_101\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__15935\,
            I => \c0.data_in_field_101\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__15928\,
            I => \c0.n18_adj_1882_cascade_\
        );

    \I__2289\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15922\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__15922\,
            I => \c0.n26_adj_1883\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__15919\,
            I => \c0.n30_adj_1897_cascade_\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__15916\,
            I => \c0.n36_cascade_\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__15913\,
            I => \c0.n5080_cascade_\
        );

    \I__2284\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15907\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__15907\,
            I => \c0.n1990\
        );

    \I__2282\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15901\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__15901\,
            I => \N__15898\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__15898\,
            I => \c0.n5192\
        );

    \I__2279\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15892\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__15892\,
            I => \c0.n5080\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15886\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__15886\,
            I => \c0.n23_adj_1931\
        );

    \I__2275\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15880\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__15880\,
            I => \c0.n21_adj_1928\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__15877\,
            I => \c0.n22_adj_1927_cascade_\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15871\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__15871\,
            I => \N__15868\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__15868\,
            I => \c0.n24_adj_1907\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__15865\,
            I => \N__15862\
        );

    \I__2268\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15858\
        );

    \I__2267\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15854\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__15858\,
            I => \N__15850\
        );

    \I__2265\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15847\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__15854\,
            I => \N__15844\
        );

    \I__2263\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15841\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__15850\,
            I => \N__15838\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__15847\,
            I => data_in_19_3
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__15844\,
            I => data_in_19_3
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__15841\,
            I => data_in_19_3
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__15838\,
            I => data_in_19_3
        );

    \I__2257\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15826\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__15826\,
            I => \c0.n3414\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__15823\,
            I => \N__15818\
        );

    \I__2254\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15813\
        );

    \I__2253\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15813\
        );

    \I__2252\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15810\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__15813\,
            I => \N__15807\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__15810\,
            I => \N__15804\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__15807\,
            I => \N__15801\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__15804\,
            I => \N__15798\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__15801\,
            I => \c0.FRAME_MATCHER_wait_for_transmission_N_909\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__15798\,
            I => \c0.FRAME_MATCHER_wait_for_transmission_N_909\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__15793\,
            I => \N__15790\
        );

    \I__2244\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15787\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__15787\,
            I => \N__15784\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__15784\,
            I => \N__15777\
        );

    \I__2241\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15772\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15772\
        );

    \I__2239\ : InMux
    port map (
            O => \N__15781\,
            I => \N__15767\
        );

    \I__2238\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15767\
        );

    \I__2237\ : Sp12to4
    port map (
            O => \N__15777\,
            I => \N__15762\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__15772\,
            I => \N__15762\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__15767\,
            I => \c0.r_SM_Main_2_N_1770_0\
        );

    \I__2234\ : Odrv12
    port map (
            O => \N__15762\,
            I => \c0.r_SM_Main_2_N_1770_0\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15753\
        );

    \I__2232\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15750\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__15753\,
            I => \N__15744\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__15750\,
            I => \N__15744\
        );

    \I__2229\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15741\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__15744\,
            I => \N__15738\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__15741\,
            I => tx2_active
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__15738\,
            I => tx2_active
        );

    \I__2225\ : CEMux
    port map (
            O => \N__15733\,
            I => \N__15730\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15727\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__15727\,
            I => \c0.n195\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__15724\,
            I => \c0.n5845_cascade_\
        );

    \I__2221\ : SRMux
    port map (
            O => \N__15721\,
            I => \N__15718\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__15718\,
            I => \N__15715\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__15715\,
            I => \N__15712\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__15712\,
            I => \c0.n2275\
        );

    \I__2217\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15706\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__15706\,
            I => \N__15703\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__2214\ : InMux
    port map (
            O => \N__15702\,
            I => \N__15690\
        );

    \I__2213\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15690\
        );

    \I__2212\ : InMux
    port map (
            O => \N__15700\,
            I => \N__15690\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__15697\,
            I => \c0.data_in_field_81\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__15690\,
            I => \c0.data_in_field_81\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__15685\,
            I => \c0.n1918_cascade_\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__15682\,
            I => \c0.n5192_cascade_\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__15679\,
            I => \c0.tx.n3507_cascade_\
        );

    \I__2206\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15670\
        );

    \I__2205\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15670\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__15670\,
            I => n2307
        );

    \I__2203\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15655\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15655\
        );

    \I__2201\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15655\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15655\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__15655\,
            I => n2200
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__15652\,
            I => \n2307_cascade_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__15649\,
            I => \N__15646\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__15646\,
            I => \N__15643\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__15643\,
            I => n805
        );

    \I__2194\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15634\
        );

    \I__2193\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15634\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15628\
        );

    \I__2191\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15625\
        );

    \I__2190\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15619\
        );

    \I__2189\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15619\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__15628\,
            I => \N__15614\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__15625\,
            I => \N__15614\
        );

    \I__2186\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15611\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__15619\,
            I => \c0.tx2.r_Bit_Index_0\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__15614\,
            I => \c0.tx2.r_Bit_Index_0\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__15611\,
            I => \c0.tx2.r_Bit_Index_0\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__15604\,
            I => \N__15599\
        );

    \I__2181\ : InMux
    port map (
            O => \N__15603\,
            I => \N__15595\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__15602\,
            I => \N__15591\
        );

    \I__2179\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15587\
        );

    \I__2178\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15584\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15581\
        );

    \I__2176\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15576\
        );

    \I__2175\ : InMux
    port map (
            O => \N__15591\,
            I => \N__15576\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__15590\,
            I => \N__15573\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__15587\,
            I => \N__15569\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__15584\,
            I => \N__15566\
        );

    \I__2171\ : Span4Mux_s2_h
    port map (
            O => \N__15581\,
            I => \N__15561\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__15576\,
            I => \N__15561\
        );

    \I__2169\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15556\
        );

    \I__2168\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15556\
        );

    \I__2167\ : Span4Mux_s3_h
    port map (
            O => \N__15569\,
            I => \N__15553\
        );

    \I__2166\ : Span4Mux_s3_h
    port map (
            O => \N__15566\,
            I => \N__15550\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__15561\,
            I => \N__15547\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__15556\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__15553\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__2162\ : Odrv4
    port map (
            O => \N__15550\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__15547\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__2160\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15534\
        );

    \I__2159\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15531\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__15534\,
            I => \N__15527\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__15531\,
            I => \N__15524\
        );

    \I__2156\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15521\
        );

    \I__2155\ : Span4Mux_s3_h
    port map (
            O => \N__15527\,
            I => \N__15518\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__15524\,
            I => \N__15515\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__15521\,
            I => \c0.tx2.r_Bit_Index_2\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__15518\,
            I => \c0.tx2.r_Bit_Index_2\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__15515\,
            I => \c0.tx2.r_Bit_Index_2\
        );

    \I__2150\ : CEMux
    port map (
            O => \N__15508\,
            I => \N__15505\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__15505\,
            I => \N__15502\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__15502\,
            I => \c0.tx2.n2218\
        );

    \I__2147\ : SRMux
    port map (
            O => \N__15499\,
            I => \N__15496\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__15496\,
            I => \c0.tx2.n2319\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__15493\,
            I => \N__15490\
        );

    \I__2144\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15487\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15483\
        );

    \I__2142\ : InMux
    port map (
            O => \N__15486\,
            I => \N__15480\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__15483\,
            I => \N__15477\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__15480\,
            I => \N__15474\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__15477\,
            I => n5153
        );

    \I__2138\ : Odrv12
    port map (
            O => \N__15474\,
            I => n5153
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__15469\,
            I => \c0.n3414_cascade_\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__15466\,
            I => \N__15463\
        );

    \I__2135\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15460\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15457\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__15457\,
            I => \N__15454\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__15454\,
            I => \c0.n9\
        );

    \I__2131\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15448\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__15448\,
            I => \N__15445\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__15445\,
            I => \c0.n5501\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__15442\,
            I => \c0.n1173_cascade_\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__15439\,
            I => \tx_data_0_N_keep_cascade_\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__15436\,
            I => \N__15432\
        );

    \I__2125\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15427\
        );

    \I__2124\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15427\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__15427\,
            I => \r_Tx_Data_0\
        );

    \I__2122\ : InMux
    port map (
            O => \N__15424\,
            I => \N__15421\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__15421\,
            I => \c0.n5531\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__15418\,
            I => \c0.n15_cascade_\
        );

    \I__2119\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15412\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__15409\,
            I => \tx_data_1_N_keep\
        );

    \I__2116\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15393\
        );

    \I__2115\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15393\
        );

    \I__2114\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15393\
        );

    \I__2113\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15393\
        );

    \I__2112\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15390\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__15393\,
            I => \c0.tx.r_SM_Main_2_N_1767_1\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__15390\,
            I => \c0.tx.r_SM_Main_2_N_1767_1\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__15385\,
            I => \N__15382\
        );

    \I__2108\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15379\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__15379\,
            I => \c0.tx.n3507\
        );

    \I__2106\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15373\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__15373\,
            I => n5156
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__15370\,
            I => \N__15367\
        );

    \I__2103\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15364\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__15364\,
            I => \N__15361\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__15361\,
            I => n5063
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__15358\,
            I => \N__15354\
        );

    \I__2099\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15351\
        );

    \I__2098\ : InMux
    port map (
            O => \N__15354\,
            I => \N__15348\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__15351\,
            I => data_out_18_3
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__15348\,
            I => data_out_18_3
        );

    \I__2095\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15339\
        );

    \I__2094\ : InMux
    port map (
            O => \N__15342\,
            I => \N__15336\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__15339\,
            I => \N__15333\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__15336\,
            I => data_out_19_7
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__15333\,
            I => data_out_19_7
        );

    \I__2090\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15325\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__15325\,
            I => \N__15322\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__15322\,
            I => n7_adj_1998
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__15319\,
            I => \N__15316\
        );

    \I__2086\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15313\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__15313\,
            I => n8_adj_1997
        );

    \I__2084\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15304\
        );

    \I__2083\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15304\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__15304\,
            I => data_out_18_7
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__15301\,
            I => \N__15298\
        );

    \I__2080\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15292\
        );

    \I__2079\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15292\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__15292\,
            I => data_out_19_3
        );

    \I__2077\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15285\
        );

    \I__2076\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15282\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__15285\,
            I => \N__15279\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__15282\,
            I => data_out_18_1
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__15279\,
            I => data_out_18_1
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__15274\,
            I => \N__15271\
        );

    \I__2071\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15268\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__15268\,
            I => n4_adj_2007
        );

    \I__2069\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15261\
        );

    \I__2068\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__15261\,
            I => \N__15255\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__15258\,
            I => \r_Tx_Data_1\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__15255\,
            I => \r_Tx_Data_1\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__15250\,
            I => \N__15246\
        );

    \I__2063\ : InMux
    port map (
            O => \N__15249\,
            I => \N__15243\
        );

    \I__2062\ : InMux
    port map (
            O => \N__15246\,
            I => \N__15240\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__15243\,
            I => data_out_19_0
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__15240\,
            I => data_out_19_0
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__15235\,
            I => \N__15232\
        );

    \I__2058\ : InMux
    port map (
            O => \N__15232\,
            I => \N__15226\
        );

    \I__2057\ : InMux
    port map (
            O => \N__15231\,
            I => \N__15226\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__15226\,
            I => \c0.delay_counter_9\
        );

    \I__2055\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15219\
        );

    \I__2054\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15216\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__15219\,
            I => \c0.delay_counter_2\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__15216\,
            I => \c0.delay_counter_2\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__15211\,
            I => \N__15207\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__15210\,
            I => \N__15204\
        );

    \I__2049\ : InMux
    port map (
            O => \N__15207\,
            I => \N__15201\
        );

    \I__2048\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15198\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__15201\,
            I => \c0.delay_counter_0\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__15198\,
            I => \c0.delay_counter_0\
        );

    \I__2045\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15189\
        );

    \I__2044\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15186\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__15189\,
            I => \c0.delay_counter_7\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__15186\,
            I => \c0.delay_counter_7\
        );

    \I__2041\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15178\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__15178\,
            I => \c0.n18_adj_1908\
        );

    \I__2039\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15172\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__15172\,
            I => \N__15169\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__15169\,
            I => n4_adj_2000
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__15166\,
            I => \n5086_cascade_\
        );

    \I__2035\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15159\
        );

    \I__2034\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15156\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__15159\,
            I => \N__15152\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15149\
        );

    \I__2031\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15146\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__15152\,
            I => \N__15143\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__15149\,
            I => \N__15140\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__15146\,
            I => \N__15137\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__15143\,
            I => n1525
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__15140\,
            I => n1525
        );

    \I__2025\ : Odrv12
    port map (
            O => \N__15137\,
            I => n1525
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__15130\,
            I => \n5156_cascade_\
        );

    \I__2023\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15123\
        );

    \I__2022\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15120\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__15123\,
            I => data_out_18_0
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__15120\,
            I => data_out_18_0
        );

    \I__2019\ : InMux
    port map (
            O => \N__15115\,
            I => \c0.n4406\
        );

    \I__2018\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15108\
        );

    \I__2017\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15105\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__15108\,
            I => \c0.delay_counter_4\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__15105\,
            I => \c0.delay_counter_4\
        );

    \I__2014\ : InMux
    port map (
            O => \N__15100\,
            I => \c0.n4407\
        );

    \I__2013\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15093\
        );

    \I__2012\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15090\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__15093\,
            I => \c0.delay_counter_5\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__15090\,
            I => \c0.delay_counter_5\
        );

    \I__2009\ : InMux
    port map (
            O => \N__15085\,
            I => \c0.n4408\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__15082\,
            I => \N__15078\
        );

    \I__2007\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15075\
        );

    \I__2006\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15072\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__15075\,
            I => \c0.delay_counter_6\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__15072\,
            I => \c0.delay_counter_6\
        );

    \I__2003\ : InMux
    port map (
            O => \N__15067\,
            I => \c0.n4409\
        );

    \I__2002\ : InMux
    port map (
            O => \N__15064\,
            I => \c0.n4410\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__15061\,
            I => \N__15058\
        );

    \I__2000\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15054\
        );

    \I__1999\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15051\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__15054\,
            I => \c0.delay_counter_8\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__15051\,
            I => \c0.delay_counter_8\
        );

    \I__1996\ : InMux
    port map (
            O => \N__15046\,
            I => \bfn_4_17_0_\
        );

    \I__1995\ : InMux
    port map (
            O => \N__15043\,
            I => \c0.n4412\
        );

    \I__1994\ : InMux
    port map (
            O => \N__15040\,
            I => \c0.n4413\
        );

    \I__1993\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15033\
        );

    \I__1992\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15030\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__15033\,
            I => \c0.delay_counter_10\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__15030\,
            I => \c0.delay_counter_10\
        );

    \I__1989\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15022\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__15022\,
            I => \N__15018\
        );

    \I__1987\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15015\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__15018\,
            I => \N__15012\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__15015\,
            I => \N__15009\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__15012\,
            I => n5077
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__15009\,
            I => n5077
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__15004\,
            I => \N__15001\
        );

    \I__1981\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14998\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__14998\,
            I => \N__14995\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__14995\,
            I => n4_adj_1988
        );

    \I__1978\ : CEMux
    port map (
            O => \N__14992\,
            I => \N__14989\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N__14985\
        );

    \I__1976\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14982\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__14985\,
            I => \c0.rx.n2213\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__14982\,
            I => \c0.rx.n2213\
        );

    \I__1973\ : SRMux
    port map (
            O => \N__14977\,
            I => \N__14974\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__14974\,
            I => \N__14971\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__14971\,
            I => \c0.rx.n2317\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14951\
        );

    \I__1969\ : InMux
    port map (
            O => \N__14967\,
            I => \N__14951\
        );

    \I__1968\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14951\
        );

    \I__1967\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14951\
        );

    \I__1966\ : InMux
    port map (
            O => \N__14964\,
            I => \N__14951\
        );

    \I__1965\ : InMux
    port map (
            O => \N__14963\,
            I => \N__14946\
        );

    \I__1964\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14946\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__14951\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__14946\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__14941\,
            I => \N__14935\
        );

    \I__1960\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14924\
        );

    \I__1959\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14924\
        );

    \I__1958\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14924\
        );

    \I__1957\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14924\
        );

    \I__1956\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14919\
        );

    \I__1955\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14919\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__14924\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__14919\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__1952\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14908\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__14913\,
            I => \N__14905\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14912\,
            I => \N__14902\
        );

    \I__1949\ : InMux
    port map (
            O => \N__14911\,
            I => \N__14899\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__14908\,
            I => \N__14896\
        );

    \I__1947\ : InMux
    port map (
            O => \N__14905\,
            I => \N__14893\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__14902\,
            I => \r_Clock_Count_0\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__14899\,
            I => \r_Clock_Count_0\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__14896\,
            I => \r_Clock_Count_0\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__14893\,
            I => \r_Clock_Count_0\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__14884\,
            I => \N__14878\
        );

    \I__1941\ : InMux
    port map (
            O => \N__14883\,
            I => \N__14875\
        );

    \I__1940\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14871\
        );

    \I__1939\ : InMux
    port map (
            O => \N__14881\,
            I => \N__14868\
        );

    \I__1938\ : InMux
    port map (
            O => \N__14878\,
            I => \N__14865\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__14875\,
            I => \N__14862\
        );

    \I__1936\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14859\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__14871\,
            I => \r_Clock_Count_6\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__14868\,
            I => \r_Clock_Count_6\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__14865\,
            I => \r_Clock_Count_6\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__14862\,
            I => \r_Clock_Count_6\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__14859\,
            I => \r_Clock_Count_6\
        );

    \I__1930\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14845\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__14845\,
            I => n8_adj_1996
        );

    \I__1928\ : IoInMux
    port map (
            O => \N__14842\,
            I => \N__14839\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__14839\,
            I => tx_enable
        );

    \I__1926\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14832\
        );

    \I__1925\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14829\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__14832\,
            I => \c0.delay_counter_1\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__14829\,
            I => \c0.delay_counter_1\
        );

    \I__1922\ : InMux
    port map (
            O => \N__14824\,
            I => \c0.n4404\
        );

    \I__1921\ : InMux
    port map (
            O => \N__14821\,
            I => \c0.n4405\
        );

    \I__1920\ : InMux
    port map (
            O => \N__14818\,
            I => \N__14814\
        );

    \I__1919\ : InMux
    port map (
            O => \N__14817\,
            I => \N__14811\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__14814\,
            I => \N__14808\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__14811\,
            I => \c0.delay_counter_3\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__14808\,
            I => \c0.delay_counter_3\
        );

    \I__1915\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14800\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__14800\,
            I => \c0.n5671\
        );

    \I__1913\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14794\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14790\
        );

    \I__1911\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14787\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__14790\,
            I => rx_data_3
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__14787\,
            I => rx_data_3
        );

    \I__1908\ : InMux
    port map (
            O => \N__14782\,
            I => \N__14779\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__14779\,
            I => \N__14775\
        );

    \I__1906\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14772\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__14775\,
            I => rx_data_5
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__14772\,
            I => rx_data_5
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__14767\,
            I => \N__14762\
        );

    \I__1902\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14757\
        );

    \I__1901\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14754\
        );

    \I__1900\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14751\
        );

    \I__1899\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14746\
        );

    \I__1898\ : InMux
    port map (
            O => \N__14760\,
            I => \N__14746\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__14757\,
            I => \N__14743\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__14754\,
            I => \N__14740\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__14751\,
            I => \r_Clock_Count_7_adj_2004\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__14746\,
            I => \r_Clock_Count_7_adj_2004\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__14743\,
            I => \r_Clock_Count_7_adj_2004\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__14740\,
            I => \r_Clock_Count_7_adj_2004\
        );

    \I__1891\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14726\
        );

    \I__1890\ : InMux
    port map (
            O => \N__14730\,
            I => \N__14721\
        );

    \I__1889\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14718\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14715\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14710\
        );

    \I__1886\ : InMux
    port map (
            O => \N__14724\,
            I => \N__14710\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__14721\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__14718\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__14715\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__14710\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__1881\ : InMux
    port map (
            O => \N__14701\,
            I => \N__14698\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__14695\,
            I => \c0.rx.n6\
        );

    \I__1878\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14686\
        );

    \I__1877\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14683\
        );

    \I__1876\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14678\
        );

    \I__1875\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14678\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__14686\,
            I => \c0.data_in_field_131\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__14683\,
            I => \c0.data_in_field_131\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__14678\,
            I => \c0.data_in_field_131\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__14671\,
            I => \c0.n2036_cascade_\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__14668\,
            I => \c0.n5273_cascade_\
        );

    \I__1869\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14662\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14658\
        );

    \I__1867\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14655\
        );

    \I__1866\ : Span4Mux_s3_h
    port map (
            O => \N__14658\,
            I => \N__14652\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__14655\,
            I => \c0.data_in_frame_18_7\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__14652\,
            I => \c0.data_in_frame_18_7\
        );

    \I__1863\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14643\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__14646\,
            I => \N__14640\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__14643\,
            I => \N__14636\
        );

    \I__1860\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14630\
        );

    \I__1859\ : InMux
    port map (
            O => \N__14639\,
            I => \N__14630\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__14636\,
            I => \N__14627\
        );

    \I__1857\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14624\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__14630\,
            I => data_in_18_3
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__14627\,
            I => data_in_18_3
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__14624\,
            I => data_in_18_3
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__14617\,
            I => \c0.n1893_cascade_\
        );

    \I__1852\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14611\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__14611\,
            I => \c0.n20_adj_1921\
        );

    \I__1850\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14605\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__14605\,
            I => \c0.n5459\
        );

    \I__1848\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14599\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__14599\,
            I => \N__14596\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__14596\,
            I => \c0.n5737\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__14593\,
            I => \N__14590\
        );

    \I__1844\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14583\
        );

    \I__1842\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14580\
        );

    \I__1841\ : Span12Mux_s2_h
    port map (
            O => \N__14583\,
            I => \N__14577\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__14580\,
            I => \c0.data_in_frame_19_1\
        );

    \I__1839\ : Odrv12
    port map (
            O => \N__14577\,
            I => \c0.data_in_frame_19_1\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__14572\,
            I => \N__14569\
        );

    \I__1837\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14566\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__14566\,
            I => \N__14563\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__14563\,
            I => \c0.n5944\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \N__14556\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__14559\,
            I => \N__14553\
        );

    \I__1832\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14550\
        );

    \I__1831\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14547\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__14550\,
            I => \c0.data_in_frame_19_6\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__14547\,
            I => \c0.data_in_frame_19_6\
        );

    \I__1828\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__14539\,
            I => \c0.n5456\
        );

    \I__1826\ : InMux
    port map (
            O => \N__14536\,
            I => \c0.n4403\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__14533\,
            I => \N__14527\
        );

    \I__1824\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14518\
        );

    \I__1823\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14518\
        );

    \I__1822\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14518\
        );

    \I__1821\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14515\
        );

    \I__1820\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14512\
        );

    \I__1819\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14506\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14500\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__14515\,
            I => \N__14500\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__14512\,
            I => \N__14497\
        );

    \I__1815\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14490\
        );

    \I__1814\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14490\
        );

    \I__1813\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14490\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__14506\,
            I => \N__14487\
        );

    \I__1811\ : InMux
    port map (
            O => \N__14505\,
            I => \N__14484\
        );

    \I__1810\ : Span4Mux_s3_h
    port map (
            O => \N__14500\,
            I => \N__14481\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__14497\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__14490\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__14487\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__14484\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__14481\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__14470\,
            I => \c0.n5785_cascade_\
        );

    \I__1803\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14464\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__14464\,
            I => \N__14461\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__14461\,
            I => \c0.n5426\
        );

    \I__1800\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14455\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__14455\,
            I => \c0.n5788\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__14452\,
            I => \N__14449\
        );

    \I__1797\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14446\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__14446\,
            I => \c0.n5968\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14440\
        );

    \I__1794\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14437\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14434\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__14434\,
            I => \c0.n5363\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__14431\,
            I => \N__14428\
        );

    \I__1790\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14424\
        );

    \I__1789\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14421\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__14424\,
            I => \N__14418\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__14421\,
            I => \N__14415\
        );

    \I__1786\ : Span4Mux_s2_h
    port map (
            O => \N__14418\,
            I => \N__14412\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__14415\,
            I => \c0.data_in_frame_19_7\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__14412\,
            I => \c0.data_in_frame_19_7\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__14407\,
            I => \N__14404\
        );

    \I__1782\ : InMux
    port map (
            O => \N__14404\,
            I => \N__14401\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__14401\,
            I => \c0.n5935\
        );

    \I__1780\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14394\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__14397\,
            I => \N__14382\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__14394\,
            I => \N__14379\
        );

    \I__1777\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14372\
        );

    \I__1776\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14372\
        );

    \I__1775\ : InMux
    port map (
            O => \N__14391\,
            I => \N__14372\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__14390\,
            I => \N__14369\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__14389\,
            I => \N__14365\
        );

    \I__1772\ : InMux
    port map (
            O => \N__14388\,
            I => \N__14362\
        );

    \I__1771\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14353\
        );

    \I__1770\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14353\
        );

    \I__1769\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14353\
        );

    \I__1768\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14353\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__14379\,
            I => \N__14350\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__14372\,
            I => \N__14347\
        );

    \I__1765\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14344\
        );

    \I__1764\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14339\
        );

    \I__1763\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14339\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__14362\,
            I => \r_SM_Main_1_adj_2010\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__14353\,
            I => \r_SM_Main_1_adj_2010\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__14350\,
            I => \r_SM_Main_1_adj_2010\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__14347\,
            I => \r_SM_Main_1_adj_2010\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__14344\,
            I => \r_SM_Main_1_adj_2010\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__14339\,
            I => \r_SM_Main_1_adj_2010\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__14326\,
            I => \c0.tx2.n2218_cascade_\
        );

    \I__1755\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14319\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__14322\,
            I => \N__14315\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__14319\,
            I => \N__14312\
        );

    \I__1752\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14309\
        );

    \I__1751\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14306\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__14312\,
            I => \N__14303\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__14309\,
            I => \c0.tx2.n3577\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__14306\,
            I => \c0.tx2.n3577\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__14303\,
            I => \c0.tx2.n3577\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__14296\,
            I => \N__14293\
        );

    \I__1745\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14290\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__14290\,
            I => \N__14287\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__14287\,
            I => \c0.n5953\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__14284\,
            I => \N__14281\
        );

    \I__1741\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14278\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__1739\ : Span4Mux_s2_h
    port map (
            O => \N__14275\,
            I => \N__14272\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__14272\,
            I => \c0.n5956\
        );

    \I__1737\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__14266\,
            I => n2392
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__14263\,
            I => \N__14245\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__14262\,
            I => \N__14242\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__14261\,
            I => \N__14229\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__14260\,
            I => \N__14226\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__14259\,
            I => \N__14223\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__14258\,
            I => \N__14220\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__14257\,
            I => \N__14217\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__14256\,
            I => \N__14214\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__14255\,
            I => \N__14211\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__14254\,
            I => \N__14208\
        );

    \I__1725\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14204\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__14252\,
            I => \N__14201\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__14251\,
            I => \N__14198\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__14250\,
            I => \N__14195\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__14249\,
            I => \N__14192\
        );

    \I__1720\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14181\
        );

    \I__1719\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14181\
        );

    \I__1718\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14181\
        );

    \I__1717\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14181\
        );

    \I__1716\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14181\
        );

    \I__1715\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14174\
        );

    \I__1714\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14174\
        );

    \I__1713\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14174\
        );

    \I__1712\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14169\
        );

    \I__1711\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14169\
        );

    \I__1710\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14162\
        );

    \I__1709\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14162\
        );

    \I__1708\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14162\
        );

    \I__1707\ : InMux
    port map (
            O => \N__14229\,
            I => \N__14153\
        );

    \I__1706\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14153\
        );

    \I__1705\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14153\
        );

    \I__1704\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14153\
        );

    \I__1703\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14144\
        );

    \I__1702\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14144\
        );

    \I__1701\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14144\
        );

    \I__1700\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14144\
        );

    \I__1699\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14141\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14138\
        );

    \I__1697\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14135\
        );

    \I__1696\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14128\
        );

    \I__1695\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14128\
        );

    \I__1694\ : InMux
    port map (
            O => \N__14192\,
            I => \N__14128\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__14181\,
            I => \N__14121\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__14174\,
            I => \N__14121\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__14169\,
            I => \N__14121\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__14162\,
            I => \N__14114\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__14153\,
            I => \N__14114\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__14144\,
            I => \N__14114\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__14141\,
            I => \r_SM_Main_2_adj_2009\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__14138\,
            I => \r_SM_Main_2_adj_2009\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__14135\,
            I => \r_SM_Main_2_adj_2009\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__14128\,
            I => \r_SM_Main_2_adj_2009\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__14121\,
            I => \r_SM_Main_2_adj_2009\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__14114\,
            I => \r_SM_Main_2_adj_2009\
        );

    \I__1681\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14098\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14093\
        );

    \I__1679\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14088\
        );

    \I__1678\ : InMux
    port map (
            O => \N__14096\,
            I => \N__14088\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__14093\,
            I => \N__14080\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__14088\,
            I => \N__14077\
        );

    \I__1675\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14068\
        );

    \I__1674\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14068\
        );

    \I__1673\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14068\
        );

    \I__1672\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14068\
        );

    \I__1671\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14065\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__14080\,
            I => n5037
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__14077\,
            I => n5037
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__14068\,
            I => n5037
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__14065\,
            I => n5037
        );

    \I__1666\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14051\
        );

    \I__1665\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14048\
        );

    \I__1664\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14045\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__14051\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__14048\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__14045\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1660\ : InMux
    port map (
            O => \N__14038\,
            I => \c0.n4400\
        );

    \I__1659\ : InMux
    port map (
            O => \N__14035\,
            I => \c0.n4401\
        );

    \I__1658\ : InMux
    port map (
            O => \N__14032\,
            I => \c0.n4402\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__14029\,
            I => \c0.tx.n12_cascade_\
        );

    \I__1656\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14019\
        );

    \I__1655\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14014\
        );

    \I__1654\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14014\
        );

    \I__1653\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14011\
        );

    \I__1652\ : InMux
    port map (
            O => \N__14022\,
            I => \N__14008\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__14019\,
            I => \r_Clock_Count_8\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__14014\,
            I => \r_Clock_Count_8\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__14011\,
            I => \r_Clock_Count_8\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__14008\,
            I => \r_Clock_Count_8\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__13999\,
            I => \n1307_cascade_\
        );

    \I__1646\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13992\
        );

    \I__1645\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__13992\,
            I => n3595
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__13989\,
            I => n3595
        );

    \I__1642\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13973\
        );

    \I__1641\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13968\
        );

    \I__1640\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13968\
        );

    \I__1639\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13963\
        );

    \I__1638\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13963\
        );

    \I__1637\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13954\
        );

    \I__1636\ : InMux
    port map (
            O => \N__13978\,
            I => \N__13954\
        );

    \I__1635\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13954\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13954\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__13973\,
            I => \N__13951\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__13968\,
            I => n4221
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__13963\,
            I => n4221
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__13954\,
            I => n4221
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__13951\,
            I => n4221
        );

    \I__1628\ : InMux
    port map (
            O => \N__13942\,
            I => \N__13939\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__13939\,
            I => n2
        );

    \I__1626\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13933\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__13933\,
            I => n1307
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__13930\,
            I => \n4_adj_2003_cascade_\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__13927\,
            I => \N__13923\
        );

    \I__1622\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13920\
        );

    \I__1621\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13917\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__13920\,
            I => n4155
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__13917\,
            I => n4155
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__13912\,
            I => \N__13909\
        );

    \I__1617\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13906\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__13906\,
            I => n2372
        );

    \I__1615\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13898\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13902\,
            I => \N__13895\
        );

    \I__1613\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13892\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__13898\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__13895\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__13892\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__13882\,
            I => n2395
        );

    \I__1607\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13874\
        );

    \I__1606\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13871\
        );

    \I__1605\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13868\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__13874\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13871\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__13868\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1601\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13857\
        );

    \I__1600\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13847\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__13857\,
            I => \N__13844\
        );

    \I__1598\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13841\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13838\
        );

    \I__1596\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13831\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13831\
        );

    \I__1594\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13831\
        );

    \I__1593\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13826\
        );

    \I__1592\ : InMux
    port map (
            O => \N__13850\,
            I => \N__13826\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__13847\,
            I => \N__13819\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__13844\,
            I => \N__13819\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__13841\,
            I => \N__13819\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13816\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__13831\,
            I => \r_SM_Main_0_adj_2011\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__13826\,
            I => \r_SM_Main_0_adj_2011\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__13819\,
            I => \r_SM_Main_0_adj_2011\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__13816\,
            I => \r_SM_Main_0_adj_2011\
        );

    \I__1583\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13796\
        );

    \I__1582\ : InMux
    port map (
            O => \N__13806\,
            I => \N__13796\
        );

    \I__1581\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13796\
        );

    \I__1580\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13790\
        );

    \I__1579\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13790\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__13796\,
            I => \N__13787\
        );

    \I__1577\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13784\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__13790\,
            I => \r_SM_Main_2_N_1767_1\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__13787\,
            I => \r_SM_Main_2_N_1767_1\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__13784\,
            I => \r_SM_Main_2_N_1767_1\
        );

    \I__1573\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13773\
        );

    \I__1572\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13770\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__13773\,
            I => \N__13765\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__13770\,
            I => \N__13765\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__13765\,
            I => data_out_19_4
        );

    \I__1568\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13756\
        );

    \I__1567\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13756\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__13756\,
            I => data_out_18_4
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__13753\,
            I => \c0.n17_cascade_\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__13750\,
            I => \tx_data_4_N_keep_cascade_\
        );

    \I__1563\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13744\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13741\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__13741\,
            I => n8_adj_2001
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__13738\,
            I => \c0.tx.r_SM_Main_2_N_1767_1_cascade_\
        );

    \I__1559\ : InMux
    port map (
            O => \N__13735\,
            I => \N__13732\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__13732\,
            I => n5041
        );

    \I__1557\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13726\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__13726\,
            I => \N__13720\
        );

    \I__1555\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13717\
        );

    \I__1554\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13714\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__13723\,
            I => \N__13711\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__13720\,
            I => \N__13703\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__13717\,
            I => \N__13703\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__13714\,
            I => \N__13703\
        );

    \I__1549\ : InMux
    port map (
            O => \N__13711\,
            I => \N__13697\
        );

    \I__1548\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13697\
        );

    \I__1547\ : Span4Mux_v
    port map (
            O => \N__13703\,
            I => \N__13694\
        );

    \I__1546\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13691\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__13697\,
            I => \c0.tx_transmit\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__13694\,
            I => \c0.tx_transmit\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__13691\,
            I => \c0.tx_transmit\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__13684\,
            I => \n4316_cascade_\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__13681\,
            I => \N__13678\
        );

    \I__1540\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13675\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__13675\,
            I => n7_adj_2002
        );

    \I__1538\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13668\
        );

    \I__1537\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13665\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__13668\,
            I => \N__13662\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__13665\,
            I => n5066
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__13662\,
            I => n5066
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__13657\,
            I => \N__13651\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13646\
        );

    \I__1531\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13646\
        );

    \I__1530\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13643\
        );

    \I__1529\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13638\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13635\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__13643\,
            I => \N__13632\
        );

    \I__1526\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13627\
        );

    \I__1525\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13627\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13638\,
            I => tx_active
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__13635\,
            I => tx_active
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__13632\,
            I => tx_active
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__13627\,
            I => tx_active
        );

    \I__1520\ : InMux
    port map (
            O => \N__13618\,
            I => \N__13614\
        );

    \I__1519\ : InMux
    port map (
            O => \N__13617\,
            I => \N__13611\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__13614\,
            I => \c0.tx_transmit_N_568_5\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__13611\,
            I => \c0.tx_transmit_N_568_5\
        );

    \I__1516\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13602\
        );

    \I__1515\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13599\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__13602\,
            I => \c0.tx_transmit_N_568_6\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__13599\,
            I => \c0.tx_transmit_N_568_6\
        );

    \I__1512\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13590\
        );

    \I__1511\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13587\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__13590\,
            I => \c0.tx_transmit_N_568_7\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__13587\,
            I => \c0.tx_transmit_N_568_7\
        );

    \I__1508\ : InMux
    port map (
            O => \N__13582\,
            I => \N__13576\
        );

    \I__1507\ : InMux
    port map (
            O => \N__13581\,
            I => \N__13571\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13571\
        );

    \I__1505\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13568\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__13576\,
            I => \c0.tx_transmit_N_568_4\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__13571\,
            I => \c0.tx_transmit_N_568_4\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__13568\,
            I => \c0.tx_transmit_N_568_4\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13557\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13554\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__13557\,
            I => \c0.n103\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__13554\,
            I => \c0.n103\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13546\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__13546\,
            I => \c0.n109\
        );

    \I__1495\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13534\
        );

    \I__1494\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13534\
        );

    \I__1493\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13529\
        );

    \I__1492\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13529\
        );

    \I__1491\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13526\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__13534\,
            I => \c0.n45\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__13529\,
            I => \c0.n45\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__13526\,
            I => \c0.n45\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__13519\,
            I => \c0.n109_cascade_\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__13516\,
            I => \n4315_cascade_\
        );

    \I__1485\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13506\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__13509\,
            I => \N__13503\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__13506\,
            I => \N__13500\
        );

    \I__1481\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13497\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__13500\,
            I => \c0.rx.n3573\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__13497\,
            I => \c0.rx.n3573\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__13492\,
            I => \c0.rx.n3573_cascade_\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__13489\,
            I => \c0.n20_adj_1918_cascade_\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__13486\,
            I => \N__13482\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__13485\,
            I => \N__13479\
        );

    \I__1474\ : InMux
    port map (
            O => \N__13482\,
            I => \N__13465\
        );

    \I__1473\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13465\
        );

    \I__1472\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13465\
        );

    \I__1471\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13465\
        );

    \I__1470\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13465\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__13465\,
            I => \c0.n87\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__13462\,
            I => \c0.n87_cascade_\
        );

    \I__1467\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13456\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__13456\,
            I => \c0.n16_adj_1909\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__13453\,
            I => \c0.rx.n4_adj_1866_cascade_\
        );

    \I__1464\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13441\
        );

    \I__1463\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13441\
        );

    \I__1462\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13441\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__13441\,
            I => \N__13436\
        );

    \I__1460\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13431\
        );

    \I__1459\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13431\
        );

    \I__1458\ : Span4Mux_s1_h
    port map (
            O => \N__13436\,
            I => \N__13428\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__13431\,
            I => \c0.rx.n4011\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__13428\,
            I => \c0.rx.n4011\
        );

    \I__1455\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13419\
        );

    \I__1454\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13416\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13411\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__13416\,
            I => \N__13411\
        );

    \I__1451\ : Span4Mux_v
    port map (
            O => \N__13411\,
            I => \N__13407\
        );

    \I__1450\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13404\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__13407\,
            I => data_in_5_1
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__13404\,
            I => data_in_5_1
        );

    \I__1447\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13393\
        );

    \I__1446\ : InMux
    port map (
            O => \N__13398\,
            I => \N__13390\
        );

    \I__1445\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13387\
        );

    \I__1444\ : InMux
    port map (
            O => \N__13396\,
            I => \N__13384\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__13393\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__13390\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__13387\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__13384\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1439\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13369\
        );

    \I__1438\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13366\
        );

    \I__1437\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13363\
        );

    \I__1436\ : InMux
    port map (
            O => \N__13372\,
            I => \N__13360\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__13369\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__13366\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__13363\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__13360\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__1431\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13348\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__13348\,
            I => \c0.rx.n37\
        );

    \I__1429\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13341\
        );

    \I__1428\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13335\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__13341\,
            I => \N__13332\
        );

    \I__1426\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13329\
        );

    \I__1425\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13326\
        );

    \I__1424\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13323\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__13335\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__13332\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__13329\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__13326\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__13323\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__13312\,
            I => \c0.rx.n37_cascade_\
        );

    \I__1417\ : InMux
    port map (
            O => \N__13309\,
            I => \N__13302\
        );

    \I__1416\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13299\
        );

    \I__1415\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13296\
        );

    \I__1414\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13291\
        );

    \I__1413\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13291\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__13302\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__13299\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__13296\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__13291\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1408\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13275\
        );

    \I__1407\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13272\
        );

    \I__1406\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13265\
        );

    \I__1405\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13265\
        );

    \I__1404\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13265\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__13275\,
            I => \r_SM_Main_2_N_1830_0\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__13272\,
            I => \r_SM_Main_2_N_1830_0\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__13265\,
            I => \r_SM_Main_2_N_1830_0\
        );

    \I__1400\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13255\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__13255\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__13252\,
            I => \n12_adj_1995_cascade_\
        );

    \I__1397\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13246\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__13246\,
            I => n5316
        );

    \I__1395\ : InMux
    port map (
            O => \N__13243\,
            I => \N__13233\
        );

    \I__1394\ : InMux
    port map (
            O => \N__13242\,
            I => \N__13233\
        );

    \I__1393\ : InMux
    port map (
            O => \N__13241\,
            I => \N__13226\
        );

    \I__1392\ : InMux
    port map (
            O => \N__13240\,
            I => \N__13226\
        );

    \I__1391\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13226\
        );

    \I__1390\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13219\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__13233\,
            I => \N__13216\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N__13213\
        );

    \I__1387\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13206\
        );

    \I__1386\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13206\
        );

    \I__1385\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13206\
        );

    \I__1384\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13203\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__13219\,
            I => n16_adj_1993
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__13216\,
            I => n16_adj_1993
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__13213\,
            I => n16_adj_1993
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__13206\,
            I => n16_adj_1993
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__13203\,
            I => n16_adj_1993
        );

    \I__1378\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13189\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__13189\,
            I => n5491
        );

    \I__1376\ : InMux
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__13183\,
            I => \c0.rx.n5535\
        );

    \I__1374\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13177\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__13177\,
            I => \c0.rx.n2157\
        );

    \I__1372\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13171\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__13171\,
            I => \c0.rx.n5538\
        );

    \I__1370\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13165\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__13165\,
            I => \c0.rx.n5539\
        );

    \I__1368\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13159\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__13159\,
            I => \c0.rx.n40\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__13156\,
            I => \c0.rx.r_SM_Main_2_N_1824_2_cascade_\
        );

    \I__1365\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13150\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__13150\,
            I => n4474
        );

    \I__1363\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13144\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__13144\,
            I => n2156
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__13141\,
            I => \n4474_cascade_\
        );

    \I__1360\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13134\
        );

    \I__1359\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13131\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__13134\,
            I => \N__13128\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__13131\,
            I => \c0.data_in_frame_18_1\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__13128\,
            I => \c0.data_in_frame_18_1\
        );

    \I__1355\ : InMux
    port map (
            O => \N__13123\,
            I => \N__13120\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__13120\,
            I => \N__13117\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__13117\,
            I => \c0.n5369\
        );

    \I__1352\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13111\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13108\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__13108\,
            I => \c0.n5869\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__13105\,
            I => \N__13102\
        );

    \I__1348\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13099\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__13099\,
            I => \c0.n5959\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__13096\,
            I => \N__13093\
        );

    \I__1345\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13090\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__13090\,
            I => \N__13087\
        );

    \I__1343\ : Odrv12
    port map (
            O => \N__13087\,
            I => \c0.n5962\
        );

    \I__1342\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13080\
        );

    \I__1341\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13077\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__13080\,
            I => \N__13074\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__13077\,
            I => \c0.data_in_frame_18_3\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__13074\,
            I => \c0.data_in_frame_18_3\
        );

    \I__1337\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13066\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__13066\,
            I => n5051
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__13063\,
            I => \c0.n5725_cascade_\
        );

    \I__1334\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13049\
        );

    \I__1333\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13049\
        );

    \I__1332\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13049\
        );

    \I__1331\ : InMux
    port map (
            O => \N__13057\,
            I => \N__13042\
        );

    \I__1330\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13039\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__13049\,
            I => \N__13036\
        );

    \I__1328\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13029\
        );

    \I__1327\ : InMux
    port map (
            O => \N__13047\,
            I => \N__13029\
        );

    \I__1326\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13029\
        );

    \I__1325\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13026\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__13042\,
            I => \N__13021\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__13039\,
            I => \N__13021\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__13036\,
            I => \c0.n1058\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__13029\,
            I => \c0.n1058\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__13026\,
            I => \c0.n1058\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__13021\,
            I => \c0.n1058\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__13012\,
            I => \c0.n5728_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__13009\,
            I => \N__13006\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__13006\,
            I => \c0.n5974\
        );

    \I__1315\ : InMux
    port map (
            O => \N__13003\,
            I => \N__13000\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__13000\,
            I => \N__12997\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__12997\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__1312\ : CEMux
    port map (
            O => \N__12994\,
            I => \N__12989\
        );

    \I__1311\ : CEMux
    port map (
            O => \N__12993\,
            I => \N__12986\
        );

    \I__1310\ : CEMux
    port map (
            O => \N__12992\,
            I => \N__12983\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__12989\,
            I => \N__12977\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12986\,
            I => \N__12977\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__12983\,
            I => \N__12974\
        );

    \I__1306\ : CEMux
    port map (
            O => \N__12982\,
            I => \N__12971\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__12977\,
            I => \N__12968\
        );

    \I__1304\ : Span4Mux_s1_h
    port map (
            O => \N__12974\,
            I => \N__12963\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__12971\,
            I => \N__12963\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__12968\,
            I => \c0.tx2.n1592\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__12963\,
            I => \c0.tx2.n1592\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__12958\,
            I => \c0.n5803_cascade_\
        );

    \I__1299\ : InMux
    port map (
            O => \N__12955\,
            I => \N__12952\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__12952\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__12949\,
            I => \c0.n5665_cascade_\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__12946\,
            I => \c0.n5372_cascade_\
        );

    \I__1295\ : InMux
    port map (
            O => \N__12943\,
            I => \N__12940\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__12940\,
            I => \c0.n5659\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__12937\,
            I => \N__12934\
        );

    \I__1292\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12931\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__12931\,
            I => \c0.n5938\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__12928\,
            I => \c0.n5971_cascade_\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__12925\,
            I => \N__12922\
        );

    \I__1288\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12919\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__12919\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__1286\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12913\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__12913\,
            I => \c0.tx2.n5947\
        );

    \I__1284\ : InMux
    port map (
            O => \N__12910\,
            I => \N__12907\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__12907\,
            I => \c0.tx2.n5950\
        );

    \I__1282\ : InMux
    port map (
            O => \N__12904\,
            I => \N__12901\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__12901\,
            I => n1345
        );

    \I__1280\ : InMux
    port map (
            O => \N__12898\,
            I => \N__12895\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__12895\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__1278\ : InMux
    port map (
            O => \N__12892\,
            I => \N__12889\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__12889\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__12886\,
            I => \N__12881\
        );

    \I__1275\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12878\
        );

    \I__1274\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12875\
        );

    \I__1273\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12872\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__12878\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__12875\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__12872\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1269\ : InMux
    port map (
            O => \N__12865\,
            I => \N__12862\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__12862\,
            I => n2399
        );

    \I__1267\ : InMux
    port map (
            O => \N__12859\,
            I => \c0.tx2.n4429\
        );

    \I__1266\ : InMux
    port map (
            O => \N__12856\,
            I => \c0.tx2.n4430\
        );

    \I__1265\ : InMux
    port map (
            O => \N__12853\,
            I => \c0.tx2.n4431\
        );

    \I__1264\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12845\
        );

    \I__1263\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12842\
        );

    \I__1262\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12839\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__12845\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__12842\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__12839\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1258\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12829\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__12829\,
            I => \N__12826\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__12826\,
            I => n2382
        );

    \I__1255\ : InMux
    port map (
            O => \N__12823\,
            I => \c0.tx2.n4432\
        );

    \I__1254\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12815\
        );

    \I__1253\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12812\
        );

    \I__1252\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12809\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__12815\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__12812\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__12809\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1248\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12799\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__12799\,
            I => \N__12796\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__12796\,
            I => n2379
        );

    \I__1245\ : InMux
    port map (
            O => \N__12793\,
            I => \c0.tx2.n4433\
        );

    \I__1244\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12785\
        );

    \I__1243\ : InMux
    port map (
            O => \N__12789\,
            I => \N__12782\
        );

    \I__1242\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12779\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__12785\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__12782\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__12779\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1238\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12769\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__12769\,
            I => \N__12766\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__12766\,
            I => n2376
        );

    \I__1235\ : InMux
    port map (
            O => \N__12763\,
            I => \c0.tx2.n4434\
        );

    \I__1234\ : InMux
    port map (
            O => \N__12760\,
            I => \c0.tx2.n4435\
        );

    \I__1233\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12752\
        );

    \I__1232\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12749\
        );

    \I__1231\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12745\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__12752\,
            I => \N__12740\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__12749\,
            I => \N__12740\
        );

    \I__1228\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12737\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__12745\,
            I => \r_Clock_Count_8_adj_2012\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__12740\,
            I => \r_Clock_Count_8_adj_2012\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__12737\,
            I => \r_Clock_Count_8_adj_2012\
        );

    \I__1224\ : InMux
    port map (
            O => \N__12730\,
            I => \bfn_2_24_0_\
        );

    \I__1223\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12724\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__12724\,
            I => \N__12721\
        );

    \I__1221\ : Odrv4
    port map (
            O => \N__12721\,
            I => n2369
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__12718\,
            I => \c0.tx2.n5_cascade_\
        );

    \I__1219\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12712\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__12712\,
            I => \c0.tx2.n3591\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__12709\,
            I => \c0.tx2.n3591_cascade_\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__12706\,
            I => \r_SM_Main_2_N_1767_1_cascade_\
        );

    \I__1215\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12699\
        );

    \I__1214\ : InMux
    port map (
            O => \N__12702\,
            I => \N__12696\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__12699\,
            I => \N__12691\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__12696\,
            I => \N__12691\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__12691\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__12688\,
            I => \N__12685\
        );

    \I__1209\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12682\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12682\,
            I => n2460
        );

    \I__1207\ : InMux
    port map (
            O => \N__12679\,
            I => \bfn_2_23_0_\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__12676\,
            I => \N__12673\
        );

    \I__1205\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12669\
        );

    \I__1204\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12666\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__12669\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__12666\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__1201\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12658\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__12658\,
            I => \c0.tx.n313\
        );

    \I__1199\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12652\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__12652\,
            I => n316
        );

    \I__1197\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12646\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__12646\,
            I => n314
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__12643\,
            I => \N__12640\
        );

    \I__1194\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12637\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__12637\,
            I => n317
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__12634\,
            I => \N__12631\
        );

    \I__1191\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12626\
        );

    \I__1190\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12623\
        );

    \I__1189\ : InMux
    port map (
            O => \N__12629\,
            I => \N__12620\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__12626\,
            I => \r_Clock_Count_2\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__12623\,
            I => \r_Clock_Count_2\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__12620\,
            I => \r_Clock_Count_2\
        );

    \I__1185\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12608\
        );

    \I__1184\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12605\
        );

    \I__1183\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12602\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__12608\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__12605\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__12602\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__12595\,
            I => \N__12591\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__12594\,
            I => \N__12587\
        );

    \I__1177\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12584\
        );

    \I__1176\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12581\
        );

    \I__1175\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12578\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__12584\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__12581\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__12578\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__1171\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12566\
        );

    \I__1170\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12561\
        );

    \I__1169\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12561\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__12566\,
            I => \r_Clock_Count_5\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__12561\,
            I => \r_Clock_Count_5\
        );

    \I__1166\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12551\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12555\,
            I => \N__12546\
        );

    \I__1164\ : InMux
    port map (
            O => \N__12554\,
            I => \N__12546\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__12551\,
            I => \r_Clock_Count_4\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__12546\,
            I => \r_Clock_Count_4\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__12541\,
            I => \c0.tx.n5_cascade_\
        );

    \I__1160\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12533\
        );

    \I__1159\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12528\
        );

    \I__1158\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12528\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__12533\,
            I => \r_Clock_Count_7\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__12528\,
            I => \r_Clock_Count_7\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__12523\,
            I => \n3595_cascade_\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__12520\,
            I => \N__12517\
        );

    \I__1153\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12514\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__12514\,
            I => \c0.tx.n5520\
        );

    \I__1151\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12506\
        );

    \I__1150\ : InMux
    port map (
            O => \N__12510\,
            I => \N__12501\
        );

    \I__1149\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12501\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__12506\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__12501\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__1146\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12493\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__12493\,
            I => n1760
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__12490\,
            I => \c0.n1529_cascade_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12484\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__12484\,
            I => \c0.n1801\
        );

    \I__1141\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12478\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__12478\,
            I => \c0.tx.n315\
        );

    \I__1139\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12472\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__12472\,
            I => n319
        );

    \I__1137\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12466\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__12466\,
            I => \c0.tx.n320\
        );

    \I__1135\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12460\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__12460\,
            I => \c0.tx.n321\
        );

    \I__1133\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12454\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__12454\,
            I => \c0.n50\
        );

    \I__1131\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12448\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__12448\,
            I => \c0.tx_active_prev\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__12445\,
            I => \c0.n5540_cascade_\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__12442\,
            I => \c0.n5977_cascade_\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__12439\,
            I => \n1760_cascade_\
        );

    \I__1126\ : InMux
    port map (
            O => \N__12436\,
            I => \c0.n4378\
        );

    \I__1125\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12427\
        );

    \I__1124\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12427\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__12427\,
            I => \c0.tx_transmit_N_568_2\
        );

    \I__1122\ : InMux
    port map (
            O => \N__12424\,
            I => \c0.n4379\
        );

    \I__1121\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12415\
        );

    \I__1120\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12415\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__12415\,
            I => \c0.tx_transmit_N_568_3\
        );

    \I__1118\ : InMux
    port map (
            O => \N__12412\,
            I => \c0.n4380\
        );

    \I__1117\ : InMux
    port map (
            O => \N__12409\,
            I => \c0.n4381\
        );

    \I__1116\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12403\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__12403\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__1114\ : InMux
    port map (
            O => \N__12400\,
            I => \c0.n4382\
        );

    \I__1113\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12394\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__12394\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__1111\ : InMux
    port map (
            O => \N__12391\,
            I => \c0.n4383\
        );

    \I__1110\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12385\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__12385\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__1108\ : InMux
    port map (
            O => \N__12382\,
            I => \c0.n4384\
        );

    \I__1107\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12376\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__12376\,
            I => n5490
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__12373\,
            I => \c0.rx.n3980_cascade_\
        );

    \I__1104\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12367\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__12367\,
            I => \c0.rx.n5532\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__12364\,
            I => \c0.rx.n5298_cascade_\
        );

    \I__1101\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12358\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__12358\,
            I => \c0.rx.n5536\
        );

    \I__1099\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12349\
        );

    \I__1098\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12349\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__12349\,
            I => \c0.rx.n5049\
        );

    \I__1096\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12343\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__12343\,
            I => n5050
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__12340\,
            I => \c0.rx.n5923_cascade_\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__12337\,
            I => \c0.rx.n5926_cascade_\
        );

    \I__1092\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12331\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__12331\,
            I => \N__12328\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__12328\,
            I => \c0.rx.n5537\
        );

    \I__1089\ : InMux
    port map (
            O => \N__12325\,
            I => \c0.rx.n4422\
        );

    \I__1088\ : InMux
    port map (
            O => \N__12322\,
            I => \c0.rx.n4423\
        );

    \I__1087\ : InMux
    port map (
            O => \N__12319\,
            I => \c0.rx.n4424\
        );

    \I__1086\ : InMux
    port map (
            O => \N__12316\,
            I => \c0.rx.n4425\
        );

    \I__1085\ : InMux
    port map (
            O => \N__12313\,
            I => \c0.rx.n4426\
        );

    \I__1084\ : InMux
    port map (
            O => \N__12310\,
            I => \c0.rx.n4427\
        );

    \I__1083\ : InMux
    port map (
            O => \N__12307\,
            I => \c0.rx.n4428\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__12304\,
            I => \n2156_cascade_\
        );

    \I__1081\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12298\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__12298\,
            I => n8
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__12295\,
            I => \N__12292\
        );

    \I__1078\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12288\
        );

    \I__1077\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12285\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__12288\,
            I => \N__12282\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__12285\,
            I => \c0.data_in_frame_19_0\
        );

    \I__1074\ : Odrv12
    port map (
            O => \N__12282\,
            I => \c0.data_in_frame_19_0\
        );

    \I__1073\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12272\
        );

    \I__1072\ : IoInMux
    port map (
            O => \N__12276\,
            I => \N__12269\
        );

    \I__1071\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12266\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__12269\,
            I => tx2_o
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__12266\,
            I => tx2_o
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__12263\,
            I => tx2_o
        );

    \I__1066\ : IoInMux
    port map (
            O => \N__12256\,
            I => \N__12253\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__12253\,
            I => tx2_enable
        );

    \I__1064\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12247\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__12247\,
            I => \c0.n5402\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__12244\,
            I => \N__12240\
        );

    \I__1061\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12237\
        );

    \I__1060\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12234\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__12237\,
            I => \c0.data_in_frame_19_3\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__12234\,
            I => \c0.data_in_frame_19_3\
        );

    \I__1057\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12226\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__12226\,
            I => \c0.n5863\
        );

    \I__1055\ : InMux
    port map (
            O => \N__12223\,
            I => \bfn_1_30_0_\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__12220\,
            I => \c0.n5920_cascade_\
        );

    \I__1053\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12214\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__12214\,
            I => \c0.n5662\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__12211\,
            I => \N__12208\
        );

    \I__1050\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12205\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__12205\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__1048\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12199\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__12199\,
            I => \c0.tx2.n5929\
        );

    \I__1046\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12193\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__12193\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__1044\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12187\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12184\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__12184\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__12181\,
            I => \c0.n5399_cascade_\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__12178\,
            I => \c0.n5857_cascade_\
        );

    \I__1039\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12172\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__12172\,
            I => \c0.n5860\
        );

    \I__1037\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12166\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__12166\,
            I => \N__12163\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__12163\,
            I => \c0.tx2.o_Tx_Serial_N_1798\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__12160\,
            I => \n3_cascade_\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__12157\,
            I => \c0.tx2.n5312_cascade_\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__12154\,
            I => \c0.n5815_cascade_\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__12151\,
            I => \N__12148\
        );

    \I__1030\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12145\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__12145\,
            I => \c0.n5818\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__12142\,
            I => \c0.tx2.n5932_cascade_\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__12139\,
            I => \c0.n5917_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__12136\,
            I => \c0.tx.n4420\
        );

    \I__1025\ : InMux
    port map (
            O => \N__12133\,
            I => \bfn_1_22_0_\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__12130\,
            I => \n5037_cascade_\
        );

    \I__1023\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12124\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__12124\,
            I => n3611
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__12121\,
            I => \n4_adj_2008_cascade_\
        );

    \I__1020\ : InMux
    port map (
            O => \N__12118\,
            I => \bfn_1_21_0_\
        );

    \I__1019\ : InMux
    port map (
            O => \N__12115\,
            I => \c0.tx.n4414\
        );

    \I__1018\ : InMux
    port map (
            O => \N__12112\,
            I => \c0.tx.n4415\
        );

    \I__1017\ : InMux
    port map (
            O => \N__12109\,
            I => \c0.tx.n4416\
        );

    \I__1016\ : InMux
    port map (
            O => \N__12106\,
            I => \c0.tx.n4417\
        );

    \I__1015\ : InMux
    port map (
            O => \N__12103\,
            I => \c0.tx.n4418\
        );

    \I__1014\ : InMux
    port map (
            O => \N__12100\,
            I => \c0.tx.n4419\
        );

    \I__1013\ : IoInMux
    port map (
            O => \N__12097\,
            I => \N__12094\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__12094\,
            I => \N__12091\
        );

    \I__1011\ : IoSpan4Mux
    port map (
            O => \N__12091\,
            I => \N__12088\
        );

    \I__1010\ : IoSpan4Mux
    port map (
            O => \N__12088\,
            I => \N__12085\
        );

    \I__1009\ : IoSpan4Mux
    port map (
            O => \N__12085\,
            I => \N__12082\
        );

    \I__1008\ : Odrv4
    port map (
            O => \N__12082\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n4436\,
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n4421\,
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n4411\,
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_6_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_17_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n4392\,
            carryinitout => \bfn_6_18_0_\
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4444,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4452,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4460,
            carryinitout => \bfn_15_28_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12097\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_937_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18977\,
            in1 => \N__20475\,
            in2 => \_gnd_net_\,
            in3 => \N__18754\,
            lcout => n5066,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16810\,
            in1 => \N__18978\,
            in2 => \N__20476\,
            in3 => \N__21076\,
            lcout => n7_adj_1998,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12672\,
            in2 => \_gnd_net_\,
            in3 => \N__12118\,
            lcout => \c0.tx.n321\,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => \c0.tx.n4414\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12590\,
            in2 => \_gnd_net_\,
            in3 => \N__12115\,
            lcout => \c0.tx.n320\,
            ltout => OPEN,
            carryin => \c0.tx.n4414\,
            carryout => \c0.tx.n4415\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12630\,
            in2 => \_gnd_net_\,
            in3 => \N__12112\,
            lcout => n319,
            ltout => OPEN,
            carryin => \c0.tx.n4415\,
            carryout => \c0.tx.n4416\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__13984\,
            in1 => \N__12511\,
            in2 => \_gnd_net_\,
            in3 => \N__12109\,
            lcout => \c0.tx.n5520\,
            ltout => OPEN,
            carryin => \c0.tx.n4416\,
            carryout => \c0.tx.n4417\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12556\,
            in2 => \_gnd_net_\,
            in3 => \N__12106\,
            lcout => n317,
            ltout => OPEN,
            carryin => \c0.tx.n4417\,
            carryout => \c0.tx.n4418\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12571\,
            in2 => \_gnd_net_\,
            in3 => \N__12103\,
            lcout => n316,
            ltout => OPEN,
            carryin => \c0.tx.n4418\,
            carryout => \c0.tx.n4419\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12612\,
            in2 => \_gnd_net_\,
            in3 => \N__12100\,
            lcout => \c0.tx.n315\,
            ltout => OPEN,
            carryin => \c0.tx.n4419\,
            carryout => \c0.tx.n4420\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12538\,
            in2 => \_gnd_net_\,
            in3 => \N__12136\,
            lcout => n314,
            ltout => OPEN,
            carryin => \c0.tx.n4420\,
            carryout => \c0.tx.n4421\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14026\,
            in2 => \_gnd_net_\,
            in3 => \N__12133\,
            lcout => \c0.tx.n313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_1010_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__13856\,
            in1 => \N__12755\,
            in2 => \N__14390\,
            in3 => \N__12127\,
            lcout => n5037,
            ltout => \n5037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i8_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12727\,
            in2 => \N__12130\,
            in3 => \N__14236\,
            lcout => \r_Clock_Count_8_adj_2012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i3366_2_lut_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14235\,
            in2 => \_gnd_net_\,
            in3 => \N__12715\,
            lcout => n3611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15537\,
            in1 => \N__15598\,
            in2 => \_gnd_net_\,
            in3 => \N__15631\,
            lcout => \c0.tx2.n3577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5286_3_lut_4_lut_4_lut_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__13851\,
            in1 => \N__14385\,
            in2 => \N__15793\,
            in3 => \N__13803\,
            lcout => OPEN,
            ltout => \n4_adj_2008_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__14387\,
            in1 => \N__15749\,
            in2 => \N__12121\,
            in3 => \N__14239\,
            lcout => tx2_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__14238\,
            in1 => \_gnd_net_\,
            in2 => \N__12688\,
            in3 => \N__14083\,
            lcout => \c0.tx2.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4968_3_lut_4_lut_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__13804\,
            in1 => \N__13850\,
            in2 => \N__14397\,
            in3 => \N__14237\,
            lcout => OPEN,
            ltout => \c0.tx2.n5312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100100"
        )
    port map (
            in0 => \N__15632\,
            in1 => \N__14386\,
            in2 => \N__12157\,
            in3 => \N__14318\,
            lcout => \c0.tx2.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14525\,
            in1 => \N__13045\,
            in2 => \N__12151\,
            in3 => \N__21532\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35295\,
            ce => \N__12982\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5450_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__32524\,
            in1 => \N__16015\,
            in2 => \N__12295\,
            in3 => \N__33221\,
            lcout => OPEN,
            ltout => \c0.n5815_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5815_bdd_4_lut_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__29539\,
            in1 => \N__32525\,
            in2 => \N__12154\,
            in3 => \N__32026\,
            lcout => \c0.n5818\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5659_bdd_4_lut_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22060\,
            in1 => \N__34807\,
            in2 => \N__14443\,
            in3 => \N__12943\,
            lcout => \c0.n5662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n5929_bdd_4_lut_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__12190\,
            in1 => \N__12898\,
            in2 => \N__15604\,
            in3 => \N__12202\,
            lcout => OPEN,
            ltout => \c0.tx2.n5932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i341524_i1_3_lut_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15538\,
            in2 => \N__12142\,
            in3 => \N__12910\,
            lcout => \c0.tx2.o_Tx_Serial_N_1798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5543_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__14665\,
            in1 => \N__32522\,
            in2 => \N__14431\,
            in3 => \N__33222\,
            lcout => OPEN,
            ltout => \c0.n5917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5917_bdd_4_lut_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32523\,
            in1 => \N__22627\,
            in2 => \N__12139\,
            in3 => \N__25677\,
            lcout => OPEN,
            ltout => \c0.n5920_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14532\,
            in1 => \N__13060\,
            in2 => \N__12220\,
            in3 => \N__12217\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => \N__12992\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_5553_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__12196\,
            in1 => \N__15603\,
            in2 => \N__12211\,
            in3 => \N__15633\,
            lcout => \c0.tx2.n5929\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__34696\,
            in2 => \N__12937\,
            in3 => \N__13059\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => \N__12992\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14530\,
            in1 => \N__13058\,
            in2 => \N__14572\,
            in3 => \N__12175\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => \N__12992\,
            sr => \_gnd_net_\
        );

    \c0.n5869_bdd_4_lut_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__13114\,
            in1 => \N__25459\,
            in2 => \N__32588\,
            in3 => \N__21631\,
            lcout => OPEN,
            ltout => \c0.n5399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5505_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__34821\,
            in1 => \N__32115\,
            in2 => \N__12181\,
            in3 => \N__12250\,
            lcout => OPEN,
            ltout => \c0.n5857_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5857_bdd_4_lut_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__34806\,
            in1 => \N__25219\,
            in2 => \N__12178\,
            in3 => \N__21682\,
            lcout => \c0.n5860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110011001"
        )
    port map (
            in0 => \N__14398\,
            in1 => \N__13861\,
            in2 => \_gnd_net_\,
            in3 => \N__12169\,
            lcout => OPEN,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__14253\,
            in1 => \_gnd_net_\,
            in2 => \N__12160\,
            in3 => \N__12277\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i153_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__36175\,
            in1 => \N__12291\,
            in2 => \N__37268\,
            in3 => \N__21462\,
            lcout => \c0.data_in_frame_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12275\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5863_bdd_4_lut_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__12229\,
            in1 => \N__17566\,
            in2 => \N__15967\,
            in3 => \N__32518\,
            lcout => \c0.n5402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i34_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29324\,
            in1 => \N__13422\,
            in2 => \_gnd_net_\,
            in3 => \N__34147\,
            lcout => data_in_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i156_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__12243\,
            in1 => \N__15857\,
            in2 => \N__37228\,
            in3 => \N__36289\,
            lcout => \c0.data_in_frame_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5568_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__13084\,
            in1 => \N__32586\,
            in2 => \N__12244\,
            in3 => \N__33273\,
            lcout => \c0.n5959\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5490_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33272\,
            in1 => \N__23068\,
            in2 => \N__32629\,
            in3 => \N__28809\,
            lcout => \c0.n5863\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010000110000"
        )
    port map (
            in0 => \N__13513\,
            in1 => \N__13180\,
            in2 => \N__18177\,
            in3 => \N__18283\,
            lcout => \c0.rx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__12301\,
            in1 => \N__14911\,
            in2 => \_gnd_net_\,
            in3 => \N__12223\,
            lcout => n5491,
            ltout => OPEN,
            carryin => \bfn_1_30_0_\,
            carryout => \c0.rx.n4422\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__13448\,
            in1 => \N__13345\,
            in2 => \_gnd_net_\,
            in3 => \N__12325\,
            lcout => \c0.rx.n5537\,
            ltout => OPEN,
            carryin => \c0.rx.n4422\,
            carryout => \c0.rx.n4423\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__13440\,
            in1 => \N__14730\,
            in2 => \_gnd_net_\,
            in3 => \N__12322\,
            lcout => \c0.rx.n5536\,
            ltout => OPEN,
            carryin => \c0.rx.n4423\,
            carryout => \c0.rx.n4424\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__13449\,
            in1 => \N__13308\,
            in2 => \_gnd_net_\,
            in3 => \N__12319\,
            lcout => \c0.rx.n5539\,
            ltout => OPEN,
            carryin => \c0.rx.n4424\,
            carryout => \c0.rx.n4425\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__13439\,
            in1 => \N__13374\,
            in2 => \_gnd_net_\,
            in3 => \N__12316\,
            lcout => \c0.rx.n5535\,
            ltout => OPEN,
            carryin => \c0.rx.n4425\,
            carryout => \c0.rx.n4426\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__13450\,
            in1 => \N__13398\,
            in2 => \_gnd_net_\,
            in3 => \N__12313\,
            lcout => \c0.rx.n5538\,
            ltout => OPEN,
            carryin => \c0.rx.n4426\,
            carryout => \c0.rx.n4427\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__12355\,
            in1 => \N__14881\,
            in2 => \_gnd_net_\,
            in3 => \N__12310\,
            lcout => n5051,
            ltout => OPEN,
            carryin => \c0.rx.n4427\,
            carryout => \c0.rx.n4428\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12354\,
            in2 => \N__14767\,
            in3 => \N__12307\,
            lcout => n5050,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i59_3_lut_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__14724\,
            in1 => \N__13338\,
            in2 => \_gnd_net_\,
            in3 => \N__13305\,
            lcout => \c0.rx.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_791_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__18109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18269\,
            lcout => n2156,
            ltout => \n2156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4941_1_lut_4_lut_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111111"
        )
    port map (
            in0 => \N__18330\,
            in1 => \N__13282\,
            in2 => \N__12304\,
            in3 => \N__13153\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4954_2_lut_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14760\,
            in2 => \_gnd_net_\,
            in3 => \N__13397\,
            lcout => OPEN,
            ltout => \c0.rx.n5298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4972_4_lut_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13339\,
            in1 => \N__13306\,
            in2 => \N__12364\,
            in3 => \N__13373\,
            lcout => n5316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13224\,
            in1 => \N__14725\,
            in2 => \_gnd_net_\,
            in3 => \N__12361\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_4_lut_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__12379\,
            in1 => \N__18046\,
            in2 => \N__18282\,
            in3 => \N__13223\,
            lcout => \c0.rx.n5049\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__13225\,
            in1 => \N__14761\,
            in2 => \_gnd_net_\,
            in3 => \N__12346\,
            lcout => \r_Clock_Count_7_adj_2004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_4_lut_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001010101010"
        )
    port map (
            in0 => \N__18130\,
            in1 => \N__18266\,
            in2 => \N__13509\,
            in3 => \N__18047\,
            lcout => OPEN,
            ltout => \c0.rx.n5923_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.n5923_bdd_4_lut_4_lut_LC_1_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011100011"
        )
    port map (
            in0 => \N__13280\,
            in1 => \N__18267\,
            in2 => \N__12340\,
            in3 => \N__20899\,
            lcout => OPEN,
            ltout => \c0.rx.n5926_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_1_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12337\,
            in3 => \N__18363\,
            lcout => \r_SM_Main_0_adj_2006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_1_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13238\,
            in1 => \N__13344\,
            in2 => \_gnd_net_\,
            in3 => \N__12334\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5253_2_lut_LC_1_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18112\,
            in2 => \_gnd_net_\,
            in3 => \N__13278\,
            lcout => n5490,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5269_3_lut_LC_1_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__13279\,
            in1 => \_gnd_net_\,
            in2 => \N__18131\,
            in3 => \N__20898\,
            lcout => \c0.rx.n5532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_795_LC_1_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18116\,
            in2 => \_gnd_net_\,
            in3 => \N__18048\,
            lcout => OPEN,
            ltout => \c0.rx.n3980_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_1_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000010101"
        )
    port map (
            in0 => \N__18362\,
            in1 => \N__18268\,
            in2 => \N__12373\,
            in3 => \N__12370\,
            lcout => \c0.rx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__13580\,
            in1 => \N__13542\,
            in2 => \N__13485\,
            in3 => \N__12433\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13478\,
            in2 => \_gnd_net_\,
            in3 => \N__13594\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_908_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12432\,
            in2 => \_gnd_net_\,
            in3 => \N__12420\,
            lcout => \c0.n103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_968_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20610\,
            in1 => \N__20718\,
            in2 => \_gnd_net_\,
            in3 => \N__16431\,
            lcout => n1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13476\,
            in2 => \_gnd_net_\,
            in3 => \N__13618\,
            lcout => \c0.byte_transmit_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__13581\,
            in1 => \N__13543\,
            in2 => \N__13486\,
            in3 => \N__12421\,
            lcout => \c0.byte_transmit_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13477\,
            in2 => \_gnd_net_\,
            in3 => \N__13606\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12457\,
            in2 => \N__20354\,
            in3 => \N__16663\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \c0.n4378\,
            clk => \N__35269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16664\,
            in1 => \N__20508\,
            in2 => \_gnd_net_\,
            in3 => \N__12436\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \c0.n4378\,
            carryout => \c0.n4379\,
            clk => \N__35269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_4_lut_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21261\,
            in2 => \_gnd_net_\,
            in3 => \N__12424\,
            lcout => \c0.tx_transmit_N_568_2\,
            ltout => OPEN,
            carryin => \c0.n4379\,
            carryout => \c0.n4380\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_5_lut_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21345\,
            in2 => \_gnd_net_\,
            in3 => \N__12412\,
            lcout => \c0.tx_transmit_N_568_3\,
            ltout => OPEN,
            carryin => \c0.n4380\,
            carryout => \c0.n4381\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_6_lut_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21148\,
            in2 => \_gnd_net_\,
            in3 => \N__12409\,
            lcout => \c0.tx_transmit_N_568_4\,
            ltout => OPEN,
            carryin => \c0.n4381\,
            carryout => \c0.n4382\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_7_lut_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12406\,
            in2 => \_gnd_net_\,
            in3 => \N__12400\,
            lcout => \c0.tx_transmit_N_568_5\,
            ltout => OPEN,
            carryin => \c0.n4382\,
            carryout => \c0.n4383\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_8_lut_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12397\,
            in2 => \_gnd_net_\,
            in3 => \N__12391\,
            lcout => \c0.tx_transmit_N_568_6\,
            ltout => OPEN,
            carryin => \c0.n4383\,
            carryout => \c0.n4384\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_9_lut_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12388\,
            in2 => \_gnd_net_\,
            in3 => \N__12382\,
            lcout => \c0.tx_transmit_N_568_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i23_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000011"
        )
    port map (
            in0 => \N__20763\,
            in1 => \N__13671\,
            in2 => \N__16291\,
            in3 => \N__16672\,
            lcout => data_out_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_985_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18967\,
            in1 => \N__18735\,
            in2 => \_gnd_net_\,
            in3 => \N__19297\,
            lcout => n5077,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_959_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12451\,
            in2 => \_gnd_net_\,
            in3 => \N__13641\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_1793_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5277_4_lut_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__21006\,
            in1 => \N__20324\,
            in2 => \N__16566\,
            in3 => \N__20509\,
            lcout => OPEN,
            ltout => \c0.n5540_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111000000"
        )
    port map (
            in0 => \N__20510\,
            in1 => \N__21379\,
            in2 => \N__12445\,
            in3 => \N__21288\,
            lcout => OPEN,
            ltout => \c0.n5977_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5977_bdd_4_lut_4_lut_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000110100101"
        )
    port map (
            in0 => \N__21380\,
            in1 => \N__20325\,
            in2 => \N__12442\,
            in3 => \N__20511\,
            lcout => \c0.n5980\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_843_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21075\,
            in2 => \_gnd_net_\,
            in3 => \N__21007\,
            lcout => n1760,
            ltout => \n1760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i18_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__15288\,
            in1 => \N__16444\,
            in2 => \N__12439\,
            in3 => \N__16677\,
            lcout => data_out_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19283\,
            in1 => \N__16284\,
            in2 => \_gnd_net_\,
            in3 => \N__20392\,
            lcout => \c0.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_935_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16570\,
            in1 => \N__18805\,
            in2 => \_gnd_net_\,
            in3 => \N__15155\,
            lcout => OPEN,
            ltout => \c0.n1529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_835_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15021\,
            in1 => \N__12496\,
            in2 => \N__12490\,
            in3 => \N__12487\,
            lcout => n5079,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20470\,
            in1 => \N__18979\,
            in2 => \_gnd_net_\,
            in3 => \N__21008\,
            lcout => n7_adj_2002,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_874_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16283\,
            in2 => \_gnd_net_\,
            in3 => \N__16371\,
            lcout => \c0.n1801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__12481\,
            in1 => \N__13978\,
            in2 => \N__16999\,
            in3 => \N__12613\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19342\,
            in1 => \N__15264\,
            in2 => \_gnd_net_\,
            in3 => \N__15415\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__16979\,
            in1 => \N__13977\,
            in2 => \N__12634\,
            in3 => \N__12475\,
            lcout => \r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__13976\,
            in1 => \N__16978\,
            in2 => \N__12595\,
            in3 => \N__12469\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__16977\,
            in1 => \N__12463\,
            in2 => \N__12676\,
            in3 => \N__13979\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__12661\,
            in1 => \N__14025\,
            in2 => \N__17001\,
            in3 => \N__13983\,
            lcout => \r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__12570\,
            in1 => \N__12655\,
            in2 => \N__16998\,
            in3 => \N__13981\,
            lcout => \r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__12537\,
            in1 => \N__12649\,
            in2 => \N__17000\,
            in3 => \N__13982\,
            lcout => \r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__16973\,
            in1 => \N__13980\,
            in2 => \N__12643\,
            in3 => \N__12555\,
            lcout => \r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_805_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__12629\,
            in1 => \N__12611\,
            in2 => \N__12594\,
            in3 => \N__12509\,
            lcout => OPEN,
            ltout => \c0.tx.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i3351_4_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__12569\,
            in1 => \N__12554\,
            in2 => \N__12541\,
            in3 => \N__12536\,
            lcout => n3595,
            ltout => \n3595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__16984\,
            in1 => \N__17051\,
            in2 => \N__12523\,
            in3 => \N__14024\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12510\,
            in1 => \_gnd_net_\,
            in2 => \N__12520\,
            in3 => \N__16985\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__13877\,
            in1 => \N__12788\,
            in2 => \N__12886\,
            in3 => \N__14054\,
            lcout => OPEN,
            ltout => \c0.tx2.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i3348_4_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__12818\,
            in1 => \N__12848\,
            in2 => \N__12718\,
            in3 => \N__13901\,
            lcout => \c0.tx2.n3591\,
            ltout => \c0.tx2.n3591_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i3380_2_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12709\,
            in3 => \N__12748\,
            lcout => \r_SM_Main_2_N_1767_1\,
            ltout => \r_SM_Main_2_N_1767_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__14388\,
            in1 => \N__13860\,
            in2 => \N__12706\,
            in3 => \N__14248\,
            lcout => \r_SM_Main_1_adj_2010\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i6_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__14087\,
            in1 => \_gnd_net_\,
            in2 => \N__14263\,
            in3 => \N__12772\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i4_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12832\,
            in1 => \N__14241\,
            in2 => \_gnd_net_\,
            in3 => \N__14085\,
            lcout => \c0.tx2.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i5_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__14086\,
            in1 => \_gnd_net_\,
            in2 => \N__14262\,
            in3 => \N__12802\,
            lcout => \c0.tx2.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i1_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12865\,
            in1 => \N__14240\,
            in2 => \_gnd_net_\,
            in3 => \N__14084\,
            lcout => \c0.tx2.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_2_lut_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__12703\,
            in1 => \N__12702\,
            in2 => \N__14254\,
            in3 => \N__12679\,
            lcout => n2460,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => \c0.tx2.n4429\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_3_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__12885\,
            in1 => \N__12884\,
            in2 => \N__14258\,
            in3 => \N__12859\,
            lcout => n2399,
            ltout => OPEN,
            carryin => \c0.tx2.n4429\,
            carryout => \c0.tx2.n4430\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_4_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__13879\,
            in1 => \N__13878\,
            in2 => \N__14255\,
            in3 => \N__12856\,
            lcout => n2395,
            ltout => OPEN,
            carryin => \c0.tx2.n4430\,
            carryout => \c0.tx2.n4431\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_5_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14056\,
            in1 => \N__14055\,
            in2 => \N__14259\,
            in3 => \N__12853\,
            lcout => n2392,
            ltout => OPEN,
            carryin => \c0.tx2.n4431\,
            carryout => \c0.tx2.n4432\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_6_lut_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__12850\,
            in1 => \N__12849\,
            in2 => \N__14256\,
            in3 => \N__12823\,
            lcout => n2382,
            ltout => OPEN,
            carryin => \c0.tx2.n4432\,
            carryout => \c0.tx2.n4433\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_7_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__12820\,
            in1 => \N__12819\,
            in2 => \N__14260\,
            in3 => \N__12793\,
            lcout => n2379,
            ltout => OPEN,
            carryin => \c0.tx2.n4433\,
            carryout => \c0.tx2.n4434\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_8_lut_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__12790\,
            in1 => \N__12789\,
            in2 => \N__14257\,
            in3 => \N__12763\,
            lcout => n2376,
            ltout => OPEN,
            carryin => \c0.tx2.n4434\,
            carryout => \c0.tx2.n4435\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_9_lut_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__13903\,
            in1 => \N__13902\,
            in2 => \N__14261\,
            in3 => \N__12760\,
            lcout => n2372,
            ltout => OPEN,
            carryin => \c0.tx2.n4435\,
            carryout => \c0.tx2.n4436\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_10_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__12756\,
            in1 => \N__12757\,
            in2 => \N__14252\,
            in3 => \N__12730\,
            lcout => n2369,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000100"
        )
    port map (
            in0 => \N__13807\,
            in1 => \N__13854\,
            in2 => \N__14250\,
            in3 => \N__12904\,
            lcout => \r_SM_Main_0_adj_2011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__12955\,
            in1 => \N__12892\,
            in2 => \N__15602\,
            in3 => \N__15624\,
            lcout => \c0.tx2.n5947\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n5947_bdd_4_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__13003\,
            in1 => \N__15594\,
            in2 => \N__12925\,
            in3 => \N__12916\,
            lcout => \c0.tx2.n5950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1104_4_lut_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__14391\,
            in1 => \N__15783\,
            in2 => \N__14322\,
            in3 => \N__13805\,
            lcout => n1345,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_4_lut_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__15782\,
            in1 => \N__13852\,
            in2 => \N__14249\,
            in3 => \N__14392\,
            lcout => \c0.tx2.n1592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i817_2_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34747\,
            in2 => \_gnd_net_\,
            in3 => \N__32079\,
            lcout => \c0.n1058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__13806\,
            in1 => \N__13853\,
            in2 => \N__14251\,
            in3 => \N__14393\,
            lcout => \r_SM_Main_2_adj_2009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5563_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__15997\,
            in1 => \N__32316\,
            in2 => \N__35440\,
            in3 => \N__33115\,
            lcout => \c0.n5953\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__13048\,
            in1 => \N__14511\,
            in2 => \N__14284\,
            in3 => \N__18916\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => \N__12993\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14509\,
            in1 => \N__13046\,
            in2 => \N__14452\,
            in3 => \N__22882\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => \N__12993\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14510\,
            in1 => \N__13047\,
            in2 => \N__13096\,
            in3 => \N__14458\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => \N__12993\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5326_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__17732\,
            in1 => \N__33287\,
            in2 => \N__32544\,
            in3 => \N__27661\,
            lcout => OPEN,
            ltout => \c0.n5665_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5665_bdd_4_lut_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__25702\,
            in1 => \N__24756\,
            in2 => \N__12949\,
            in3 => \N__32444\,
            lcout => OPEN,
            ltout => \c0.n5372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5331_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__32099\,
            in1 => \N__34805\,
            in2 => \N__12946\,
            in3 => \N__13123\,
            lcout => \c0.n5659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5310_4_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100111111"
        )
    port map (
            in0 => \N__33288\,
            in1 => \N__13056\,
            in2 => \N__14533\,
            in3 => \N__32443\,
            lcout => \c0.FRAME_MATCHER_wait_for_transmission_N_909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5935_bdd_4_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32445\,
            in1 => \N__27139\,
            in2 => \N__14407\,
            in3 => \N__19681\,
            lcout => \c0.n5938\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i140_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__34362\,
            in1 => \N__14639\,
            in2 => \N__17534\,
            in3 => \_gnd_net_\,
            lcout => data_in_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i148_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15861\,
            in2 => \N__14646\,
            in3 => \N__34361\,
            lcout => data_in_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__33246\,
            in1 => \N__13138\,
            in2 => \N__14593\,
            in3 => \N__32526\,
            lcout => OPEN,
            ltout => \c0.n5971_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5971_bdd_4_lut_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32527\,
            in1 => \N__30872\,
            in2 => \N__12928\,
            in3 => \N__19939\,
            lcout => \c0.n5974\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5395_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__32108\,
            in1 => \N__16051\,
            in2 => \N__34827\,
            in3 => \N__14608\,
            lcout => OPEN,
            ltout => \c0.n5725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5725_bdd_4_lut_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__25822\,
            in1 => \N__34811\,
            in2 => \N__13063\,
            in3 => \N__14542\,
            lcout => OPEN,
            ltout => \c0.n5728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__14526\,
            in1 => \N__13057\,
            in2 => \N__13012\,
            in3 => \N__13009\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => \N__12994\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i132_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26831\,
            in1 => \N__17535\,
            in2 => \_gnd_net_\,
            in3 => \N__34294\,
            lcout => data_in_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i42_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36787\,
            in1 => \N__36041\,
            in2 => \N__17436\,
            in3 => \N__13423\,
            lcout => \c0.data_in_field_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5440_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__33274\,
            in1 => \N__26271\,
            in2 => \N__24964\,
            in3 => \N__32516\,
            lcout => OPEN,
            ltout => \c0.n5803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5803_bdd_4_lut_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32517\,
            in1 => \N__25057\,
            in2 => \N__12958\,
            in3 => \N__19984\,
            lcout => \c0.n5426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i22_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__16111\,
            in1 => \N__36040\,
            in2 => \N__37000\,
            in3 => \N__23739\,
            lcout => \c0.data_in_field_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i149_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26795\,
            in1 => \N__37334\,
            in2 => \_gnd_net_\,
            in3 => \N__34295\,
            lcout => data_in_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_909_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32022\,
            in1 => \N__29535\,
            in2 => \_gnd_net_\,
            in3 => \N__22245\,
            lcout => \c0.n16_adj_1922\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i146_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__13137\,
            in1 => \N__37124\,
            in2 => \N__36261\,
            in3 => \N__20086\,
            lcout => \c0.data_in_frame_18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i156_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34151\,
            in1 => \N__14797\,
            in2 => \_gnd_net_\,
            in3 => \N__15853\,
            lcout => data_in_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5671_bdd_4_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__14803\,
            in1 => \N__17509\,
            in2 => \N__32593\,
            in3 => \N__25501\,
            lcout => \c0.n5369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5495_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33236\,
            in1 => \N__23623\,
            in2 => \N__32594\,
            in3 => \N__26953\,
            lcout => \c0.n5869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5959_bdd_4_lut_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32587\,
            in1 => \N__14692\,
            in2 => \N__13105\,
            in3 => \N__25009\,
            lcout => \c0.n5962\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i148_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__13083\,
            in1 => \N__37125\,
            in2 => \N__36262\,
            in3 => \N__14647\,
            lcout => \c0.data_in_frame_18_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__13240\,
            in1 => \N__14882\,
            in2 => \_gnd_net_\,
            in3 => \N__13069\,
            lcout => \r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__18138\,
            in2 => \N__18355\,
            in3 => \N__18281\,
            lcout => \r_SM_Main_2_adj_2005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_878_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19800\,
            in1 => \N__22573\,
            in2 => \N__24434\,
            in3 => \N__28030\,
            lcout => \c0.n15_adj_1894\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14912\,
            in1 => \N__13192\,
            in2 => \_gnd_net_\,
            in3 => \N__13241\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13186\,
            in1 => \N__13243\,
            in2 => \_gnd_net_\,
            in3 => \N__13375\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_4_lut_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__18055\,
            in1 => \N__18137\,
            in2 => \N__18354\,
            in3 => \N__18280\,
            lcout => \c0.rx.n2157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13239\,
            in1 => \N__13399\,
            in2 => \_gnd_net_\,
            in3 => \N__13174\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13242\,
            in1 => \N__13309\,
            in2 => \_gnd_net_\,
            in3 => \N__13168\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_794_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__14766\,
            in1 => \N__13162\,
            in2 => \N__14884\,
            in3 => \N__13351\,
            lcout => \c0.rx.r_SM_Main_2_N_1824_2\,
            ltout => \c0.rx.r_SM_Main_2_N_1824_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18328\,
            in2 => \N__13156\,
            in3 => \N__18276\,
            lcout => n4474,
            ltout => \n4474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_796_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__18329\,
            in1 => \N__13147\,
            in2 => \N__13141\,
            in3 => \N__13281\,
            lcout => OPEN,
            ltout => \c0.rx.n4_adj_1866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3748_2_lut_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13453\,
            in3 => \N__13222\,
            lcout => \c0.rx.n4011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i42_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23956\,
            in1 => \_gnd_net_\,
            in2 => \N__34363\,
            in3 => \N__13410\,
            lcout => data_in_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_793_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13396\,
            in2 => \_gnd_net_\,
            in3 => \N__13372\,
            lcout => \c0.rx.n37\,
            ltout => \c0.rx.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i4_4_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14701\,
            in1 => \N__13340\,
            in2 => \N__13312\,
            in3 => \N__13307\,
            lcout => \r_SM_Main_2_N_1830_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__18247\,
            in1 => \N__18111\,
            in2 => \N__18356\,
            in3 => \N__18049\,
            lcout => \c0.rx.n2213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13258\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_29_i4_2_lut_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14934\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5_4_lut_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18110\,
            in1 => \N__18246\,
            in2 => \N__20915\,
            in3 => \N__14729\,
            lcout => OPEN,
            ltout => \n12_adj_1995_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_1012_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__18337\,
            in1 => \N__14848\,
            in2 => \N__13252\,
            in3 => \N__13249\,
            lcout => n16_adj_1993,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_3_lut_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14933\,
            in1 => \N__18176\,
            in2 => \_gnd_net_\,
            in3 => \N__14962\,
            lcout => \c0.rx.n3573\,
            ltout => \c0.rx.n3573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2073_2_lut_3_lut_LC_2_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__18248\,
            in1 => \_gnd_net_\,
            in2 => \N__13492\,
            in3 => \N__14988\,
            lcout => \c0.rx.n2317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i36_LC_2_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34152\,
            in1 => \N__26584\,
            in2 => \_gnd_net_\,
            in3 => \N__17669\,
            lcout => data_in_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20639\,
            in1 => \N__20739\,
            in2 => \N__18817\,
            in3 => \N__16430\,
            lcout => n4_adj_1988,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_1794_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13549\,
            in1 => \N__13541\,
            in2 => \N__13723\,
            in3 => \N__13656\,
            lcout => \c0.tx_transmit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_902_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14818\,
            in1 => \N__15036\,
            in2 => \N__15082\,
            in3 => \N__15181\,
            lcout => OPEN,
            ltout => \c0.n20_adj_1918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_906_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15057\,
            in1 => \N__15111\,
            in2 => \N__13489\,
            in3 => \N__13459\,
            lcout => n21_adj_1999,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_939_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13710\,
            in1 => \N__19167\,
            in2 => \_gnd_net_\,
            in3 => \N__13655\,
            lcout => \c0.n87\,
            ltout => \c0.n87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__13540\,
            in1 => \N__13582\,
            in2 => \N__13462\,
            in3 => \N__13561\,
            lcout => \c0.byte_transmit_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15096\,
            in2 => \_gnd_net_\,
            in3 => \N__14835\,
            lcout => \c0.n16_adj_1909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i14_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19174\,
            in1 => \N__20730\,
            in2 => \N__18406\,
            in3 => \N__19033\,
            lcout => data_out_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_913_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13617\,
            in1 => \N__13605\,
            in2 => \_gnd_net_\,
            in3 => \N__13593\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i119_2_lut_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13579\,
            in2 => \_gnd_net_\,
            in3 => \N__13560\,
            lcout => \c0.n109\,
            ltout => \c0.n109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5298_3_lut_4_lut_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__13702\,
            in1 => \N__13539\,
            in2 => \N__13519\,
            in3 => \N__13654\,
            lcout => n4315,
            ltout => \n4315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i12_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__18427\,
            in1 => \N__16565\,
            in2 => \N__13516\,
            in3 => \N__19175\,
            lcout => data_out_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i29_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__16711\,
            in1 => \N__13777\,
            in2 => \N__16144\,
            in3 => \N__16673\,
            lcout => data_out_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i15_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19034\,
            in1 => \N__18382\,
            in2 => \N__20640\,
            in3 => \N__19176\,
            lcout => data_out_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i10_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__19029\,
            in1 => \N__16807\,
            in2 => \N__18472\,
            in3 => \N__19179\,
            lcout => data_out_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i6_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19178\,
            in1 => \N__21109\,
            in2 => \N__18535\,
            in3 => \N__19032\,
            lcout => data_out_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i5_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19031\,
            in1 => \N__18553\,
            in2 => \N__18749\,
            in3 => \N__19181\,
            lcout => data_out_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i27_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__16227\,
            in1 => \N__16186\,
            in2 => \N__15493\,
            in3 => \N__16666\,
            lcout => data_out_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i4_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__19030\,
            in1 => \N__21012\,
            in2 => \N__18574\,
            in3 => \N__19180\,
            lcout => data_out_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_943_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__19177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19028\,
            lcout => n4316,
            ltout => \n4316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i20_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011000101"
        )
    port map (
            in0 => \N__20979\,
            in1 => \N__15357\,
            in2 => \N__13684\,
            in3 => \N__15163\,
            lcout => data_out_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i25_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__15249\,
            in1 => \N__13747\,
            in2 => \N__13681\,
            in3 => \N__16665\,
            lcout => data_out_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_4_lut_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__13724\,
            in1 => \N__17121\,
            in2 => \N__17002\,
            in3 => \N__17062\,
            lcout => n1442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i21_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100101"
        )
    port map (
            in0 => \N__13672\,
            in1 => \N__13762\,
            in2 => \N__15274\,
            in3 => \N__16671\,
            lcout => data_out_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110100"
        )
    port map (
            in0 => \N__17122\,
            in1 => \N__13735\,
            in2 => \N__13657\,
            in3 => \N__16996\,
            lcout => tx_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13776\,
            in1 => \N__20393\,
            in2 => \_gnd_net_\,
            in3 => \N__13761\,
            lcout => OPEN,
            ltout => \c0.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__21186\,
            in1 => \N__18706\,
            in2 => \N__13753\,
            in3 => \N__20683\,
            lcout => OPEN,
            ltout => \tx_data_4_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__16827\,
            in1 => \_gnd_net_\,
            in2 => \N__13750\,
            in3 => \N__19340\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i16_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__16416\,
            in1 => \N__19220\,
            in2 => \N__18628\,
            in3 => \N__19058\,
            lcout => data_out_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16474\,
            in1 => \N__19300\,
            in2 => \N__16378\,
            in3 => \N__21079\,
            lcout => n8_adj_2001,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14022\,
            in2 => \_gnd_net_\,
            in3 => \N__13995\,
            lcout => \c0.tx.r_SM_Main_2_N_1767_1\,
            ltout => \c0.tx.r_SM_Main_2_N_1767_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5288_3_lut_4_lut_4_lut_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000100010"
        )
    port map (
            in0 => \N__13725\,
            in1 => \N__17116\,
            in2 => \N__13738\,
            in3 => \N__17058\,
            lcout => n5041,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17120\,
            in1 => \N__17049\,
            in2 => \N__16997\,
            in3 => \N__15405\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__15404\,
            in1 => \N__16972\,
            in2 => \N__17060\,
            in3 => \N__17119\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i29_4_lut_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__13729\,
            in1 => \N__17098\,
            in2 => \N__15385\,
            in3 => \N__15403\,
            lcout => OPEN,
            ltout => \c0.tx.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100110000"
        )
    port map (
            in0 => \N__15406\,
            in1 => \N__16967\,
            in2 => \N__14029\,
            in3 => \N__17059\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1066_2_lut_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17097\,
            in2 => \_gnd_net_\,
            in3 => \N__17044\,
            lcout => n1307,
            ltout => \n1307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_802_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__16949\,
            in1 => \N__14023\,
            in2 => \N__13999\,
            in3 => \N__13996\,
            lcout => n4221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011100000"
        )
    port map (
            in0 => \N__17118\,
            in1 => \N__17045\,
            in2 => \N__13927\,
            in3 => \N__13942\,
            lcout => OPEN,
            ltout => \n4_adj_2003_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Done_44_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111110000"
        )
    port map (
            in0 => \N__13926\,
            in1 => \N__13936\,
            in2 => \N__13930\,
            in3 => \N__16968\,
            lcout => n4155,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i7_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__14097\,
            in1 => \_gnd_net_\,
            in2 => \N__13912\,
            in3 => \N__14234\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i2_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__14233\,
            in1 => \N__13885\,
            in2 => \_gnd_net_\,
            in3 => \N__14096\,
            lcout => \c0.tx2.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_3_lut_4_lut_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__13855\,
            in1 => \N__14232\,
            in2 => \N__14389\,
            in3 => \N__13795\,
            lcout => \c0.tx2.n2218\,
            ltout => \c0.tx2.n2218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2075_2_lut_3_lut_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14368\,
            in2 => \N__14326\,
            in3 => \N__14323\,
            lcout => \c0.tx2.n2319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5953_bdd_4_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32319\,
            in1 => \N__28861\,
            in2 => \N__14296\,
            in3 => \N__27433\,
            lcout => \c0.n5956\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i3_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__14269\,
            in1 => \N__14207\,
            in2 => \_gnd_net_\,
            in3 => \N__14101\,
            lcout => \c0.tx2.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23864\,
            in1 => \N__34283\,
            in2 => \_gnd_net_\,
            in3 => \N__27892\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i93_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34282\,
            in1 => \N__28708\,
            in2 => \_gnd_net_\,
            in3 => \N__27038\,
            lcout => data_in_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_525_526__i1_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33116\,
            in2 => \N__15823\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => \c0.n4400\,
            clk => \N__35307\,
            ce => \N__15733\,
            sr => \N__15721\
        );

    \c0.byte_transmit_counter2_525_526__i2_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32320\,
            in2 => \_gnd_net_\,
            in3 => \N__14038\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \c0.n4400\,
            carryout => \c0.n4401\,
            clk => \N__35307\,
            ce => \N__15733\,
            sr => \N__15721\
        );

    \c0.byte_transmit_counter2_525_526__i3_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32098\,
            in2 => \_gnd_net_\,
            in3 => \N__14035\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \c0.n4401\,
            carryout => \c0.n4402\,
            clk => \N__35307\,
            ce => \N__15733\,
            sr => \N__15721\
        );

    \c0.byte_transmit_counter2_525_526__i4_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34762\,
            in2 => \_gnd_net_\,
            in3 => \N__14032\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \c0.n4402\,
            carryout => \c0.n4403\,
            clk => \N__35307\,
            ce => \N__15733\,
            sr => \N__15721\
        );

    \c0.byte_transmit_counter2_525_526__i5_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14505\,
            in2 => \_gnd_net_\,
            in3 => \N__14536\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => \N__15733\,
            sr => \N__15721\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5455_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__32097\,
            in1 => \N__21751\,
            in2 => \N__34800\,
            in3 => \N__21775\,
            lcout => OPEN,
            ltout => \c0.n5785_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5785_bdd_4_lut_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__21853\,
            in1 => \N__34761\,
            in2 => \N__14470\,
            in3 => \N__14467\,
            lcout => \c0.n5788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5965_bdd_4_lut_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32318\,
            in1 => \N__28396\,
            in2 => \N__17386\,
            in3 => \N__28438\,
            lcout => \c0.n5968\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34219\,
            in1 => \N__17686\,
            in2 => \_gnd_net_\,
            in3 => \N__23305\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35311\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5809_bdd_4_lut_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32317\,
            in1 => \N__30358\,
            in2 => \N__19417\,
            in3 => \N__20119\,
            lcout => \c0.n5363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i160_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__14427\,
            in1 => \N__20164\,
            in2 => \N__37003\,
            in3 => \N__36199\,
            lcout => \c0.data_in_frame_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5548_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__16129\,
            in1 => \N__33181\,
            in2 => \N__14559\,
            in3 => \N__32446\,
            lcout => \c0.n5935\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i102_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36798\,
            in1 => \N__36198\,
            in2 => \N__16039\,
            in3 => \N__15963\,
            lcout => \c0.data_in_field_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i158_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34215\,
            in1 => \N__14782\,
            in2 => \_gnd_net_\,
            in3 => \N__24505\,
            lcout => data_in_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i94_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__16035\,
            in1 => \N__34216\,
            in2 => \N__26983\,
            in3 => \_gnd_net_\,
            lcout => data_in_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5941_bdd_4_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32447\,
            in1 => \N__23932\,
            in2 => \N__18904\,
            in3 => \N__20050\,
            lcout => \c0.n5944\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i86_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26978\,
            in1 => \N__34217\,
            in2 => \_gnd_net_\,
            in3 => \N__27528\,
            lcout => data_in_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_3_lut_4_lut_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14614\,
            in1 => \N__22198\,
            in2 => \N__22399\,
            in3 => \N__22165\,
            lcout => \c0.n23_adj_1931\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i14_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__24154\,
            in1 => \N__36272\,
            in2 => \N__37002\,
            in3 => \N__21707\,
            lcout => \c0.data_in_field_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i12_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__21875\,
            in1 => \N__22375\,
            in2 => \N__37001\,
            in3 => \N__36273\,
            lcout => \c0.data_in_field_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i159_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36271\,
            in1 => \N__36791\,
            in2 => \N__14560\,
            in3 => \N__17370\,
            lcout => \c0.data_in_frame_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5743_bdd_4_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32543\,
            in1 => \N__17422\,
            in2 => \N__19852\,
            in3 => \N__29302\,
            lcout => \c0.n5456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_975_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__21579\,
            in2 => \_gnd_net_\,
            in3 => \N__19935\,
            lcout => \c0.n1893\,
            ltout => \c0.n1893_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_907_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19503\,
            in1 => \N__14635\,
            in2 => \N__14617\,
            in3 => \N__28395\,
            lcout => \c0.n20_adj_1921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_849_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17421\,
            in1 => \N__21874\,
            in2 => \N__17508\,
            in3 => \N__17277\,
            lcout => \c0.n1821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_846_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15958\,
            in1 => \N__31344\,
            in2 => \_gnd_net_\,
            in3 => \N__14689\,
            lcout => \c0.n5072\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_891_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19518\,
            in1 => \N__23638\,
            in2 => \N__19804\,
            in3 => \N__25810\,
            lcout => \c0.n24_adj_1907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i132_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36786\,
            in1 => \N__36013\,
            in2 => \N__26835\,
            in3 => \N__14690\,
            lcout => \c0.data_in_field_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5737_bdd_4_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__14602\,
            in1 => \N__30271\,
            in2 => \N__32595\,
            in3 => \N__20017\,
            lcout => \c0.n5459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24640\,
            in1 => \N__17435\,
            in2 => \N__24223\,
            in3 => \N__28437\,
            lcout => \c0.n22_adj_1881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5385_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33237\,
            in1 => \N__23554\,
            in2 => \N__32545\,
            in3 => \N__15701\,
            lcout => \c0.n5737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i82_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__15702\,
            in1 => \N__28573\,
            in2 => \N__36200\,
            in3 => \N__37123\,
            lcout => \c0.data_in_field_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i154_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__14586\,
            in1 => \N__36006\,
            in2 => \N__37226\,
            in3 => \N__17878\,
            lcout => \c0.data_in_frame_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i120_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36005\,
            in1 => \N__37116\,
            in2 => \N__21667\,
            in3 => \N__17725\,
            lcout => \c0.data_in_field_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i20_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23354\,
            in1 => \N__17845\,
            in2 => \N__37227\,
            in3 => \N__36010\,
            lcout => \c0.data_in_field_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_832_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15700\,
            in1 => \N__23353\,
            in2 => \N__23740\,
            in3 => \N__14691\,
            lcout => \c0.n2036\,
            ltout => \c0.n2036_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_834_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14671\,
            in3 => \N__24956\,
            lcout => OPEN,
            ltout => \c0.n5273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19470\,
            in1 => \N__24579\,
            in2 => \N__14668\,
            in3 => \N__25939\,
            lcout => \c0.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34030\,
            in1 => \N__31731\,
            in2 => \_gnd_net_\,
            in3 => \N__22371\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i152_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__14661\,
            in1 => \N__36146\,
            in2 => \N__37203\,
            in3 => \N__26043\,
            lcout => \c0.data_in_frame_18_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i151_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34029\,
            in1 => \N__17359\,
            in2 => \_gnd_net_\,
            in3 => \N__24211\,
            lcout => data_in_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i127_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23672\,
            in1 => \N__34031\,
            in2 => \_gnd_net_\,
            in3 => \N__17934\,
            lcout => data_in_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5336_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33117\,
            in1 => \N__19834\,
            in2 => \N__32589\,
            in3 => \N__23007\,
            lcout => \c0.n5671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31439\,
            in1 => \N__31528\,
            in2 => \_gnd_net_\,
            in3 => \N__33881\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__14793\,
            in1 => \N__20859\,
            in2 => \N__20930\,
            in3 => \N__17964\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i138_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33880\,
            in1 => \N__20798\,
            in2 => \_gnd_net_\,
            in3 => \N__20084\,
            lcout => data_in_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33885\,
            in1 => \N__16107\,
            in2 => \_gnd_net_\,
            in3 => \N__27967\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33882\,
            in1 => \N__23312\,
            in2 => \_gnd_net_\,
            in3 => \N__17837\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__20911\,
            in1 => \N__14778\,
            in2 => \N__20863\,
            in3 => \N__16170\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__14874\,
            in1 => \N__14765\,
            in2 => \N__14913\,
            in3 => \N__14731\,
            lcout => \c0.rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_26_i4_2_lut_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__14965\,
            in1 => \N__14938\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n4_adj_1990,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__14940\,
            in1 => \_gnd_net_\,
            in2 => \N__18184\,
            in3 => \N__14967\,
            lcout => \c0.rx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35352\,
            ce => \N__14992\,
            sr => \N__14977\
        );

    \c0.rx.r_Bit_Index_i1_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__14968\,
            in1 => \N__18180\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35352\,
            ce => \N__14992\,
            sr => \N__14977\
        );

    \c0.rx.equal_27_i4_2_lut_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14941\,
            in3 => \N__14964\,
            lcout => n4_adj_1986,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3101_2_lut_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14966\,
            in1 => \N__14939\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n3342,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_797_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14914\,
            in2 => \_gnd_net_\,
            in3 => \N__14883\,
            lcout => n8_adj_1996,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4002_1_lut_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16891\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i0_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19027\,
            in2 => \N__15211\,
            in3 => \_gnd_net_\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \c0.n4404\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i1_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14836\,
            in2 => \_gnd_net_\,
            in3 => \N__14824\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \c0.n4404\,
            carryout => \c0.n4405\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i2_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15223\,
            in2 => \_gnd_net_\,
            in3 => \N__14821\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \c0.n4405\,
            carryout => \c0.n4406\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i3_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14817\,
            in2 => \_gnd_net_\,
            in3 => \N__15115\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \c0.n4406\,
            carryout => \c0.n4407\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i4_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15112\,
            in2 => \_gnd_net_\,
            in3 => \N__15100\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \c0.n4407\,
            carryout => \c0.n4408\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i5_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15097\,
            in2 => \_gnd_net_\,
            in3 => \N__15085\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \c0.n4408\,
            carryout => \c0.n4409\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i6_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15081\,
            in2 => \_gnd_net_\,
            in3 => \N__15067\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \c0.n4409\,
            carryout => \c0.n4410\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i7_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15193\,
            in2 => \_gnd_net_\,
            in3 => \N__15064\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \c0.n4410\,
            carryout => \c0.n4411\,
            clk => \N__35280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i8_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15061\,
            in3 => \N__15046\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => \c0.n4412\,
            clk => \N__35273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i9_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15235\,
            in3 => \N__15043\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \c0.n4412\,
            carryout => \c0.n4413\,
            clk => \N__35273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i10_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15037\,
            in2 => \_gnd_net_\,
            in3 => \N__15040\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i19_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__15025\,
            in1 => \N__16246\,
            in2 => \N__15004\,
            in3 => \N__16678\,
            lcout => data_out_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_944_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16796\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16273\,
            lcout => n4_adj_2000,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_894_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16797\,
            in2 => \_gnd_net_\,
            in3 => \N__21077\,
            lcout => n5063,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5267_4_lut_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__15126\,
            in1 => \N__20679\,
            in2 => \N__15250\,
            in3 => \N__20391\,
            lcout => \c0.n5501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_893_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15231\,
            in1 => \N__15222\,
            in2 => \N__15210\,
            in3 => \N__15192\,
            lcout => \c0.n18_adj_1908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_942_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16469\,
            in2 => \_gnd_net_\,
            in3 => \N__19299\,
            lcout => OPEN,
            ltout => \n5086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i31_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__16669\,
            in1 => \N__15175\,
            in2 => \N__15166\,
            in3 => \N__20784\,
            lcout => data_out_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i22_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__16204\,
            in1 => \N__16198\,
            in2 => \N__20983\,
            in3 => \N__16668\,
            lcout => data_out_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_967_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18806\,
            in1 => \N__15162\,
            in2 => \N__16513\,
            in3 => \N__16558\,
            lcout => n5156,
            ltout => \n5156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i17_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__19240\,
            in1 => \N__15127\,
            in2 => \N__15130\,
            in3 => \N__16667\,
            lcout => data_out_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15376\,
            in1 => \N__21108\,
            in2 => \_gnd_net_\,
            in3 => \N__19298\,
            lcout => n8_adj_1997,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i32_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101101000001"
        )
    port map (
            in0 => \N__16670\,
            in1 => \N__16470\,
            in2 => \N__15370\,
            in3 => \N__15342\,
            lcout => data_out_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5254_4_lut_4_lut_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__20409\,
            in1 => \N__15297\,
            in2 => \N__15358\,
            in3 => \N__20572\,
            lcout => \c0.n5519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15343\,
            in1 => \N__20407\,
            in2 => \_gnd_net_\,
            in3 => \N__15309\,
            lcout => \c0.n17_adj_1961\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i24_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__15310\,
            in1 => \N__15328\,
            in2 => \N__15319\,
            in3 => \N__16679\,
            lcout => data_out_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i28_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010110001"
        )
    port map (
            in0 => \N__16680\,
            in1 => \N__15486\,
            in2 => \N__15301\,
            in3 => \N__16690\,
            lcout => data_out_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5227_4_lut_4_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__20408\,
            in1 => \N__15289\,
            in2 => \N__16308\,
            in3 => \N__20571\,
            lcout => \c0.n5531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_934_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20638\,
            in1 => \N__19296\,
            in2 => \_gnd_net_\,
            in3 => \N__16415\,
            lcout => n4_adj_2007,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n5719_bdd_4_lut_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__15265\,
            in1 => \N__17234\,
            in2 => \N__15436\,
            in3 => \N__17158\,
            lcout => \c0.tx.n5722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i932_4_lut_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100100010"
        )
    port map (
            in0 => \N__20412\,
            in1 => \N__21408\,
            in2 => \N__15466\,
            in3 => \N__20580\,
            lcout => OPEN,
            ltout => \c0.n1173_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__21189\,
            in1 => \N__15451\,
            in2 => \N__15442\,
            in3 => \N__21313\,
            lcout => OPEN,
            ltout => \tx_data_0_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15435\,
            in1 => \_gnd_net_\,
            in2 => \N__15439\,
            in3 => \N__19341\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_4_lut_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010010011001"
        )
    port map (
            in0 => \N__21407\,
            in1 => \N__21312\,
            in2 => \N__16765\,
            in3 => \N__20579\,
            lcout => OPEN,
            ltout => \c0.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__21230\,
            in1 => \N__15424\,
            in2 => \N__15418\,
            in3 => \N__21188\,
            lcout => \tx_data_1_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__15676\,
            in1 => \N__17237\,
            in2 => \N__17191\,
            in3 => \N__15666\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__15665\,
            in1 => \N__17186\,
            in2 => \_gnd_net_\,
            in3 => \N__15675\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_799_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__17050\,
            in1 => \N__17099\,
            in2 => \N__16983\,
            in3 => \N__15402\,
            lcout => n2200,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_3_lut_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17150\,
            in1 => \N__17235\,
            in2 => \_gnd_net_\,
            in3 => \N__17185\,
            lcout => \c0.tx.n3507\,
            ltout => \c0.tx.n3507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2063_3_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17100\,
            in2 => \N__15679\,
            in3 => \N__15664\,
            lcout => n2307,
            ltout => \n2307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__15667\,
            in1 => \N__15649\,
            in2 => \N__15652\,
            in3 => \N__17152\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i573_2_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17236\,
            in2 => \_gnd_net_\,
            in3 => \N__17190\,
            lcout => n805,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15572\,
            in2 => \_gnd_net_\,
            in3 => \N__15639\,
            lcout => \c0.tx2.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35302\,
            ce => \N__15508\,
            sr => \N__15499\
        );

    \c0.tx2.r_Bit_Index_i2_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__15640\,
            in1 => \_gnd_net_\,
            in2 => \N__15590\,
            in3 => \N__15530\,
            lcout => \c0.tx2.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35302\,
            ce => \N__15508\,
            sr => \N__15499\
        );

    \c0.i1_2_lut_adj_847_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20471\,
            in2 => \_gnd_net_\,
            in3 => \N__21123\,
            lcout => n5153,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3173_2_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15756\,
            in2 => \_gnd_net_\,
            in3 => \N__15781\,
            lcout => \c0.n3414\,
            ltout => \c0.n3414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_1801_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__36482\,
            in1 => \N__15822\,
            in2 => \N__15469\,
            in3 => \N__17320\,
            lcout => \c0.r_SM_Main_2_N_1770_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5430_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33138\,
            in1 => \N__26101\,
            in2 => \N__32506\,
            in3 => \N__31348\,
            lcout => \c0.n5791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011101111"
        )
    port map (
            in0 => \N__15829\,
            in1 => \N__15821\,
            in2 => \N__36636\,
            in3 => \N__17319\,
            lcout => \c0.FRAME_MATCHER_wait_for_transmission\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i489_3_lut_4_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__15780\,
            in1 => \N__15757\,
            in2 => \N__36635\,
            in3 => \N__17318\,
            lcout => \c0.n195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5475_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33139\,
            in1 => \N__28024\,
            in2 => \N__32507\,
            in3 => \N__31069\,
            lcout => OPEN,
            ltout => \c0.n5845_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5845_bdd_4_lut_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32315\,
            in1 => \N__31585\,
            in2 => \N__15724\,
            in3 => \N__21997\,
            lcout => \c0.n5411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i118_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34075\,
            in1 => \N__20218\,
            in2 => \_gnd_net_\,
            in3 => \N__19433\,
            lcout => data_in_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5293_2_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__36437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17317\,
            lcout => \c0.n2275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_810_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23432\,
            in2 => \_gnd_net_\,
            in3 => \N__15709\,
            lcout => \c0.n1918\,
            ltout => \c0.n1918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_995_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22622\,
            in1 => \N__17754\,
            in2 => \N__15685\,
            in3 => \N__31954\,
            lcout => \c0.n5192\,
            ltout => \c0.n5192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_adj_881_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23750\,
            in2 => \N__15682\,
            in3 => \N__23372\,
            lcout => OPEN,
            ltout => \c0.n30_adj_1897_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_923_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17578\,
            in1 => \N__25774\,
            in2 => \N__15919\,
            in3 => \N__25809\,
            lcout => OPEN,
            ltout => \c0.n36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26284\,
            in1 => \N__19387\,
            in2 => \N__15916\,
            in3 => \N__22009\,
            lcout => \c0.n5277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_917_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15910\,
            in1 => \N__21624\,
            in2 => \N__26113\,
            in3 => \N__30511\,
            lcout => \c0.n21_adj_1928\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25885\,
            in1 => \N__25381\,
            in2 => \N__23023\,
            in3 => \N__24081\,
            lcout => \c0.n5080\,
            ltout => \c0.n5080_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_911_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29890\,
            in1 => \N__19669\,
            in2 => \N__15913\,
            in3 => \N__21993\,
            lcout => \c0.n24_adj_1924\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_853_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32913\,
            in2 => \_gnd_net_\,
            in3 => \N__22830\,
            lcout => \c0.n1990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_916_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24913\,
            in1 => \N__15904\,
            in2 => \N__30267\,
            in3 => \N__15895\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1927_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_921_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__15889\,
            in1 => \N__15883\,
            in2 => \N__15877\,
            in3 => \N__15973\,
            lcout => \c0.n23_adj_1932\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_904_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15874\,
            in1 => \N__24580\,
            in2 => \N__15865\,
            in3 => \N__27225\,
            lcout => \c0.n27_adj_1919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i72_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__36058\,
            in1 => \N__22468\,
            in2 => \N__36650\,
            in3 => \N__17499\,
            lcout => \c0.data_in_field_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i83_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__22769\,
            in1 => \N__36501\,
            in2 => \N__31639\,
            in3 => \N__36061\,
            lcout => \c0.data_in_field_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i145_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__36057\,
            in1 => \N__16011\,
            in2 => \N__36649\,
            in3 => \N__33477\,
            lcout => \c0.data_in_frame_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i100_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__21581\,
            in1 => \N__36500\,
            in2 => \N__31840\,
            in3 => \N__36060\,
            lcout => \c0.data_in_field_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_851_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21580\,
            in2 => \_gnd_net_\,
            in3 => \N__22768\,
            lcout => \c0.n5225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i149_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__15993\,
            in1 => \N__36059\,
            in2 => \N__26808\,
            in3 => \N__36508\,
            lcout => \c0.data_in_frame_18_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_918_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15979\,
            in1 => \N__22078\,
            in2 => \N__17896\,
            in3 => \N__15925\,
            lcout => \c0.n5266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i104_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34074\,
            in1 => \N__24779\,
            in2 => \_gnd_net_\,
            in3 => \N__25725\,
            lcout => data_in_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_4_lut_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32990\,
            in1 => \N__29367\,
            in2 => \N__24757\,
            in3 => \N__22946\,
            lcout => OPEN,
            ltout => \c0.n18_adj_1882_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_866_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24709\,
            in1 => \N__15959\,
            in2 => \N__15928\,
            in3 => \N__25018\,
            lcout => \c0.n26_adj_1883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_120_2_lut_3_lut_4_lut_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22823\,
            in1 => \N__32985\,
            in2 => \N__32914\,
            in3 => \N__29366\,
            lcout => \c0.n6103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i87_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__29977\,
            in1 => \N__36011\,
            in2 => \N__32994\,
            in3 => \N__36638\,
            lcout => \c0.data_in_field_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_859_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21733\,
            in2 => \_gnd_net_\,
            in3 => \N__32986\,
            lcout => \c0.n5201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i31_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__21734\,
            in1 => \N__36637\,
            in2 => \N__27850\,
            in3 => \N__36012\,
            lcout => \c0.data_in_field_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i110_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34218\,
            in1 => \N__19440\,
            in2 => \_gnd_net_\,
            in3 => \N__17594\,
            lcout => data_in_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5731_bdd_4_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__21947\,
            in1 => \N__32791\,
            in2 => \N__17905\,
            in3 => \N__29800\,
            lcout => \c0.n5462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i102_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17595\,
            in1 => \N__34073\,
            in2 => \_gnd_net_\,
            in3 => \N__16029\,
            lcout => data_in_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i84_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__35991\,
            in1 => \N__37127\,
            in2 => \N__26473\,
            in3 => \N__23422\,
            lcout => \c0.data_in_field_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i106_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37126\,
            in1 => \N__35992\,
            in2 => \N__21954\,
            in3 => \N__30979\,
            lcout => \c0.data_in_field_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i121_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23468\,
            in1 => \N__19629\,
            in2 => \N__36196\,
            in3 => \N__37128\,
            lcout => \c0.data_in_field_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_986_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22161\,
            in1 => \N__21946\,
            in2 => \_gnd_net_\,
            in3 => \N__23467\,
            lcout => \c0.n5222\,
            ltout => \c0.n5222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_3_lut_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17506\,
            in2 => \N__16069\,
            in3 => \N__21882\,
            lcout => OPEN,
            ltout => \c0.n33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28333\,
            in1 => \N__16066\,
            in2 => \N__16060\,
            in3 => \N__25414\,
            lcout => \c0.n45_adj_1885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i96_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24789\,
            in1 => \N__34082\,
            in2 => \_gnd_net_\,
            in3 => \N__22721\,
            lcout => data_in_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i152_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__26039\,
            in1 => \N__20159\,
            in2 => \N__34284\,
            in3 => \_gnd_net_\,
            lcout => data_in_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_825_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20185\,
            in2 => \_gnd_net_\,
            in3 => \N__24841\,
            lcout => \c0.n2008\,
            ltout => \c0.n2008_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_867_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24635\,
            in1 => \N__23553\,
            in2 => \N__16057\,
            in3 => \N__22870\,
            lcout => OPEN,
            ltout => \c0.n38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24853\,
            in1 => \N__26038\,
            in2 => \N__16054\,
            in3 => \N__26264\,
            lcout => \c0.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i112_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34076\,
            in1 => \N__21663\,
            in2 => \_gnd_net_\,
            in3 => \N__25718\,
            lcout => data_in_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i121_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27613\,
            in1 => \N__34081\,
            in2 => \_gnd_net_\,
            in3 => \N__19614\,
            lcout => data_in_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i159_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34077\,
            in1 => \N__16084\,
            in2 => \_gnd_net_\,
            in3 => \N__17360\,
            lcout => data_in_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_124_2_lut_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28789\,
            in2 => \_gnd_net_\,
            in3 => \N__20042\,
            lcout => \c0.n6107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34035\,
            in1 => \N__16103\,
            in2 => \_gnd_net_\,
            in3 => \N__24146\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i151_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__16125\,
            in1 => \N__24212\,
            in2 => \N__36193\,
            in3 => \N__36639\,
            lcout => \c0.data_in_frame_18_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_949_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31730\,
            in1 => \N__16102\,
            in2 => \N__31440\,
            in3 => \N__17836\,
            lcout => \c0.n26_adj_1955\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i62_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34036\,
            in1 => \N__22497\,
            in2 => \_gnd_net_\,
            in3 => \N__24234\,
            lcout => data_in_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i157_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16156\,
            in1 => \N__34037\,
            in2 => \_gnd_net_\,
            in3 => \N__37315\,
            lcout => data_in_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__16080\,
            in1 => \N__20935\,
            in2 => \N__17953\,
            in3 => \N__20835\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i72_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23845\,
            in1 => \N__33874\,
            in2 => \_gnd_net_\,
            in3 => \N__22457\,
            lcout => data_in_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33872\,
            in1 => \N__22671\,
            in2 => \_gnd_net_\,
            in3 => \N__27577\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_4_lut_4_lut_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100100010001"
        )
    port map (
            in0 => \N__18136\,
            in1 => \N__18278\,
            in2 => \N__18364\,
            in3 => \N__18066\,
            lcout => OPEN,
            ltout => \c0.rx.n2151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__33873\,
            in1 => \N__18279\,
            in2 => \N__16177\,
            in3 => \N__18361\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_4_lut_adj_792_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__18179\,
            in1 => \N__18190\,
            in2 => \N__18139\,
            in3 => \N__18065\,
            lcout => n1709,
            ltout => \n1709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__20933\,
            in1 => \N__16155\,
            in2 => \N__16174\,
            in3 => \N__16171\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__18015\,
            in1 => \N__17948\,
            in2 => \N__21480\,
            in3 => \N__20934\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i8_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__16354\,
            in1 => \N__19207\,
            in2 => \N__18508\,
            in3 => \N__19078\,
            lcout => data_out_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_973_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20468\,
            in1 => \N__20748\,
            in2 => \N__18813\,
            in3 => \N__16582\,
            lcout => n4_adj_1992,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i972_2_lut_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21318\,
            in2 => \_gnd_net_\,
            in3 => \N__20586\,
            lcout => \c0.n1227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2006_4_lut_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__18976\,
            in1 => \N__21417\,
            in2 => \N__16514\,
            in3 => \N__20403\,
            lcout => \c0.n2249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i11_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__16512\,
            in1 => \N__19221\,
            in2 => \N__18448\,
            in3 => \N__19056\,
            lcout => data_out_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_971_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16809\,
            in1 => \N__16344\,
            in2 => \N__16515\,
            in3 => \N__16271\,
            lcout => n5135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i9_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__16272\,
            in1 => \N__19222\,
            in2 => \N__18490\,
            in3 => \N__19057\,
            lcout => data_out_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5249_4_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__16245\,
            in1 => \N__20678\,
            in2 => \N__16234\,
            in3 => \N__20404\,
            lcout => OPEN,
            ltout => \c0.n5522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__18657\,
            in1 => \N__16213\,
            in2 => \N__16207\,
            in3 => \N__21187\,
            lcout => \tx_data_2_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_845_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16363\,
            in2 => \_gnd_net_\,
            in3 => \N__16435\,
            lcout => n4_adj_1991,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5257_4_lut_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__16197\,
            in1 => \N__20677\,
            in2 => \N__16600\,
            in3 => \N__20413\,
            lcout => \c0.n5489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_940_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16703\,
            in1 => \N__18748\,
            in2 => \_gnd_net_\,
            in3 => \N__16580\,
            lcout => n4_adj_1994,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_941_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__18792\,
            in1 => \_gnd_net_\,
            in2 => \N__16710\,
            in3 => \N__16581\,
            lcout => n5117,
            ltout => \n5117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i30_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__16599\,
            in1 => \N__20692\,
            in2 => \N__16684\,
            in3 => \N__16681\,
            lcout => data_out_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19368\,
            in1 => \N__16588\,
            in2 => \_gnd_net_\,
            in3 => \N__17256\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_936_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18781\,
            in1 => \N__20744\,
            in2 => \_gnd_net_\,
            in3 => \N__16579\,
            lcout => \c0.n1805\,
            ltout => \c0.n1805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_965_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16519\,
            in1 => \N__20641\,
            in2 => \N__16477\,
            in3 => \N__16433\,
            lcout => n135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21119\,
            in1 => \N__20743\,
            in2 => \_gnd_net_\,
            in3 => \N__20410\,
            lcout => \c0.n9_adj_1890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_933_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16450\,
            in1 => \N__20642\,
            in2 => \_gnd_net_\,
            in3 => \N__16434\,
            lcout => n5173,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2004_4_lut_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__16432\,
            in1 => \N__21415\,
            in2 => \N__16370\,
            in3 => \N__20411\,
            lcout => \c0.n2247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i26_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110000"
        )
    port map (
            in0 => \N__19208\,
            in1 => \N__16318\,
            in2 => \N__16309\,
            in3 => \N__19079\,
            lcout => data_out_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__16849\,
            in1 => \N__16843\,
            in2 => \N__21238\,
            in3 => \N__21190\,
            lcout => \tx_data_3_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_5365_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__18639\,
            in1 => \N__19311\,
            in2 => \N__17242\,
            in3 => \N__17184\,
            lcout => OPEN,
            ltout => \c0.tx.n5713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n5713_bdd_4_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__17233\,
            in1 => \N__16831\,
            in2 => \N__16813\,
            in3 => \N__16728\,
            lcout => \c0.tx.n5716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16808\,
            in1 => \N__21044\,
            in2 => \_gnd_net_\,
            in3 => \N__20405\,
            lcout => \c0.n9_adj_1880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i750_4_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100100010"
        )
    port map (
            in0 => \N__20406\,
            in1 => \N__21416\,
            in2 => \N__16756\,
            in3 => \N__20587\,
            lcout => OPEN,
            ltout => \c0.n991_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__21191\,
            in1 => \N__16744\,
            in2 => \N__16735\,
            in3 => \N__21314\,
            lcout => OPEN,
            ltout => \tx_data_5_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19369\,
            in2 => \N__16732\,
            in3 => \N__16729\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i2_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__21059\,
            in1 => \N__19224\,
            in2 => \N__18601\,
            in3 => \N__19083\,
            lcout => data_out_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19370\,
            in1 => \N__16720\,
            in2 => \_gnd_net_\,
            in3 => \N__17266\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__17265\,
            in1 => \N__17257\,
            in2 => \N__17238\,
            in3 => \N__17183\,
            lcout => \c0.tx.n5719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i342127_i1_3_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17151\,
            in1 => \N__17134\,
            in2 => \_gnd_net_\,
            in3 => \N__17128\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_N_1798_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17117\,
            in2 => \N__17065\,
            in3 => \N__17061\,
            lcout => OPEN,
            ltout => \c0.tx.n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16992\,
            in1 => \_gnd_net_\,
            in2 => \N__16894\,
            in3 => \N__16869\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_811_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29030\,
            in2 => \_gnd_net_\,
            in3 => \N__25998\,
            lcout => \c0.n2018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_870_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19746\,
            in1 => \N__29534\,
            in2 => \N__16858\,
            in3 => \N__23757\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i147_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__17398\,
            in1 => \N__36496\,
            in2 => \N__31251\,
            in3 => \N__36321\,
            lcout => \c0.data_in_frame_18_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_857_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30381\,
            in2 => \_gnd_net_\,
            in3 => \N__30849\,
            lcout => \c0.n5147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i108_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__30382\,
            in1 => \N__36494\,
            in2 => \N__31870\,
            in3 => \N__36319\,
            lcout => \c0.data_in_field_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i130_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__30850\,
            in1 => \N__36495\,
            in2 => \N__30223\,
            in3 => \N__36320\,
            lcout => \c0.data_in_field_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5573_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__17397\,
            in1 => \N__32412\,
            in2 => \N__18889\,
            in3 => \N__33212\,
            lcout => \c0.n5965\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_885_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19378\,
            in1 => \N__28029\,
            in2 => \N__17371\,
            in3 => \N__28756\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1901_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_928_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19951\,
            in1 => \N__23179\,
            in2 => \N__17332\,
            in3 => \N__34684\,
            lcout => \c0.n5280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_931_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17635\,
            in1 => \N__17329\,
            in2 => \N__19549\,
            in3 => \N__17776\,
            lcout => OPEN,
            ltout => \c0.n30_adj_1940_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3321_4_lut_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35838\,
            in1 => \N__17290\,
            in2 => \N__17323\,
            in3 => \N__17446\,
            lcout => \c0.n3563\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_932_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__19690\,
            in1 => \N__17302\,
            in2 => \N__19402\,
            in3 => \N__17296\,
            lcout => \c0.n25_adj_1941\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_900_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23335\,
            in1 => \N__17284\,
            in2 => \N__17626\,
            in3 => \N__17695\,
            lcout => OPEN,
            ltout => \c0.n26_adj_1915_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_903_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19603\,
            in1 => \N__24484\,
            in2 => \N__17542\,
            in3 => \N__22441\,
            lcout => \c0.n5250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i140_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__17539\,
            in1 => \N__36314\,
            in2 => \N__25008\,
            in3 => \N__36509\,
            lcout => \c0.data_in_field_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19602\,
            in1 => \N__22522\,
            in2 => \_gnd_net_\,
            in3 => \N__17608\,
            lcout => OPEN,
            ltout => \c0.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_901_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30316\,
            in1 => \N__17507\,
            in2 => \N__17464\,
            in3 => \N__22315\,
            lcout => OPEN,
            ltout => \c0.n28_adj_1917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_930_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101101"
        )
    port map (
            in0 => \N__17461\,
            in1 => \N__17455\,
            in2 => \N__17449\,
            in3 => \N__19717\,
            lcout => \c0.n26_adj_1939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_886_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17440\,
            in1 => \N__31203\,
            in2 => \N__17877\,
            in3 => \N__25161\,
            lcout => \c0.n28_adj_1902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i127_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__23692\,
            in1 => \N__36315\,
            in2 => \N__33360\,
            in3 => \N__36951\,
            lcout => \c0.data_in_field_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i135_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__36950\,
            in1 => \N__19680\,
            in2 => \N__36330\,
            in3 => \N__17935\,
            lcout => \c0.data_in_field_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_873_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23492\,
            in1 => \N__19670\,
            in2 => \N__19584\,
            in3 => \N__33346\,
            lcout => OPEN,
            ltout => \c0.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24280\,
            in2 => \N__17401\,
            in3 => \N__23575\,
            lcout => OPEN,
            ltout => \c0.n16_adj_1893_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_920_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001111011"
        )
    port map (
            in0 => \N__17653\,
            in1 => \N__19891\,
            in2 => \N__17638\,
            in3 => \N__23161\,
            lcout => \c0.n22_adj_1930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_830_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29608\,
            in2 => \_gnd_net_\,
            in3 => \N__28025\,
            lcout => \c0.n2058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21735\,
            in1 => \N__17561\,
            in2 => \N__22623\,
            in3 => \N__26901\,
            lcout => \c0.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_858_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27296\,
            in2 => \_gnd_net_\,
            in3 => \N__23546\,
            lcout => OPEN,
            ltout => \c0.n5096_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_861_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19825\,
            in1 => \N__20284\,
            in2 => \N__17614\,
            in3 => \N__22023\,
            lcout => \c0.n1785\,
            ltout => \c0.n1785_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_862_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30673\,
            in1 => \N__28304\,
            in2 => \N__17611\,
            in3 => \N__25052\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i110_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36937\,
            in1 => \N__35996\,
            in2 => \N__17599\,
            in3 => \N__17562\,
            lcout => \c0.data_in_field_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_981_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19826\,
            lcout => \c0.n5150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_962_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19824\,
            in1 => \N__17559\,
            in2 => \_gnd_net_\,
            in3 => \N__25004\,
            lcout => \c0.n2033\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_896_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29739\,
            in1 => \N__24328\,
            in2 => \N__33476\,
            in3 => \N__17764\,
            lcout => \c0.n12_adj_1911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17815\,
            in1 => \N__17809\,
            in2 => \N__17803\,
            in3 => \N__17740\,
            lcout => OPEN,
            ltout => \c0.n5275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_919_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__17701\,
            in1 => \N__17791\,
            in2 => \N__17779\,
            in3 => \N__20227\,
            lcout => \c0.n24_adj_1929\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_998_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27657\,
            in1 => \N__27297\,
            in2 => \N__17733\,
            in3 => \N__19641\,
            lcout => \c0.n5182\,
            ltout => \c0.n5182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17758\,
            in1 => \N__31554\,
            in2 => \N__17743\,
            in3 => \N__23571\,
            lcout => \c0.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_872_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23928\,
            in1 => \N__30757\,
            in2 => \N__17734\,
            in3 => \N__26730\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26260\,
            in1 => \N__26111\,
            in2 => \_gnd_net_\,
            in3 => \N__19870\,
            lcout => \c0.n20_adj_1906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i36_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__35649\,
            in1 => \N__37132\,
            in2 => \N__19983\,
            in3 => \N__17685\,
            lcout => \c0.data_in_field_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i11_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__27466\,
            in1 => \N__35650\,
            in2 => \N__37229\,
            in3 => \N__22822\,
            lcout => \c0.data_in_field_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i135_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24183\,
            in1 => \N__34220\,
            in2 => \_gnd_net_\,
            in3 => \N__17921\,
            lcout => data_in_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5380_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33286\,
            in1 => \N__22571\,
            in2 => \N__32630\,
            in3 => \N__24085\,
            lcout => \c0.n5731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i134_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__20041\,
            in1 => \N__24475\,
            in2 => \N__37230\,
            in3 => \N__35651\,
            lcout => \c0.data_in_field_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_989_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20005\,
            in1 => \N__21711\,
            in2 => \N__28788\,
            in3 => \N__20040\,
            lcout => \c0.n5264\,
            ltout => \c0.n5264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_990_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20186\,
            in2 => \N__17881\,
            in3 => \N__22821\,
            lcout => \c0.n14_adj_1967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i154_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33884\,
            in1 => \N__17998\,
            in2 => \_gnd_net_\,
            in3 => \N__17866\,
            lcout => data_in_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i26_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__23788\,
            in1 => \N__35645\,
            in2 => \N__37231\,
            in3 => \N__20188\,
            lcout => \c0.data_in_field_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i146_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33883\,
            in1 => \N__20085\,
            in2 => \_gnd_net_\,
            in3 => \N__17867\,
            lcout => data_in_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33878\,
            in1 => \N__17844\,
            in2 => \_gnd_net_\,
            in3 => \N__22363\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i8_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__35644\,
            in1 => \N__17982\,
            in2 => \N__20115\,
            in3 => \N__37142\,
            lcout => \c0.data_in_field_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i126_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33877\,
            in1 => \N__24474\,
            in2 => \_gnd_net_\,
            in3 => \N__20207\,
            lcout => data_in_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_948_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23111\,
            in1 => \N__24139\,
            in2 => \N__27585\,
            in3 => \N__17981\,
            lcout => \c0.n28_adj_1954\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33879\,
            in1 => \N__23891\,
            in2 => \_gnd_net_\,
            in3 => \N__23112\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_798_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18357\,
            in2 => \_gnd_net_\,
            in3 => \N__18277\,
            lcout => \c0.rx.n5058\,
            ltout => \c0.rx.n5058_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_4_lut_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__18178\,
            in1 => \N__18132\,
            in2 => \N__18070\,
            in3 => \N__18067\,
            lcout => n1714,
            ltout => \n1714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__17994\,
            in1 => \N__18016\,
            in2 => \N__18001\,
            in3 => \N__20931\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33876\,
            in1 => \N__17983\,
            in2 => \_gnd_net_\,
            in3 => \N__27578\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__17968\,
            in1 => \N__17952\,
            in2 => \N__22416\,
            in3 => \N__20932\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i145_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33875\,
            in1 => \N__33454\,
            in2 => \_gnd_net_\,
            in3 => \N__21463\,
            lcout => data_in_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i0_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18486\,
            in2 => \_gnd_net_\,
            in3 => \N__18475\,
            lcout => data_0,
            ltout => OPEN,
            carryin => \bfn_6_17_0_\,
            carryout => \c0.n4385\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i1_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18462\,
            in2 => \_gnd_net_\,
            in3 => \N__18451\,
            lcout => data_1,
            ltout => OPEN,
            carryin => \c0.n4385\,
            carryout => \c0.n4386\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i2_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18441\,
            in2 => \_gnd_net_\,
            in3 => \N__18430\,
            lcout => data_2,
            ltout => OPEN,
            carryin => \c0.n4386\,
            carryout => \c0.n4387\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i3_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18423\,
            in2 => \_gnd_net_\,
            in3 => \N__18412\,
            lcout => data_3,
            ltout => OPEN,
            carryin => \c0.n4387\,
            carryout => \c0.n4388\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i4_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18843\,
            in2 => \_gnd_net_\,
            in3 => \N__18409\,
            lcout => data_4,
            ltout => OPEN,
            carryin => \c0.n4388\,
            carryout => \c0.n4389\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i5_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18396\,
            in2 => \_gnd_net_\,
            in3 => \N__18385\,
            lcout => data_5,
            ltout => OPEN,
            carryin => \c0.n4389\,
            carryout => \c0.n4390\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i6_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18378\,
            in2 => \_gnd_net_\,
            in3 => \N__18367\,
            lcout => data_6,
            ltout => OPEN,
            carryin => \c0.n4390\,
            carryout => \c0.n4391\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i7_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18618\,
            in2 => \_gnd_net_\,
            in3 => \N__18607\,
            lcout => data_7,
            ltout => OPEN,
            carryin => \c0.n4391\,
            carryout => \c0.n4392\,
            clk => \N__35282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i8_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18696\,
            in2 => \_gnd_net_\,
            in3 => \N__18604\,
            lcout => data_8,
            ltout => OPEN,
            carryin => \bfn_6_18_0_\,
            carryout => \c0.n4393\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i9_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18591\,
            in2 => \_gnd_net_\,
            in3 => \N__18580\,
            lcout => data_9,
            ltout => OPEN,
            carryin => \c0.n4393\,
            carryout => \c0.n4394\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i10_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19098\,
            in2 => \_gnd_net_\,
            in3 => \N__18577\,
            lcout => data_10,
            ltout => OPEN,
            carryin => \c0.n4394\,
            carryout => \c0.n4395\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i11_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18567\,
            in2 => \_gnd_net_\,
            in3 => \N__18556\,
            lcout => data_11,
            ltout => OPEN,
            carryin => \c0.n4395\,
            carryout => \c0.n4396\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i12_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18549\,
            in2 => \_gnd_net_\,
            in3 => \N__18538\,
            lcout => data_12,
            ltout => OPEN,
            carryin => \c0.n4396\,
            carryout => \c0.n4397\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i13_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18528\,
            in2 => \_gnd_net_\,
            in3 => \N__18517\,
            lcout => data_13,
            ltout => OPEN,
            carryin => \c0.n4397\,
            carryout => \c0.n4398\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i14_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18828\,
            in2 => \_gnd_net_\,
            in3 => \N__18514\,
            lcout => data_14,
            ltout => OPEN,
            carryin => \c0.n4398\,
            carryout => \c0.n4399\,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i15_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \_gnd_net_\,
            in3 => \N__18511\,
            lcout => data_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i13_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__18780\,
            in1 => \N__19209\,
            in2 => \N__18850\,
            in3 => \N__19080\,
            lcout => data_out_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i7_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__19082\,
            in1 => \N__20459\,
            in2 => \N__18832\,
            in3 => \N__19213\,
            lcout => data_out_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18779\,
            in1 => \N__18750\,
            in2 => \_gnd_net_\,
            in3 => \N__20415\,
            lcout => OPEN,
            ltout => \c0.n9_adj_1887_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i15_3_lut_3_lut_4_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100001110111"
        )
    port map (
            in0 => \N__21414\,
            in1 => \N__21321\,
            in2 => \N__18709\,
            in3 => \N__20584\,
            lcout => \c0.n15_adj_1889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i1_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__19282\,
            in1 => \N__18697\,
            in2 => \N__19223\,
            in3 => \N__19081\,
            lcout => data_out_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i980_2_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21413\,
            in2 => \_gnd_net_\,
            in3 => \N__21320\,
            lcout => \c0.n1236\,
            ltout => \c0.n1236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5231_3_lut_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__18685\,
            in1 => \_gnd_net_\,
            in2 => \N__18673\,
            in3 => \N__20585\,
            lcout => OPEN,
            ltout => \c0.n5511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111011"
        )
    port map (
            in0 => \N__18670\,
            in1 => \N__18664\,
            in2 => \N__18646\,
            in3 => \N__21196\,
            lcout => OPEN,
            ltout => \tx_data_7_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19372\,
            in1 => \_gnd_net_\,
            in2 => \N__18643\,
            in3 => \N__18640\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19371\,
            in1 => \N__21130\,
            in2 => \_gnd_net_\,
            in3 => \N__19312\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_833_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18954\,
            lcout => n1748,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i3_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__18955\,
            in1 => \N__19225\,
            in2 => \N__19105\,
            in3 => \N__19087\,
            lcout => data_out_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5827_bdd_4_lut_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__34820\,
            in1 => \N__18928\,
            in2 => \N__24595\,
            in3 => \N__20941\,
            lcout => \c0.n5830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5558_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18870\,
            in1 => \N__32483\,
            in2 => \N__18862\,
            in3 => \N__33186\,
            lcout => \c0.n5941\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i155_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__35857\,
            in1 => \N__18888\,
            in2 => \N__24442\,
            in3 => \N__36607\,
            lcout => \c0.data_in_frame_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i150_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__36605\,
            in1 => \N__21523\,
            in2 => \N__18874\,
            in3 => \N__35861\,
            lcout => \c0.data_in_frame_18_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i158_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__35858\,
            in1 => \N__18861\,
            in2 => \N__24529\,
            in3 => \N__36608\,
            lcout => \c0.data_in_frame_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i118_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36604\,
            in1 => \N__35859\,
            in2 => \N__19447\,
            in3 => \N__23047\,
            lcout => \c0.data_in_field_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19793\,
            in1 => \N__21517\,
            in2 => \N__23054\,
            in3 => \N__23256\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i55_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36606\,
            in1 => \N__35860\,
            in2 => \N__26218\,
            in3 => \N__22864\,
            lcout => \c0.data_in_field_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5445_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33185\,
            in1 => \N__22160\,
            in2 => \N__32572\,
            in3 => \N__20272\,
            lcout => \c0.n5809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i98_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34286\,
            in1 => \N__30975\,
            in2 => \_gnd_net_\,
            in3 => \N__25331\,
            lcout => data_in_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_927_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28305\,
            in1 => \N__19567\,
            in2 => \N__34636\,
            in3 => \N__21637\,
            lcout => \c0.n5241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_field_143__I_0_1808_2_lut_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27137\,
            in2 => \_gnd_net_\,
            in3 => \N__25678\,
            lcout => \c0.tx2_transmit_N_1031\,
            ltout => \c0.tx2_transmit_N_1031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21496\,
            in1 => \N__21826\,
            in2 => \N__19390\,
            in3 => \N__21901\,
            lcout => \c0.n38_adj_1934\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34285\,
            in1 => \N__26155\,
            in2 => \_gnd_net_\,
            in3 => \N__22265\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_979_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29140\,
            in1 => \N__24675\,
            in2 => \N__29218\,
            in3 => \N__27426\,
            lcout => \c0.n14_adj_1900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i150_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24528\,
            in1 => \N__34287\,
            in2 => \_gnd_net_\,
            in3 => \N__21521\,
            lcout => data_in_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i113_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34460\,
            in1 => \N__19630\,
            in2 => \_gnd_net_\,
            in3 => \N__24351\,
            lcout => data_in_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_855_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20013\,
            in2 => \_gnd_net_\,
            in3 => \N__29139\,
            lcout => \c0.n5210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_883_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30664\,
            in1 => \N__19591\,
            in2 => \N__37338\,
            in3 => \N__19585\,
            lcout => \c0.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_914_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26416\,
            in1 => \N__30481\,
            in2 => \N__31030\,
            in3 => \N__19453\,
            lcout => OPEN,
            ltout => \c0.n5259_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_922_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111001"
        )
    port map (
            in0 => \N__23449\,
            in1 => \N__19561\,
            in2 => \N__19552\,
            in3 => \N__21781\,
            lcout => \c0.n21_adj_1933\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_895_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19540\,
            in1 => \N__21811\,
            in2 => \N__19531\,
            in3 => \N__19507\,
            lcout => \c0.n18_adj_1910\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_850_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21918\,
            lcout => \c0.n5198\,
            ltout => \c0.n5198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19486\,
            in1 => \N__23211\,
            in2 => \N__19477\,
            in3 => \N__19474\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_888_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21810\,
            in1 => \N__21598\,
            in2 => \N__24279\,
            in3 => \N__26629\,
            lcout => \c0.n31_adj_1904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_897_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19762\,
            in1 => \N__19885\,
            in2 => \N__19756\,
            in3 => \N__27391\,
            lcout => OPEN,
            ltout => \c0.n17_adj_1912_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_905_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__27064\,
            in1 => \N__19732\,
            in2 => \N__19726\,
            in3 => \N__19723\,
            lcout => \c0.n19_adj_1920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_4_lut_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19905\,
            in1 => \N__22033\,
            in2 => \N__24960\,
            in3 => \N__19711\,
            lcout => \c0.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_889_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30404\,
            in1 => \N__25315\,
            in2 => \N__23437\,
            in3 => \N__19642\,
            lcout => OPEN,
            ltout => \c0.n29_adj_1905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_929_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19861\,
            in1 => \N__19705\,
            in2 => \N__19699\,
            in3 => \N__19696\,
            lcout => \c0.n5278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19668\,
            in1 => \N__33339\,
            in2 => \_gnd_net_\,
            in3 => \N__26295\,
            lcout => OPEN,
            ltout => \c0.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22778\,
            in1 => \N__29885\,
            in2 => \N__19645\,
            in3 => \N__23080\,
            lcout => \c0.n1880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_876_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22437\,
            in1 => \N__20163\,
            in2 => \N__19909\,
            in3 => \N__22102\,
            lcout => \c0.n20_adj_1892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_983_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30865\,
            in1 => \N__19884\,
            in2 => \N__28924\,
            in3 => \N__25957\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1963_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_960_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25676\,
            in1 => \N__29031\,
            in2 => \N__19873\,
            in3 => \N__26004\,
            lcout => \c0.n5114\,
            ltout => \c0.n5114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_887_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28351\,
            in1 => \N__21894\,
            in2 => \N__19864\,
            in3 => \N__25396\,
            lcout => \c0.n30_adj_1903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i91_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36038\,
            in1 => \N__37089\,
            in2 => \N__27310\,
            in3 => \N__31672\,
            lcout => \c0.data_in_field_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5390_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__26005\,
            in1 => \N__33289\,
            in2 => \N__32789\,
            in3 => \N__19791\,
            lcout => \c0.n5743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i88_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36037\,
            in1 => \N__37088\,
            in2 => \N__22705\,
            in3 => \N__19830\,
            lcout => \c0.data_in_field_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i58_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37087\,
            in1 => \N__36039\,
            in2 => \N__23986\,
            in3 => \N__19792\,
            lcout => \c0.data_in_field_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1000_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21976\,
            in1 => \N__19969\,
            in2 => \N__32950\,
            in3 => \N__22995\,
            lcout => \c0.n5162\,
            ltout => \c0.n5162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_819_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20105\,
            in2 => \N__20089\,
            in3 => \N__25250\,
            lcout => \c0.n1825\,
            ltout => \c0.n1825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_869_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20071\,
            in1 => \N__26380\,
            in2 => \N__20053\,
            in3 => \N__20043\,
            lcout => \c0.n28_adj_1886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i95_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__32938\,
            in1 => \N__36992\,
            in2 => \N__31288\,
            in3 => \N__35653\,
            lcout => \c0.data_in_field_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i96_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36990\,
            in1 => \N__35643\,
            in2 => \N__22735\,
            in3 => \N__22997\,
            lcout => \c0.data_in_field_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i74_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__35641\,
            in1 => \N__36991\,
            in2 => \N__26554\,
            in3 => \N__20012\,
            lcout => \c0.data_in_field_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i23_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__27891\,
            in1 => \N__35642\,
            in2 => \N__37161\,
            in3 => \N__22238\,
            lcout => \c0.data_in_field_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22996\,
            in1 => \N__25084\,
            in2 => \N__19979\,
            in3 => \N__31555\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i80_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23828\,
            in1 => \_gnd_net_\,
            in2 => \N__34296\,
            in3 => \N__22695\,
            lcout => data_in_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i138_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__20812\,
            in1 => \N__37285\,
            in2 => \N__35837\,
            in3 => \N__19923\,
            lcout => \c0.data_in_field_137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_829_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19922\,
            in1 => \N__20263\,
            in2 => \_gnd_net_\,
            in3 => \N__22303\,
            lcout => \c0.n2043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_860_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25143\,
            lcout => \c0.n6_adj_1877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i32_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__35768\,
            in1 => \N__24052\,
            in2 => \N__37290\,
            in3 => \N__20265\,
            lcout => \c0.data_in_field_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_871_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22389\,
            in1 => \N__20248\,
            in2 => \N__20242\,
            in3 => \N__22504\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_956_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__23275\,
            in1 => \N__27811\,
            in2 => \N__22639\,
            in3 => \N__22321\,
            lcout => \c0.n1686\,
            ltout => \c0.n1686_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i126_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__20217\,
            in1 => \N__37281\,
            in2 => \N__20191\,
            in3 => \N__28810\,
            lcout => \c0.data_in_field_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5400_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33309\,
            in1 => \N__20187\,
            in2 => \N__32735\,
            in3 => \N__22307\,
            lcout => \c0.n5749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34010\,
            in1 => \N__24048\,
            in2 => \_gnd_net_\,
            in3 => \N__22670\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i114_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37201\,
            in1 => \N__35640\,
            in2 => \N__31012\,
            in3 => \N__22567\,
            lcout => \c0.data_in_field_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i160_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34009\,
            in1 => \N__20820\,
            in2 => \_gnd_net_\,
            in3 => \N__20149\,
            lcout => data_in_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__20916\,
            in1 => \N__20850\,
            in2 => \N__20824\,
            in3 => \N__20839\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i130_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20811\,
            in1 => \N__34011\,
            in2 => \_gnd_net_\,
            in3 => \N__30203\,
            lcout => data_in_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i136_LC_6_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__35639\,
            in1 => \N__37202\,
            in2 => \N__25618\,
            in3 => \N__22603\,
            lcout => \c0.data_in_field_135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3325_2_lut_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20530\,
            in2 => \_gnd_net_\,
            in3 => \N__20355\,
            lcout => \c0.n3567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5247_4_lut_4_lut_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111110101"
        )
    port map (
            in0 => \N__20582\,
            in1 => \N__20785\,
            in2 => \N__20770\,
            in3 => \N__20416\,
            lcout => \c0.n5515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_892_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20647\,
            in2 => \_gnd_net_\,
            in3 => \N__20749\,
            lcout => n5176,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_972_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21412\,
            in1 => \N__21319\,
            in2 => \_gnd_net_\,
            in3 => \N__20581\,
            lcout => \c0.n1590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5259_4_lut_4_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__20643\,
            in1 => \N__20583\,
            in2 => \N__20469\,
            in3 => \N__20414\,
            lcout => OPEN,
            ltout => \c0.n5523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5256_4_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010001"
        )
    port map (
            in0 => \N__21427\,
            in1 => \N__21418\,
            in2 => \N__21325\,
            in3 => \N__21322\,
            lcout => OPEN,
            ltout => \c0.n5513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__21231\,
            in1 => \N__21205\,
            in2 => \N__21199\,
            in3 => \N__21195\,
            lcout => \tx_data_6_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_980_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21124\,
            in1 => \N__21078\,
            in2 => \_gnd_net_\,
            in3 => \N__21016\,
            lcout => n5132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5470_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33275\,
            in1 => \N__30546\,
            in2 => \N__32777\,
            in3 => \N__27016\,
            lcout => OPEN,
            ltout => \c0.n5839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5839_bdd_4_lut_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32775\,
            in1 => \N__26379\,
            in2 => \N__20956\,
            in3 => \N__29686\,
            lcout => \c0.n5414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5465_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33276\,
            in1 => \N__31114\,
            in2 => \N__32778\,
            in3 => \N__25117\,
            lcout => OPEN,
            ltout => \c0.n5833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5833_bdd_4_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32776\,
            in1 => \N__27187\,
            in2 => \N__20953\,
            in3 => \N__28669\,
            lcout => OPEN,
            ltout => \c0.n5417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5480_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__34813\,
            in1 => \N__32122\,
            in2 => \N__20950\,
            in3 => \N__20947\,
            lcout => \c0.n5827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5351_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33201\,
            in1 => \N__29889\,
            in2 => \N__32582\,
            in3 => \N__25162\,
            lcout => \c0.n5695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5341_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__23500\,
            in1 => \N__33202\,
            in2 => \N__24327\,
            in3 => \N__32502\,
            lcout => OPEN,
            ltout => \c0.n5683_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5683_bdd_4_lut_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32503\,
            in1 => \N__22950\,
            in2 => \N__21553\,
            in3 => \N__23149\,
            lcout => \c0.n5483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5695_bdd_4_lut_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__21550\,
            in1 => \N__29032\,
            in2 => \N__29467\,
            in3 => \N__32504\,
            lcout => OPEN,
            ltout => \c0.n5480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5370_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__34804\,
            in1 => \N__32123\,
            in2 => \N__21544\,
            in3 => \N__21541\,
            lcout => OPEN,
            ltout => \c0.n5677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5677_bdd_4_lut_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__34812\,
            in1 => \N__24865\,
            in2 => \N__21535\,
            in3 => \N__28207\,
            lcout => \c0.n5680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i90_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34543\,
            in1 => \N__25332\,
            in2 => \_gnd_net_\,
            in3 => \N__28589\,
            lcout => data_in_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i142_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34367\,
            in1 => \N__24003\,
            in2 => \_gnd_net_\,
            in3 => \N__21522\,
            lcout => data_in_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21445\,
            in2 => \_gnd_net_\,
            in3 => \N__25056\,
            lcout => \c0.n24_adj_1895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i153_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21446\,
            in1 => \_gnd_net_\,
            in2 => \N__34505\,
            in3 => \N__21490\,
            lcout => data_in_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5797_bdd_4_lut_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__23392\,
            in1 => \N__24898\,
            in2 => \N__23260\,
            in3 => \N__32454\,
            lcout => \c0.n5429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5791_bdd_4_lut_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000010"
        )
    port map (
            in0 => \N__21592\,
            in1 => \N__21763\,
            in2 => \N__32571\,
            in3 => \N__30405\,
            lcout => \c0.n5432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5530_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33285\,
            in1 => \N__21742\,
            in2 => \N__32546\,
            in3 => \N__22246\,
            lcout => \c0.n5911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5881_bdd_4_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32476\,
            in1 => \N__21715\,
            in2 => \N__23707\,
            in3 => \N__25534\,
            lcout => \c0.n5393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i120_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34378\,
            in1 => \N__27688\,
            in2 => \_gnd_net_\,
            in3 => \N__21648\,
            lcout => data_in_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_882_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27085\,
            in1 => \N__26112\,
            in2 => \N__26272\,
            in3 => \N__26905\,
            lcout => \c0.n10_adj_1898\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i70_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__21617\,
            in1 => \N__36691\,
            in2 => \N__22498\,
            in3 => \N__36201\,
            lcout => \c0.data_in_field_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_997_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21616\,
            in2 => \_gnd_net_\,
            in3 => \N__22865\,
            lcout => \c0.n5159\,
            ltout => \c0.n5159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1001_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26365\,
            in1 => \N__21588\,
            in2 => \N__21556\,
            in3 => \N__22785\,
            lcout => \c0.n1978\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_827_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21955\,
            in2 => \_gnd_net_\,
            in3 => \N__23491\,
            lcout => OPEN,
            ltout => \c0.n2095_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_880_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22089\,
            in1 => \N__22897\,
            in2 => \N__21925\,
            in3 => \N__21922\,
            lcout => \c0.n34_adj_1896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5460_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__21837\,
            in2 => \N__32790\,
            in3 => \N__23380\,
            lcout => OPEN,
            ltout => \c0.n5821_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5821_bdd_4_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32755\,
            in1 => \N__21895\,
            in2 => \N__21856\,
            in3 => \N__31714\,
            lcout => \c0.n5423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i28_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__36227\,
            in1 => \N__21838\,
            in2 => \N__23323\,
            in3 => \N__36785\,
            lcout => \c0.data_in_field_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i13_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__24617\,
            in1 => \N__22272\,
            in2 => \N__36999\,
            in3 => \N__36228\,
            lcout => \c0.data_in_field_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_977_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21836\,
            in2 => \_gnd_net_\,
            in3 => \N__24616\,
            lcout => \c0.n2080\,
            ltout => \c0.n2080_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_978_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26375\,
            in1 => \N__26325\,
            in2 => \N__21814\,
            in3 => \N__32830\,
            lcout => \c0.n5243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_915_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30826\,
            in1 => \N__28326\,
            in2 => \N__21802\,
            in3 => \N__22077\,
            lcout => \c0.n25_adj_1926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_969_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24340\,
            in2 => \_gnd_net_\,
            in3 => \N__22090\,
            lcout => \c0.n5261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5346_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__33294\,
            in1 => \N__22193\,
            in2 => \N__26740\,
            in3 => \N__32785\,
            lcout => OPEN,
            ltout => \c0.n5689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5689_bdd_4_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32756\,
            in1 => \N__27721\,
            in2 => \N__22063\,
            in3 => \N__25564\,
            lcout => \c0.n5366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i56_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36017\,
            in1 => \N__36881\,
            in2 => \N__23812\,
            in3 => \N__22194\,
            lcout => \c0.data_in_field_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i133_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36880\,
            in1 => \N__36018\,
            in2 => \N__28195\,
            in3 => \N__27424\,
            lcout => \c0.data_in_field_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_993_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22045\,
            in1 => \N__29422\,
            in2 => \N__29743\,
            in3 => \N__22171\,
            lcout => \c0.n5276\,
            ltout => \c0.n5276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_924_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22027\,
            in1 => \N__27262\,
            in2 => \N__22012\,
            in3 => \N__25938\,
            lcout => \c0.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i37_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36030\,
            in1 => \N__37070\,
            in2 => \N__21992\,
            in3 => \N__30073\,
            lcout => \c0.data_in_field_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i86_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37069\,
            in1 => \N__36032\,
            in2 => \N__27550\,
            in3 => \N__23600\,
            lcout => \c0.data_in_field_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_818_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__24661\,
            in1 => \N__27414\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n2005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_820_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22231\,
            in1 => \N__31048\,
            in2 => \N__22210\,
            in3 => \N__23239\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1873_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_821_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__28250\,
            in1 => \_gnd_net_\,
            in2 => \N__22207\,
            in3 => \N__22204\,
            lcout => \c0.n5111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i53_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37068\,
            in1 => \N__36031\,
            in2 => \N__30037\,
            in3 => \N__31049\,
            lcout => \c0.data_in_field_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25410\,
            in1 => \N__22189\,
            in2 => \_gnd_net_\,
            in3 => \N__22141\,
            lcout => \c0.n13_adj_1951\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i21_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__24668\,
            in1 => \N__26154\,
            in2 => \N__37200\,
            in3 => \N__36033\,
            lcout => \c0.data_in_field_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i24_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__35646\,
            in1 => \N__22145\,
            in2 => \N__22678\,
            in3 => \N__36998\,
            lcout => \c0.data_in_field_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i54_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__24246\,
            in2 => \_gnd_net_\,
            in3 => \N__28100\,
            lcout => data_in_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_875_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23921\,
            in1 => \N__33403\,
            in2 => \N__22117\,
            in3 => \N__33359\,
            lcout => \c0.n18_adj_1891\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_945_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22534\,
            in1 => \N__26946\,
            in2 => \_gnd_net_\,
            in3 => \N__25493\,
            lcout => \c0.n5249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i68_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__35647\,
            in1 => \N__36996\,
            in2 => \N__33535\,
            in3 => \N__23248\,
            lcout => \c0.data_in_field_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i155_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34166\,
            in1 => \N__22423\,
            in2 => \_gnd_net_\,
            in3 => \N__24416\,
            lcout => data_in_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i89_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__35648\,
            in1 => \N__36997\,
            in2 => \N__28543\,
            in3 => \N__25150\,
            lcout => \c0.data_in_field_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_946_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25668\,
            in1 => \N__26945\,
            in2 => \_gnd_net_\,
            in3 => \N__25492\,
            lcout => \c0.n5255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_951_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22364\,
            in1 => \N__29239\,
            in2 => \N__22282\,
            in3 => \N__31416\,
            lcout => OPEN,
            ltout => \c0.n25_adj_1957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_954_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22342\,
            in1 => \N__22333\,
            in2 => \N__22324\,
            in3 => \N__22645\,
            lcout => \c0.n4465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i18_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__30187\,
            in1 => \N__35652\,
            in2 => \N__37291\,
            in3 => \N__22308\,
            lcout => \c0.data_in_field_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34168\,
            in1 => \N__22281\,
            in2 => \_gnd_net_\,
            in3 => \N__26394\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_854_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27012\,
            in1 => \N__25452\,
            in2 => \_gnd_net_\,
            in3 => \N__31786\,
            lcout => \c0.n1772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i88_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22734\,
            in1 => \_gnd_net_\,
            in2 => \N__34379\,
            in3 => \N__22694\,
            lcout => data_in_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_950_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30153\,
            in1 => \N__26393\,
            in2 => \N__29656\,
            in3 => \N__22663\,
            lcout => \c0.n27_adj_1956\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34012\,
            in1 => \N__29412\,
            in2 => \_gnd_net_\,
            in3 => \N__29246\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_952_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24047\,
            in1 => \N__23892\,
            in2 => \N__25912\,
            in3 => \N__23773\,
            lcout => \c0.n26_adj_1958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_856_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27650\,
            in1 => \N__22597\,
            in2 => \N__22572\,
            in3 => \N__22533\,
            lcout => \c0.n5144\,
            ltout => \c0.n5144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23215\,
            in1 => \N__25201\,
            in2 => \N__22507\,
            in3 => \N__22954\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i70_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34015\,
            in1 => \N__27517\,
            in2 => \_gnd_net_\,
            in3 => \N__22484\,
            lcout => data_in_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i64_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34013\,
            in1 => \N__22464\,
            in2 => \_gnd_net_\,
            in3 => \N__24101\,
            lcout => data_in_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_7_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34014\,
            in1 => \N__29335\,
            in2 => \_gnd_net_\,
            in3 => \N__23774\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5761_bdd_4_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__25770\,
            in1 => \N__22741\,
            in2 => \N__32698\,
            in3 => \N__24840\,
            lcout => OPEN,
            ltout => \c0.n5447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5420_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__34828\,
            in1 => \N__32124\,
            in2 => \N__22888\,
            in3 => \N__22747\,
            lcout => OPEN,
            ltout => \c0.n5755_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5755_bdd_4_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__34829\,
            in1 => \N__28219\,
            in2 => \N__22885\,
            in3 => \N__22795\,
            lcout => \c0.n5758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5525_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__33184\,
            in1 => \N__22869\,
            in2 => \N__26671\,
            in3 => \N__32667\,
            lcout => \c0.n5905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5779_bdd_4_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__27226\,
            in1 => \N__32674\,
            in2 => \N__24394\,
            in3 => \N__22834\,
            lcout => \c0.n5438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5410_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33182\,
            in1 => \N__22789\,
            in2 => \N__32697\,
            in3 => \N__27319\,
            lcout => OPEN,
            ltout => \c0.n5767_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5767_bdd_4_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32505\,
            in1 => \N__31204\,
            in2 => \N__22750\,
            in3 => \N__30580\,
            lcout => \c0.n5444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5405_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33183\,
            in1 => \N__30668\,
            in2 => \N__32696\,
            in3 => \N__31953\,
            lcout => \c0.n5761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i55_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34466\,
            in1 => \N__26523\,
            in2 => \_gnd_net_\,
            in3 => \N__26195\,
            lcout => data_in_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i97_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36953\,
            in1 => \N__35862\,
            in2 => \N__23098\,
            in3 => \N__22925\,
            lcout => \c0.data_in_field_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28456\,
            in1 => \N__23138\,
            in2 => \N__22936\,
            in3 => \N__30572\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i85_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27054\,
            in1 => \N__34467\,
            in2 => \_gnd_net_\,
            in3 => \N__26489\,
            lcout => data_in_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_957_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23539\,
            in1 => \N__29294\,
            in2 => \N__27318\,
            in3 => \N__28257\,
            lcout => \c0.n2074\,
            ltout => \c0.n2074_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_996_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23067\,
            in1 => \N__25533\,
            in2 => \N__23026\,
            in3 => \N__25292\,
            lcout => \c0.n5213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_970_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25251\,
            in1 => \N__29799\,
            in2 => \N__22971\,
            in3 => \N__32964\,
            lcout => \c0.n10_adj_1888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_848_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25560\,
            in1 => \N__22926\,
            in2 => \_gnd_net_\,
            in3 => \N__23008\,
            lcout => \c0.n1851\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_966_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22927\,
            in1 => \N__28457\,
            in2 => \N__24740\,
            in3 => \N__24970\,
            lcout => \c0.n5099\,
            ltout => \c0.n5099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_877_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23191\,
            in1 => \N__23175\,
            in2 => \N__23164\,
            in3 => \N__30260\,
            lcout => \c0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i105_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36194\,
            in1 => \N__37222\,
            in2 => \N__23148\,
            in3 => \N__24382\,
            lcout => \c0.data_in_field_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i7_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__28458\,
            in1 => \N__23122\,
            in2 => \N__37272\,
            in3 => \N__36195\,
            lcout => \c0.data_in_field_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i97_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34464\,
            in1 => \N__24381\,
            in2 => \_gnd_net_\,
            in3 => \N__23093\,
            lcout => data_in_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i89_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23094\,
            in1 => \N__34465\,
            in2 => \_gnd_net_\,
            in3 => \N__28523\,
            lcout => data_in_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i65_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36814\,
            in1 => \N__36226\,
            in2 => \N__27772\,
            in3 => \N__29015\,
            lcout => \c0.data_in_field_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i41_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28046\,
            in1 => \N__34474\,
            in2 => \_gnd_net_\,
            in3 => \N__26861\,
            lcout => data_in_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i57_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27768\,
            in1 => \_gnd_net_\,
            in2 => \N__34546\,
            in3 => \N__30929\,
            lcout => data_in_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i49_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__30930\,
            in1 => \_gnd_net_\,
            in2 => \N__28050\,
            in3 => \N__34478\,
            lcout => data_in_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i107_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34473\,
            in1 => \N__29078\,
            in2 => \_gnd_net_\,
            in3 => \N__30699\,
            lcout => data_in_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i90_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36225\,
            in1 => \N__36815\,
            in2 => \N__28609\,
            in3 => \N__23535\,
            lcout => \c0.data_in_field_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_912_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25763\,
            in1 => \N__27130\,
            in2 => \N__30672\,
            in3 => \N__23499\,
            lcout => \c0.n23_adj_1925\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5435_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33263\,
            in1 => \N__23436\,
            in2 => \N__32678\,
            in3 => \N__31785\,
            lcout => \c0.n5797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_890_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23379\,
            in1 => \N__31710\,
            in2 => \N__25080\,
            in3 => \N__24894\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_955_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26150\,
            in1 => \N__23319\,
            in2 => \N__29399\,
            in3 => \N__27353\,
            lcout => \c0.n25_adj_1960\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29398\,
            in1 => \N__34532\,
            in2 => \_gnd_net_\,
            in3 => \N__30615\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34531\,
            in1 => \N__31417\,
            in2 => \_gnd_net_\,
            in3 => \N__27354\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_852_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25367\,
            in1 => \N__29790\,
            in2 => \N__24836\,
            in3 => \N__23255\,
            lcout => \c0.n5093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i59_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__36197\,
            in1 => \N__30001\,
            in2 => \N__37079\,
            in3 => \N__28294\,
            lcout => \c0.data_in_field_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i58_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34533\,
            in1 => \N__30297\,
            in2 => \_gnd_net_\,
            in3 => \N__23972\,
            lcout => data_in_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5510_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33298\,
            in1 => \N__23652\,
            in2 => \N__32666\,
            in3 => \N__23758\,
            lcout => \c0.n5881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i30_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36034\,
            in1 => \N__36955\,
            in2 => \N__23656\,
            in3 => \N__27966\,
            lcout => \c0.data_in_field_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i143_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36954\,
            in1 => \N__36036\,
            in2 => \N__24184\,
            in3 => \N__27113\,
            lcout => \c0.data_in_field_142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i6_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36035\,
            in1 => \N__36956\,
            in2 => \N__27493\,
            in3 => \N__25526\,
            lcout => \c0.data_in_field_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i119_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34319\,
            in1 => \N__23691\,
            in2 => \_gnd_net_\,
            in3 => \N__28725\,
            lcout => data_in_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_988_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25652\,
            in1 => \N__23651\,
            in2 => \N__27126\,
            in3 => \N__23911\,
            lcout => \c0.n2046\,
            ltout => \c0.n2046_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_824_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23619\,
            in1 => \N__27370\,
            in2 => \N__23578\,
            in3 => \N__25392\,
            lcout => \c0.n5108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i50_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37148\,
            in1 => \N__35990\,
            in2 => \N__25997\,
            in3 => \N__23949\,
            lcout => \c0.data_in_field_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i50_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__34497\,
            in2 => \_gnd_net_\,
            in3 => \N__23979\,
            lcout => data_in_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i142_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37147\,
            in1 => \N__35989\,
            in2 => \N__24019\,
            in3 => \N__23920\,
            lcout => \c0.data_in_field_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i15_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__35986\,
            in1 => \N__23893\,
            in2 => \N__28509\,
            in3 => \N__37151\,
            lcout => \c0.data_in_field_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i48_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34495\,
            in1 => \N__27737\,
            in2 => \_gnd_net_\,
            in3 => \N__23802\,
            lcout => data_in_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i80_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__35988\,
            in1 => \N__37150\,
            in2 => \N__25497\,
            in3 => \N__23844\,
            lcout => \c0.data_in_field_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i56_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34496\,
            in1 => \N__24114\,
            in2 => \_gnd_net_\,
            in3 => \N__23801\,
            lcout => data_in_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i38_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__35987\,
            in1 => \N__37149\,
            in2 => \N__27802\,
            in3 => \N__25249\,
            lcout => \c0.data_in_field_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34493\,
            in1 => \N__30181\,
            in2 => \_gnd_net_\,
            in3 => \N__23787\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i122_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37143\,
            in1 => \N__36025\,
            in2 => \N__31168\,
            in3 => \N__24068\,
            lcout => \c0.data_in_field_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i62_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36024\,
            in1 => \N__37146\,
            in2 => \N__25294\,
            in3 => \N__24250\,
            lcout => \c0.data_in_field_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i143_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34320\,
            in1 => \N__24170\,
            in2 => \_gnd_net_\,
            in3 => \N__24222\,
            lcout => data_in_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34494\,
            in1 => \N__24150\,
            in2 => \_gnd_net_\,
            in3 => \N__27488\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i64_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37144\,
            in1 => \N__36026\,
            in2 => \N__24118\,
            in3 => \N__26715\,
            lcout => \c0.data_in_field_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i2_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__25836\,
            in1 => \N__37145\,
            in2 => \N__36204\,
            in3 => \N__29655\,
            lcout => \c0.data_in_field_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_822_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25282\,
            in1 => \N__24067\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \c0.n1830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i40_LC_9_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34140\,
            in1 => \N__27744\,
            in2 => \_gnd_net_\,
            in3 => \N__25577\,
            lcout => data_in_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_9_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25578\,
            in1 => \N__34141\,
            in2 => \_gnd_net_\,
            in3 => \N__24043\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i33_LC_9_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34139\,
            in1 => \N__26874\,
            in2 => \_gnd_net_\,
            in3 => \N__29151\,
            lcout => data_in_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i134_LC_9_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34138\,
            in1 => \N__24015\,
            in2 => \_gnd_net_\,
            in3 => \N__24461\,
            lcout => data_in_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i147_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__34545\,
            in1 => \N__24435\,
            in2 => \N__31237\,
            in3 => \_gnd_net_\,
            lcout => data_in_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i133_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34523\,
            in1 => \N__26764\,
            in2 => \_gnd_net_\,
            in3 => \N__28178\,
            lcout => data_in_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5425_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33270\,
            in1 => \N__29374\,
            in2 => \N__32712\,
            in3 => \N__29217\,
            lcout => \c0.n5779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i105_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34544\,
            in1 => \N__24375\,
            in2 => \_gnd_net_\,
            in3 => \N__24363\,
            lcout => data_in_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i113_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36989\,
            in1 => \N__36205\,
            in2 => \N__24323\,
            in3 => \N__24364\,
            lcout => \c0.data_in_field_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i29_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__24699\,
            in1 => \N__27928\,
            in2 => \N__37271\,
            in3 => \N__36207\,
            lcout => \c0.data_in_field_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_808_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30529\,
            in2 => \_gnd_net_\,
            in3 => \N__24829\,
            lcout => \c0.n1929\,
            ltout => \c0.n1929_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_809_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24316\,
            in1 => \N__32889\,
            in2 => \N__24286\,
            in3 => \N__28844\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30916\,
            in2 => \N__24283\,
            in3 => \N__24697\,
            lcout => \c0.n5204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5485_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__24698\,
            in1 => \N__33315\,
            in2 => \N__32570\,
            in3 => \N__24682\,
            lcout => OPEN,
            ltout => \c0.n5851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5851_bdd_4_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__28916\,
            in1 => \N__24639\,
            in2 => \N__24598\,
            in3 => \N__32475\,
            lcout => \c0.n5408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_984_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26656\,
            in1 => \N__24887\,
            in2 => \_gnd_net_\,
            in3 => \N__27720\,
            lcout => \c0.n5267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i85_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36206\,
            in1 => \N__37218\,
            in2 => \N__26497\,
            in3 => \N__30530\,
            lcout => \c0.data_in_field_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5905_bdd_4_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__28959\,
            in1 => \N__32580\,
            in2 => \N__24550\,
            in3 => \N__25377\,
            lcout => \c0.n5381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_899_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24535\,
            in1 => \N__31093\,
            in2 => \N__24524\,
            in3 => \N__26729\,
            lcout => \c0.n22_adj_1914\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i52_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37152\,
            in1 => \N__36208\,
            in2 => \N__26620\,
            in3 => \N__24932\,
            lcout => \c0.data_in_field_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i67_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__30571\,
            in1 => \N__30721\,
            in2 => \N__36290\,
            in3 => \N__37153\,
            lcout => \c0.data_in_field_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_831_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26655\,
            in2 => \_gnd_net_\,
            in3 => \N__24885\,
            lcout => OPEN,
            ltout => \c0.n1947_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25003\,
            in1 => \N__24909\,
            in2 => \N__24973\,
            in3 => \N__25311\,
            lcout => \c0.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24931\,
            in2 => \_gnd_net_\,
            in3 => \N__30570\,
            lcout => \c0.n1922\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i76_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__24886\,
            in1 => \N__26442\,
            in2 => \N__36291\,
            in3 => \N__37154\,
            lcout => \c0.data_in_field_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5707_bdd_4_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__27340\,
            in1 => \N__32657\,
            in2 => \N__26914\,
            in3 => \N__30753\,
            lcout => \c0.n5474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_826_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25185\,
            in2 => \_gnd_net_\,
            in3 => \N__25106\,
            lcout => \c0.n5105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_974_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25107\,
            in1 => \N__26355\,
            in2 => \N__25196\,
            in3 => \N__28914\,
            lcout => \c0.n26_adj_1884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i99_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36310\,
            in1 => \N__36806\,
            in2 => \N__29065\,
            in3 => \N__24828\,
            lcout => \c0.data_in_field_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i104_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36804\,
            in1 => \N__36311\,
            in2 => \N__24793\,
            in3 => \N__24739\,
            lcout => \c0.data_in_field_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i109_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36309\,
            in1 => \N__36805\,
            in2 => \N__26182\,
            in3 => \N__27179\,
            lcout => \c0.data_in_field_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5500_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33310\,
            in1 => \N__25192\,
            in2 => \N__32628\,
            in3 => \N__25293\,
            lcout => OPEN,
            ltout => \c0.n5875_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5875_bdd_4_lut_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32581\,
            in1 => \N__29607\,
            in2 => \N__25261\,
            in3 => \N__25258\,
            lcout => \c0.n5396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i54_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__28108\,
            in1 => \N__36062\,
            in2 => \N__25200\,
            in3 => \N__37199\,
            lcout => \c0.data_in_field_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i44_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__26574\,
            in1 => \N__36251\,
            in2 => \N__37267\,
            in3 => \N__25039\,
            lcout => \c0.data_in_field_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i125_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__25105\,
            in1 => \N__37195\,
            in2 => \N__28162\,
            in3 => \N__36063\,
            lcout => \c0.data_in_field_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_839_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25160\,
            in2 => \_gnd_net_\,
            in3 => \N__25104\,
            lcout => \c0.n1944\,
            ltout => \c0.n1944_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_864_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33394\,
            in1 => \N__31542\,
            in2 => \N__25063\,
            in3 => \N__28854\,
            lcout => OPEN,
            ltout => \c0.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_865_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27381\,
            in1 => \N__28284\,
            in2 => \N__25060\,
            in3 => \N__25038\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i78_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36085\,
            in1 => \N__37208\,
            in2 => \N__25451\,
            in3 => \N__27513\,
            lcout => \c0.data_in_field_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i40_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37207\,
            in1 => \N__36087\,
            in2 => \N__25588\,
            in3 => \N__25553\,
            lcout => \c0.data_in_field_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_814_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25552\,
            in1 => \N__25519\,
            in2 => \N__25491\,
            in3 => \N__28631\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1871_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_879_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25435\,
            in1 => \N__25870\,
            in2 => \N__25417\,
            in3 => \N__25365\,
            lcout => \c0.n5234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28955\,
            in1 => \N__30451\,
            in2 => \N__28505\,
            in3 => \N__25780\,
            lcout => \c0.n1975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i10_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__30157\,
            in1 => \N__36086\,
            in2 => \N__37269\,
            in3 => \N__25871\,
            lcout => \c0.data_in_field_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i39_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__25366\,
            in1 => \N__28078\,
            in2 => \N__36224\,
            in3 => \N__37212\,
            lcout => \c0.data_in_field_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i128_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25608\,
            in1 => \_gnd_net_\,
            in2 => \N__34547\,
            in3 => \N__27677\,
            lcout => data_in_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i98_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36230\,
            in1 => \N__37276\,
            in2 => \N__29795\,
            in3 => \N__25342\,
            lcout => \c0.data_in_field_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_807_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25691\,
            in2 => \_gnd_net_\,
            in3 => \N__27706\,
            lcout => \c0.n2062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_823_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25749\,
            in2 => \_gnd_net_\,
            in3 => \N__25791\,
            lcout => \c0.n5141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i107_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__37274\,
            in1 => \N__25759\,
            in2 => \N__29095\,
            in3 => \N__36235\,
            lcout => \c0.data_in_field_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i112_LC_10_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__25692\,
            in1 => \N__25726\,
            in2 => \N__36293\,
            in3 => \N__37277\,
            lcout => \c0.data_in_field_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i144_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37273\,
            in1 => \N__36231\,
            in2 => \N__25672\,
            in3 => \N__26020\,
            lcout => \c0.data_in_field_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i129_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36229\,
            in1 => \N__37275\,
            in2 => \N__27612\,
            in3 => \N__29515\,
            lcout => \c0.data_in_field_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i136_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34492\,
            in1 => \N__26019\,
            in2 => \_gnd_net_\,
            in3 => \N__25601\,
            lcout => data_in_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i3_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__25911\,
            in1 => \N__35964\,
            in2 => \N__37289\,
            in3 => \N__27217\,
            lcout => \c0.data_in_field_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i101_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26178\,
            in1 => \N__34491\,
            in2 => \_gnd_net_\,
            in3 => \N__28685\,
            lcout => data_in_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i61_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37261\,
            in1 => \N__35965\,
            in2 => \N__34591\,
            in3 => \N__28003\,
            lcout => \c0.data_in_field_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i144_LC_10_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34498\,
            in1 => \N__26018\,
            in2 => \_gnd_net_\,
            in3 => \N__26050\,
            lcout => data_in_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_828_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30100\,
            in2 => \_gnd_net_\,
            in3 => \N__26702\,
            lcout => OPEN,
            ltout => \c0.n2092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_836_LC_10_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25981\,
            in1 => \N__27973\,
            in2 => \N__25960\,
            in3 => \N__25956\,
            lcout => \c0.n5246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i68_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34490\,
            in1 => \N__26443\,
            in2 => \_gnd_net_\,
            in3 => \N__33518\,
            lcout => data_in_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i52_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34499\,
            in1 => \N__26600\,
            in2 => \_gnd_net_\,
            in3 => \N__33501\,
            lcout => data_in_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_10_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33918\,
            in1 => \N__27455\,
            in2 => \_gnd_net_\,
            in3 => \N__29250\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_10_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27456\,
            in1 => \N__33921\,
            in2 => \_gnd_net_\,
            in3 => \N__25907\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i39_LC_10_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33919\,
            in1 => \N__27240\,
            in2 => \_gnd_net_\,
            in3 => \N__28073\,
            lcout => data_in_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5749_bdd_4_lut_LC_10_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32733\,
            in1 => \N__25881\,
            in2 => \N__25852\,
            in3 => \N__25837\,
            lcout => \c0.n5453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i60_LC_10_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37053\,
            in1 => \N__36312\,
            in2 => \N__26247\,
            in3 => \N__33505\,
            lcout => \c0.data_in_field_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i47_LC_10_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33920\,
            in1 => \N__27239\,
            in2 => \_gnd_net_\,
            in3 => \N__26214\,
            lcout => data_in_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i63_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28131\,
            in1 => \_gnd_net_\,
            in2 => \N__34561\,
            in3 => \N__26510\,
            lcout => data_in_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i109_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31137\,
            in1 => \N__34553\,
            in2 => \_gnd_net_\,
            in3 => \N__26166\,
            lcout => data_in_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i91_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34552\,
            in1 => \N__29055\,
            in2 => \_gnd_net_\,
            in3 => \N__31652\,
            lcout => data_in_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27926\,
            in1 => \N__26143\,
            in2 => \_gnd_net_\,
            in3 => \N__34560\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i116_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34557\,
            in1 => \N__31371\,
            in2 => \_gnd_net_\,
            in3 => \N__31883\,
            lcout => data_in_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i71_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36222\,
            in1 => \N__36705\,
            in2 => \N__28132\,
            in3 => \N__32893\,
            lcout => \c0.data_in_field_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i116_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36704\,
            in1 => \N__36223\,
            in2 => \N__26091\,
            in3 => \N__31884\,
            lcout => \c0.data_in_field_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i66_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26538\,
            in1 => \N__34559\,
            in2 => \_gnd_net_\,
            in3 => \N__30284\,
            lcout => data_in_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i74_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34558\,
            in1 => \N__26537\,
            in2 => \_gnd_net_\,
            in3 => \N__28563\,
            lcout => data_in_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i63_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36952\,
            in1 => \N__35863\,
            in2 => \N__26524\,
            in3 => \N__26663\,
            lcout => \c0.data_in_field_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i77_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34528\,
            in1 => \N__29702\,
            in2 => \_gnd_net_\,
            in3 => \N__26496\,
            lcout => data_in_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i84_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34529\,
            in1 => \N__31810\,
            in2 => \_gnd_net_\,
            in3 => \N__26456\,
            lcout => data_in_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i76_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__34530\,
            in2 => \_gnd_net_\,
            in3 => \N__26432\,
            lcout => data_in_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28882\,
            in1 => \N__31946\,
            in2 => \N__26809\,
            in3 => \N__27178\,
            lcout => \c0.n26_adj_1878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i5_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__26404\,
            in1 => \N__36323\,
            in2 => \N__37086\,
            in3 => \N__28917\,
            lcout => \c0.data_in_field_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i69_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36322\,
            in1 => \N__36889\,
            in2 => \N__34617\,
            in3 => \N__26364\,
            lcout => \c0.data_in_field_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_926_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28867\,
            in1 => \N__27154\,
            in2 => \N__26329\,
            in3 => \N__26302\,
            lcout => \c0.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i87_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34526\,
            in1 => \N__31284\,
            in2 => \_gnd_net_\,
            in3 => \N__29957\,
            lcout => data_in_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i124_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31364\,
            in1 => \N__34527\,
            in2 => \_gnd_net_\,
            in3 => \N__26845\,
            lcout => data_in_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i141_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26807\,
            in1 => \_gnd_net_\,
            in2 => \N__26763\,
            in3 => \N__34525\,
            lcout => data_in_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i141_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__36888\,
            in1 => \N__26759\,
            in2 => \N__36331\,
            in3 => \N__28853\,
            lcout => \c0.data_in_field_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_958_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26728\,
            in1 => \N__28975\,
            in2 => \N__30119\,
            in3 => \N__26664\,
            lcout => \c0.n1795\,
            ltout => \c0.n1795_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_114_2_lut_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26632\,
            in3 => \N__26894\,
            lcout => \c0.n6097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i79_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__36807\,
            in2 => \N__29941\,
            in3 => \N__36327\,
            lcout => \c0.data_in_field_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26930\,
            in1 => \N__26998\,
            in2 => \_gnd_net_\,
            in3 => \N__32852\,
            lcout => \c0.n5179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i44_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34524\,
            in1 => \N__26619\,
            in2 => \_gnd_net_\,
            in3 => \N__26570\,
            lcout => data_in_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_898_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27138\,
            in1 => \N__33393\,
            in2 => \N__27081\,
            in3 => \N__28849\,
            lcout => \c0.n11_adj_1913\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i93_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__26999\,
            in1 => \N__27055\,
            in2 => \N__37005\,
            in3 => \N__36328\,
            lcout => \c0.data_in_field_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i94_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__36329\,
            in1 => \N__26982\,
            in2 => \N__37004\,
            in3 => \N__26936\,
            lcout => \c0.data_in_field_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5375_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33256\,
            in1 => \N__31488\,
            in2 => \N__32679\,
            in3 => \N__29483\,
            lcout => \c0.n5707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i119_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36845\,
            in1 => \N__36083\,
            in2 => \N__28741\,
            in3 => \N__33398\,
            lcout => \c0.data_in_field_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i17_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__36081\,
            in1 => \N__29484\,
            in2 => \N__31459\,
            in3 => \N__36848\,
            lcout => \c0.data_in_field_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_963_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28424\,
            in1 => \N__28714\,
            in2 => \N__28382\,
            in3 => \N__27150\,
            lcout => \c0.n1838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i73_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36082\,
            in1 => \N__36847\,
            in2 => \N__29569\,
            in3 => \N__29457\,
            lcout => \c0.data_in_field_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i41_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36846\,
            in1 => \N__36084\,
            in2 => \N__26878\,
            in3 => \N__28635\,
            lcout => \c0.data_in_field_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_837_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29456\,
            in2 => \_gnd_net_\,
            in3 => \N__29794\,
            lcout => OPEN,
            ltout => \c0.n6_adj_1876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_838_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30450\,
            in1 => \N__30497\,
            in2 => \N__27436\,
            in3 => \N__27425\,
            lcout => \c0.n5129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_987_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27334\,
            in1 => \N__34667\,
            in2 => \_gnd_net_\,
            in3 => \N__34647\,
            lcout => \c0.n6_adj_1874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i1_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__27361\,
            in1 => \N__36256\,
            in2 => \N__37270\,
            in3 => \N__27336\,
            lcout => \c0.data_in_field_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_999_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27335\,
            in1 => \N__27640\,
            in2 => \_gnd_net_\,
            in3 => \N__27311\,
            lcout => \c0.n22_adj_1935\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i35_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36255\,
            in1 => \N__37214\,
            in2 => \N__30616\,
            in3 => \N__28249\,
            lcout => \c0.data_in_field_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i47_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37213\,
            in1 => \N__36257\,
            in2 => \N__27250\,
            in3 => \N__28954\,
            lcout => \c0.data_in_field_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34406\,
            in1 => \N__29169\,
            in2 => \_gnd_net_\,
            in3 => \N__31513\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_815_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27218\,
            in1 => \N__27180\,
            in2 => \N__29284\,
            in3 => \N__29176\,
            lcout => \c0.n5102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i48_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37278\,
            in1 => \N__36254\,
            in2 => \N__27748\,
            in3 => \N__27713\,
            lcout => \c0.data_in_field_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i128_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36252\,
            in1 => \N__37279\,
            in2 => \N__27687\,
            in3 => \N__27641\,
            lcout => \c0.data_in_field_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i129_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34415\,
            in1 => \N__33432\,
            in2 => \_gnd_net_\,
            in3 => \N__27608\,
            lcout => data_in_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i16_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__36253\,
            in1 => \N__27586\,
            in2 => \N__30353\,
            in3 => \N__37280\,
            lcout => \c0.data_in_field_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34416\,
            in1 => \N__30072\,
            in2 => \_gnd_net_\,
            in3 => \N__27919\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i78_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27546\,
            in1 => \N__34417\,
            in2 => \_gnd_net_\,
            in3 => \N__27509\,
            lcout => data_in_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27795\,
            in1 => \_gnd_net_\,
            in2 => \N__34535\,
            in3 => \N__27956\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i53_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34421\,
            in1 => \N__34587\,
            in2 => \_gnd_net_\,
            in3 => \N__30012\,
            lcout => data_in_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27454\,
            lcout => \c0.n22_adj_1952\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i46_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28107\,
            in1 => \_gnd_net_\,
            in2 => \N__34534\,
            in3 => \N__29624\,
            lcout => data_in_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27836\,
            in1 => \N__34408\,
            in2 => \_gnd_net_\,
            in3 => \N__27869\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34407\,
            in1 => \N__28074\,
            in2 => \_gnd_net_\,
            in3 => \N__27837\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i49_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37265\,
            in1 => \N__36101\,
            in2 => \N__30123\,
            in3 => \N__28057\,
            lcout => \c0.data_in_field_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_982_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29590\,
            in1 => \N__27994\,
            in2 => \_gnd_net_\,
            in3 => \N__30337\,
            lcout => \c0.n6_adj_1875\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_947_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31517\,
            in1 => \N__27949\,
            in2 => \N__27927\,
            in3 => \N__27868\,
            lcout => OPEN,
            ltout => \c0.n28_adj_1953_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_953_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30185\,
            in1 => \N__27835\,
            in2 => \N__27820\,
            in3 => \N__27817\,
            lcout => \c0.n30_adj_1959\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i38_LC_11_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33922\,
            in1 => \N__29625\,
            in2 => \_gnd_net_\,
            in3 => \N__27788\,
            lcout => data_in_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35405\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i65_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34538\,
            in1 => \N__29562\,
            in2 => \_gnd_net_\,
            in3 => \N__27759\,
            lcout => data_in_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5415_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33271\,
            in1 => \N__28306\,
            in2 => \N__32627\,
            in3 => \N__30793\,
            lcout => OPEN,
            ltout => \c0.n5773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5773_bdd_4_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32576\,
            in1 => \N__30448\,
            in2 => \N__28261\,
            in3 => \N__28258\,
            lcout => \c0.n5441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i117_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28148\,
            in2 => \N__34536\,
            in3 => \N__31130\,
            lcout => data_in_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5701_bdd_4_lut_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32464\,
            in1 => \N__29129\,
            in2 => \N__30082\,
            in3 => \N__28636\,
            lcout => \c0.n5477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i123_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34428\,
            in1 => \N__33630\,
            in2 => \_gnd_net_\,
            in3 => \N__31967\,
            lcout => data_in_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i125_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28188\,
            in1 => \_gnd_net_\,
            in2 => \N__28155\,
            in3 => \N__34429\,
            lcout => data_in_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i69_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29703\,
            in1 => \_gnd_net_\,
            in2 => \N__34537\,
            in3 => \N__34613\,
            lcout => data_in_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i71_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28130\,
            in1 => \N__29928\,
            in2 => \_gnd_net_\,
            in3 => \N__34430\,
            lcout => data_in_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i115_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34427\,
            in1 => \N__31968\,
            in2 => \_gnd_net_\,
            in3 => \N__30686\,
            lcout => data_in_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i82_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28562\,
            in1 => \N__28608\,
            in2 => \_gnd_net_\,
            in3 => \N__34431\,
            lcout => data_in_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i81_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34449\,
            in1 => \N__28536\,
            in2 => \_gnd_net_\,
            in3 => \N__29906\,
            lcout => data_in_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5911_bdd_4_lut_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32659\,
            in1 => \N__28510\,
            in2 => \N__28480\,
            in3 => \N__28462\,
            lcout => \c0.n5378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_964_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29857\,
            in1 => \N__28366\,
            in2 => \_gnd_net_\,
            in3 => \N__28409\,
            lcout => \c0.n1899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i139_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__28410\,
            in1 => \N__33658\,
            in2 => \N__36313\,
            in3 => \N__36894\,
            lcout => \c0.data_in_field_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i131_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36893\,
            in1 => \N__36266\,
            in2 => \N__33634\,
            in3 => \N__28367\,
            lcout => \c0.data_in_field_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_812_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__30259\,
            in1 => \_gnd_net_\,
            in2 => \N__30787\,
            in3 => \_gnd_net_\,
            lcout => \c0.n5123\,
            ltout => \c0.n5123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_991_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28974\,
            in1 => \N__29029\,
            in2 => \N__28336\,
            in3 => \N__29437\,
            lcout => \c0.n5231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_813_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31480\,
            in2 => \_gnd_net_\,
            in3 => \N__30742\,
            lcout => \c0.n5188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i99_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34541\,
            in1 => \N__29091\,
            in2 => \_gnd_net_\,
            in3 => \N__29043\,
            lcout => data_in_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30258\,
            in1 => \N__29019\,
            in2 => \N__30788\,
            in3 => \N__28973\,
            lcout => OPEN,
            ltout => \c0.n1767_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_994_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28960\,
            in1 => \N__28915\,
            in2 => \N__28885\,
            in3 => \N__28878\,
            lcout => \c0.n5126\,
            ltout => \c0.n5126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_884_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28848\,
            in1 => \N__31083\,
            in2 => \N__28813\,
            in3 => \N__28808\,
            lcout => \c0.n20_adj_1899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i111_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34549\,
            in1 => \N__28737\,
            in2 => \_gnd_net_\,
            in3 => \N__29837\,
            lcout => data_in_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_816_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31575\,
            in1 => \N__31330\,
            in2 => \N__31932\,
            in3 => \N__28654\,
            lcout => \c0.n10_adj_1872\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i101_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36171\,
            in1 => \N__37167\,
            in2 => \N__28707\,
            in3 => \N__28665\,
            lcout => \c0.data_in_field_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_841_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28655\,
            in2 => \_gnd_net_\,
            in3 => \N__28630\,
            lcout => \c0.n1969\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i103_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34548\,
            in1 => \N__31299\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => data_in_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29527\,
            in1 => \N__31999\,
            in2 => \N__29488\,
            in3 => \N__29455\,
            lcout => \c0.n5138\,
            ltout => \c0.n5138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_992_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29361\,
            in1 => \N__29436\,
            in2 => \N__29425\,
            in3 => \N__32162\,
            lcout => \c0.n15_adj_1968\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i27_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__29365\,
            in1 => \N__29413\,
            in2 => \N__37250\,
            in3 => \N__36170\,
            lcout => \c0.data_in_field_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i34_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37054\,
            in1 => \N__36163\,
            in2 => \N__29298\,
            in3 => \N__29334\,
            lcout => \c0.data_in_field_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i19_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__29195\,
            in1 => \N__37060\,
            in2 => \N__29257\,
            in3 => \N__36202\,
            lcout => \c0.data_in_field_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_868_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31693\,
            in1 => \N__29194\,
            in2 => \_gnd_net_\,
            in3 => \N__29113\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i33_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__29114\,
            in1 => \N__29170\,
            in2 => \N__37194\,
            in3 => \N__36203\,
            lcout => \c0.data_in_field_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_844_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29674\,
            in1 => \N__31184\,
            in2 => \_gnd_net_\,
            in3 => \N__31767\,
            lcout => \c0.n5219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i111_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__37059\,
            in1 => \N__29839\,
            in2 => \N__36270\,
            in3 => \N__32166\,
            lcout => \c0.data_in_field_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4988_4_lut_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011000100"
        )
    port map (
            in0 => \N__37438\,
            in1 => \N__37413\,
            in2 => \N__37387\,
            in3 => \N__37462\,
            lcout => n5332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4987_4_lut_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000100010"
        )
    port map (
            in0 => \N__37461\,
            in1 => \N__37383\,
            in2 => \N__37414\,
            in3 => \N__37437\,
            lcout => OPEN,
            ltout => \n5331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4989_3_lut_LC_12_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29824\,
            in2 => \N__29818\,
            in3 => \N__37357\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29675\,
            in1 => \N__31768\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \c0.n1972\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i77_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37058\,
            in1 => \N__36174\,
            in2 => \N__29713\,
            in3 => \N__29676\,
            lcout => \c0.data_in_field_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34413\,
            in1 => \N__30149\,
            in2 => \_gnd_net_\,
            in3 => \N__29645\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i46_LC_12_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37188\,
            in1 => \N__35966\,
            in2 => \N__29629\,
            in3 => \N__29597\,
            lcout => \c0.data_in_field_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i73_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34414\,
            in1 => \N__29550\,
            in2 => \_gnd_net_\,
            in3 => \N__29911\,
            lcout => data_in_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_12_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34412\,
            in1 => \N__30186\,
            in2 => \_gnd_net_\,
            in3 => \N__30148\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i51_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34540\,
            in1 => \N__30806\,
            in2 => \_gnd_net_\,
            in3 => \N__29994\,
            lcout => data_in_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i43_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34539\,
            in1 => \N__30807\,
            in2 => \_gnd_net_\,
            in3 => \N__30462\,
            lcout => data_in_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5356_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__33299\,
            in1 => \N__30915\,
            in2 => \N__30127\,
            in3 => \N__32465\,
            lcout => \c0.n5701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i37_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31599\,
            in1 => \N__34425\,
            in2 => \_gnd_net_\,
            in3 => \N__30053\,
            lcout => data_in_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i45_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34422\,
            in1 => \N__31598\,
            in2 => \_gnd_net_\,
            in3 => \N__30030\,
            lcout => data_in_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i59_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30714\,
            in1 => \N__34426\,
            in2 => \_gnd_net_\,
            in3 => \N__29993\,
            lcout => data_in_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i79_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34424\,
            in1 => \N__29927\,
            in2 => \_gnd_net_\,
            in3 => \N__29970\,
            lcout => data_in_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i81_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37009\,
            in1 => \N__35864\,
            in2 => \N__29875\,
            in3 => \N__29910\,
            lcout => \c0.data_in_field_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i67_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34423\,
            in1 => \N__33558\,
            in2 => \_gnd_net_\,
            in3 => \N__30713\,
            lcout => data_in_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i115_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37006\,
            in1 => \N__36265\,
            in2 => \N__30700\,
            in3 => \N__30648\,
            lcout => \c0.data_in_field_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i35_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34448\,
            in1 => \N__30468\,
            in2 => \_gnd_net_\,
            in3 => \N__30596\,
            lcout => data_in_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32010\,
            in1 => \N__30579\,
            in2 => \N__30547\,
            in3 => \N__30504\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i43_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__36263\,
            in1 => \N__37007\,
            in2 => \N__30449\,
            in3 => \N__30469\,
            lcout => \c0.data_in_field_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_976_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30886\,
            in1 => \N__31936\,
            in2 => \N__30409\,
            in3 => \N__30354\,
            lcout => \c0.n20_adj_1916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i66_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36264\,
            in1 => \N__37008\,
            in2 => \N__30301\,
            in3 => \N__30257\,
            lcout => \c0.data_in_field_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i122_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34446\,
            in1 => \N__30216\,
            in2 => \_gnd_net_\,
            in3 => \N__31154\,
            lcout => data_in_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i114_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31155\,
            in1 => \N__34447\,
            in2 => \_gnd_net_\,
            in3 => \N__30992\,
            lcout => data_in_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i117_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__31107\,
            in1 => \N__37189\,
            in2 => \N__31141\,
            in3 => \N__36217\,
            lcout => \c0.data_in_field_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_842_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31106\,
            in2 => \_gnd_net_\,
            in3 => \N__32960\,
            lcout => \c0.n1815\,
            ltout => \c0.n1815_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30907\,
            in1 => \N__31481\,
            in2 => \N__31072\,
            in3 => \N__31068\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i106_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34542\,
            in1 => \N__30956\,
            in2 => \_gnd_net_\,
            in3 => \N__30999\,
            lcout => data_in_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i57_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__30908\,
            in1 => \N__37190\,
            in2 => \N__30940\,
            in3 => \N__36218\,
            lcout => \c0.data_in_field_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_910_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31247\,
            in2 => \_gnd_net_\,
            in3 => \N__30885\,
            lcout => \c0.n15_adj_1923\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i51_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__30814\,
            in1 => \N__36216\,
            in2 => \N__30792\,
            in3 => \N__36803\,
            lcout => \c0.data_in_field_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i9_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36215\,
            in1 => \N__36802\,
            in2 => \N__31409\,
            in3 => \N__30749\,
            lcout => \c0.data_in_field_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i103_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37184\,
            in1 => \N__36162\,
            in2 => \N__32829\,
            in3 => \N__31306\,
            lcout => \c0.data_in_field_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i45_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36161\,
            in1 => \N__37186\,
            in2 => \N__31609\,
            in3 => \N__31574\,
            lcout => \c0.data_in_field_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_840_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32809\,
            in2 => \_gnd_net_\,
            in3 => \N__32161\,
            lcout => \c0.n1962\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i25_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__36160\,
            in1 => \N__31524\,
            in2 => \N__31489\,
            in3 => \N__37187\,
            lcout => \c0.data_in_field_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31402\,
            in1 => \N__31458\,
            in2 => \_gnd_net_\,
            in3 => \N__34451\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i124_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__36159\,
            in1 => \N__37185\,
            in2 => \N__31378\,
            in3 => \N__31331\,
            lcout => \c0.data_in_field_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i95_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34550\,
            in1 => \N__31305\,
            in2 => \_gnd_net_\,
            in3 => \N__31274\,
            lcout => data_in_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i139_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34450\,
            in1 => \N__33650\,
            in2 => \N__31252\,
            in3 => \_gnd_net_\,
            lcout => data_in_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i75_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__31190\,
            in1 => \N__36168\,
            in2 => \N__33559\,
            in3 => \N__37163\,
            lcout => \c0.data_in_field_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i137_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37165\,
            in1 => \N__36172\,
            in2 => \N__33433\,
            in3 => \N__32006\,
            lcout => \c0.data_in_field_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i123_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__31931\,
            in1 => \N__36167\,
            in2 => \N__31978\,
            in3 => \N__37162\,
            lcout => \c0.data_in_field_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i108_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34500\,
            in1 => \N__31853\,
            in2 => \_gnd_net_\,
            in3 => \N__31894\,
            lcout => data_in_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i100_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31854\,
            in1 => \N__34501\,
            in2 => \_gnd_net_\,
            in3 => \N__31823\,
            lcout => data_in_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i92_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__31824\,
            in1 => \_gnd_net_\,
            in2 => \N__34551\,
            in3 => \N__31799\,
            lcout => data_in_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i92_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__31775\,
            in1 => \N__36169\,
            in2 => \N__31806\,
            in3 => \N__37164\,
            lcout => \c0.data_in_field_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i4_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__37166\,
            in1 => \N__31744\,
            in2 => \N__31709\,
            in3 => \N__36173\,
            lcout => \c0.data_in_field_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i83_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34281\,
            in1 => \N__31671\,
            in2 => \_gnd_net_\,
            in3 => \N__31622\,
            lcout => data_in_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i75_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34280\,
            in1 => \N__33551\,
            in2 => \_gnd_net_\,
            in3 => \N__31623\,
            lcout => data_in_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i60_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34279\,
            in1 => \N__33531\,
            in2 => \_gnd_net_\,
            in3 => \N__33489\,
            lcout => data_in_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i137_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34278\,
            in1 => \N__33419\,
            in2 => \_gnd_net_\,
            in3 => \N__33478\,
            lcout => data_in_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5515_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33316\,
            in1 => \N__33402\,
            in2 => \N__32564\,
            in3 => \N__33361\,
            lcout => \c0.n5893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5520_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__33311\,
            in1 => \N__33001\,
            in2 => \N__32658\,
            in3 => \N__32965\,
            lcout => OPEN,
            ltout => \c0.n5899_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5899_bdd_4_lut_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32713\,
            in1 => \N__32909\,
            in2 => \N__32863\,
            in3 => \N__32860\,
            lcout => \c0.n5384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5893_bdd_4_lut_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__32839\,
            in1 => \N__32825\,
            in2 => \N__32734\,
            in3 => \N__32170\,
            lcout => OPEN,
            ltout => \c0.n5387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__34830\,
            in1 => \N__32140\,
            in2 => \N__32134\,
            in3 => \N__32131\,
            lcout => OPEN,
            ltout => \c0.n5887_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5887_bdd_4_lut_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__32047\,
            in1 => \N__32038\,
            in2 => \N__34834\,
            in3 => \N__34831\,
            lcout => \c0.n5890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_817_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34680\,
            in2 => \_gnd_net_\,
            in3 => \N__34651\,
            lcout => \c0.n1896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i61_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34459\,
            in1 => \N__34618\,
            in2 => \_gnd_net_\,
            in3 => \N__34572\,
            lcout => data_in_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i131_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34458\,
            in1 => \N__33651\,
            in2 => \_gnd_net_\,
            in3 => \N__33615\,
            lcout => data_in_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i0_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33604\,
            in2 => \_gnd_net_\,
            in3 => \N__33598\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => n4437,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i1_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33595\,
            in2 => \_gnd_net_\,
            in3 => \N__33589\,
            lcout => n25,
            ltout => OPEN,
            carryin => n4437,
            carryout => n4438,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i2_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33586\,
            in2 => \_gnd_net_\,
            in3 => \N__33580\,
            lcout => n24,
            ltout => OPEN,
            carryin => n4438,
            carryout => n4439,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i3_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33577\,
            in2 => \_gnd_net_\,
            in3 => \N__33571\,
            lcout => n23,
            ltout => OPEN,
            carryin => n4439,
            carryout => n4440,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i4_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33568\,
            in2 => \_gnd_net_\,
            in3 => \N__33562\,
            lcout => n22,
            ltout => OPEN,
            carryin => n4440,
            carryout => n4441,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i5_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34906\,
            in2 => \_gnd_net_\,
            in3 => \N__34900\,
            lcout => n21,
            ltout => OPEN,
            carryin => n4441,
            carryout => n4442,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i6_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34897\,
            in2 => \_gnd_net_\,
            in3 => \N__34891\,
            lcout => n20,
            ltout => OPEN,
            carryin => n4442,
            carryout => n4443,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i7_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34888\,
            in2 => \_gnd_net_\,
            in3 => \N__34882\,
            lcout => n19,
            ltout => OPEN,
            carryin => n4443,
            carryout => n4444,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i8_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34879\,
            in2 => \_gnd_net_\,
            in3 => \N__34873\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => n4445,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i9_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34870\,
            in2 => \_gnd_net_\,
            in3 => \N__34864\,
            lcout => n17,
            ltout => OPEN,
            carryin => n4445,
            carryout => n4446,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i10_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34861\,
            in2 => \_gnd_net_\,
            in3 => \N__34855\,
            lcout => n16,
            ltout => OPEN,
            carryin => n4446,
            carryout => n4447,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i11_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34852\,
            in2 => \_gnd_net_\,
            in3 => \N__34846\,
            lcout => n15,
            ltout => OPEN,
            carryin => n4447,
            carryout => n4448,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i12_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34843\,
            in2 => \_gnd_net_\,
            in3 => \N__34837\,
            lcout => n14,
            ltout => OPEN,
            carryin => n4448,
            carryout => n4449,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i13_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34978\,
            in2 => \_gnd_net_\,
            in3 => \N__34972\,
            lcout => n13,
            ltout => OPEN,
            carryin => n4449,
            carryout => n4450,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i14_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34969\,
            in2 => \_gnd_net_\,
            in3 => \N__34963\,
            lcout => n12,
            ltout => OPEN,
            carryin => n4450,
            carryout => n4451,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i15_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34960\,
            in2 => \_gnd_net_\,
            in3 => \N__34954\,
            lcout => n11,
            ltout => OPEN,
            carryin => n4451,
            carryout => n4452,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i16_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34951\,
            in2 => \_gnd_net_\,
            in3 => \N__34945\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => n4453,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i17_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34942\,
            in2 => \_gnd_net_\,
            in3 => \N__34936\,
            lcout => n9,
            ltout => OPEN,
            carryin => n4453,
            carryout => n4454,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i18_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34933\,
            in2 => \_gnd_net_\,
            in3 => \N__34927\,
            lcout => n8_adj_1989,
            ltout => OPEN,
            carryin => n4454,
            carryout => n4455,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i19_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34924\,
            in2 => \_gnd_net_\,
            in3 => \N__34918\,
            lcout => n7,
            ltout => OPEN,
            carryin => n4455,
            carryout => n4456,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i20_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34915\,
            in2 => \_gnd_net_\,
            in3 => \N__34909\,
            lcout => n6,
            ltout => OPEN,
            carryin => n4456,
            carryout => n4457,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i21_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37452\,
            in2 => \_gnd_net_\,
            in3 => \N__37441\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n4457,
            carryout => n4458,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i22_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37428\,
            in2 => \_gnd_net_\,
            in3 => \N__37417\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n4458,
            carryout => n4459,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i23_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37401\,
            in2 => \_gnd_net_\,
            in3 => \N__37390\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n4459,
            carryout => n4460,
            clk => \N__35404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i24_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37374\,
            in2 => \_gnd_net_\,
            in3 => \N__37363\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_15_28_0_\,
            carryout => n4461,
            clk => \N__35408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i25_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37350\,
            in2 => \_gnd_net_\,
            in3 => \N__37360\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i157_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__35424\,
            in1 => \N__37339\,
            in2 => \N__37266\,
            in3 => \N__36292\,
            lcout => \c0.data_in_frame_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
