-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jun 29 2019 15:10:02

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    pin9 : out std_logic;
    pin8 : out std_logic;
    pin7 : out std_logic;
    pin6 : in std_logic;
    pin5 : in std_logic;
    pin4 : in std_logic;
    pin3_clk_16mhz : in std_logic;
    pin2_usb_dn : out std_logic;
    pin24 : out std_logic;
    pin23 : out std_logic;
    pin22 : out std_logic;
    pin21 : out std_logic;
    pin20 : out std_logic;
    pin1_usb_dp : out std_logic;
    pin19 : out std_logic;
    pin18 : out std_logic;
    pin17_ss : out std_logic;
    pin16_sck : out std_logic;
    pin15_sdi : out std_logic;
    pin14_sdo : out std_logic;
    pin13 : out std_logic;
    pin12 : out std_logic;
    pin11 : out std_logic;
    pin10 : out std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__69497\ : std_logic;
signal \N__69496\ : std_logic;
signal \N__69495\ : std_logic;
signal \N__69488\ : std_logic;
signal \N__69487\ : std_logic;
signal \N__69486\ : std_logic;
signal \N__69479\ : std_logic;
signal \N__69478\ : std_logic;
signal \N__69477\ : std_logic;
signal \N__69470\ : std_logic;
signal \N__69469\ : std_logic;
signal \N__69468\ : std_logic;
signal \N__69461\ : std_logic;
signal \N__69460\ : std_logic;
signal \N__69459\ : std_logic;
signal \N__69452\ : std_logic;
signal \N__69451\ : std_logic;
signal \N__69450\ : std_logic;
signal \N__69443\ : std_logic;
signal \N__69442\ : std_logic;
signal \N__69441\ : std_logic;
signal \N__69434\ : std_logic;
signal \N__69433\ : std_logic;
signal \N__69432\ : std_logic;
signal \N__69425\ : std_logic;
signal \N__69424\ : std_logic;
signal \N__69423\ : std_logic;
signal \N__69416\ : std_logic;
signal \N__69415\ : std_logic;
signal \N__69414\ : std_logic;
signal \N__69407\ : std_logic;
signal \N__69406\ : std_logic;
signal \N__69405\ : std_logic;
signal \N__69398\ : std_logic;
signal \N__69397\ : std_logic;
signal \N__69396\ : std_logic;
signal \N__69389\ : std_logic;
signal \N__69388\ : std_logic;
signal \N__69387\ : std_logic;
signal \N__69380\ : std_logic;
signal \N__69379\ : std_logic;
signal \N__69378\ : std_logic;
signal \N__69371\ : std_logic;
signal \N__69370\ : std_logic;
signal \N__69369\ : std_logic;
signal \N__69362\ : std_logic;
signal \N__69361\ : std_logic;
signal \N__69360\ : std_logic;
signal \N__69353\ : std_logic;
signal \N__69352\ : std_logic;
signal \N__69351\ : std_logic;
signal \N__69344\ : std_logic;
signal \N__69343\ : std_logic;
signal \N__69342\ : std_logic;
signal \N__69335\ : std_logic;
signal \N__69334\ : std_logic;
signal \N__69333\ : std_logic;
signal \N__69326\ : std_logic;
signal \N__69325\ : std_logic;
signal \N__69324\ : std_logic;
signal \N__69317\ : std_logic;
signal \N__69316\ : std_logic;
signal \N__69315\ : std_logic;
signal \N__69298\ : std_logic;
signal \N__69295\ : std_logic;
signal \N__69294\ : std_logic;
signal \N__69293\ : std_logic;
signal \N__69288\ : std_logic;
signal \N__69285\ : std_logic;
signal \N__69282\ : std_logic;
signal \N__69279\ : std_logic;
signal \N__69276\ : std_logic;
signal \N__69273\ : std_logic;
signal \N__69268\ : std_logic;
signal \N__69265\ : std_logic;
signal \N__69262\ : std_logic;
signal \N__69259\ : std_logic;
signal \N__69256\ : std_logic;
signal \N__69253\ : std_logic;
signal \N__69252\ : std_logic;
signal \N__69251\ : std_logic;
signal \N__69246\ : std_logic;
signal \N__69243\ : std_logic;
signal \N__69240\ : std_logic;
signal \N__69237\ : std_logic;
signal \N__69234\ : std_logic;
signal \N__69231\ : std_logic;
signal \N__69226\ : std_logic;
signal \N__69223\ : std_logic;
signal \N__69220\ : std_logic;
signal \N__69217\ : std_logic;
signal \N__69214\ : std_logic;
signal \N__69211\ : std_logic;
signal \N__69208\ : std_logic;
signal \N__69205\ : std_logic;
signal \N__69204\ : std_logic;
signal \N__69203\ : std_logic;
signal \N__69200\ : std_logic;
signal \N__69197\ : std_logic;
signal \N__69194\ : std_logic;
signal \N__69191\ : std_logic;
signal \N__69186\ : std_logic;
signal \N__69183\ : std_logic;
signal \N__69180\ : std_logic;
signal \N__69175\ : std_logic;
signal \N__69172\ : std_logic;
signal \N__69169\ : std_logic;
signal \N__69166\ : std_logic;
signal \N__69163\ : std_logic;
signal \N__69160\ : std_logic;
signal \N__69157\ : std_logic;
signal \N__69156\ : std_logic;
signal \N__69155\ : std_logic;
signal \N__69150\ : std_logic;
signal \N__69147\ : std_logic;
signal \N__69144\ : std_logic;
signal \N__69141\ : std_logic;
signal \N__69136\ : std_logic;
signal \N__69133\ : std_logic;
signal \N__69130\ : std_logic;
signal \N__69127\ : std_logic;
signal \N__69124\ : std_logic;
signal \N__69121\ : std_logic;
signal \N__69118\ : std_logic;
signal \N__69115\ : std_logic;
signal \N__69112\ : std_logic;
signal \N__69109\ : std_logic;
signal \N__69108\ : std_logic;
signal \N__69107\ : std_logic;
signal \N__69102\ : std_logic;
signal \N__69099\ : std_logic;
signal \N__69096\ : std_logic;
signal \N__69093\ : std_logic;
signal \N__69090\ : std_logic;
signal \N__69087\ : std_logic;
signal \N__69084\ : std_logic;
signal \N__69081\ : std_logic;
signal \N__69076\ : std_logic;
signal \N__69073\ : std_logic;
signal \N__69072\ : std_logic;
signal \N__69071\ : std_logic;
signal \N__69068\ : std_logic;
signal \N__69067\ : std_logic;
signal \N__69064\ : std_logic;
signal \N__69063\ : std_logic;
signal \N__69060\ : std_logic;
signal \N__69059\ : std_logic;
signal \N__69046\ : std_logic;
signal \N__69045\ : std_logic;
signal \N__69044\ : std_logic;
signal \N__69043\ : std_logic;
signal \N__69040\ : std_logic;
signal \N__69037\ : std_logic;
signal \N__69032\ : std_logic;
signal \N__69025\ : std_logic;
signal \N__69022\ : std_logic;
signal \N__69019\ : std_logic;
signal \N__69016\ : std_logic;
signal \N__69013\ : std_logic;
signal \N__69010\ : std_logic;
signal \N__69007\ : std_logic;
signal \N__69006\ : std_logic;
signal \N__69003\ : std_logic;
signal \N__69000\ : std_logic;
signal \N__68997\ : std_logic;
signal \N__68994\ : std_logic;
signal \N__68991\ : std_logic;
signal \N__68988\ : std_logic;
signal \N__68983\ : std_logic;
signal \N__68980\ : std_logic;
signal \N__68977\ : std_logic;
signal \N__68974\ : std_logic;
signal \N__68971\ : std_logic;
signal \N__68968\ : std_logic;
signal \N__68965\ : std_logic;
signal \N__68962\ : std_logic;
signal \N__68961\ : std_logic;
signal \N__68958\ : std_logic;
signal \N__68955\ : std_logic;
signal \N__68952\ : std_logic;
signal \N__68949\ : std_logic;
signal \N__68944\ : std_logic;
signal \N__68943\ : std_logic;
signal \N__68942\ : std_logic;
signal \N__68937\ : std_logic;
signal \N__68936\ : std_logic;
signal \N__68933\ : std_logic;
signal \N__68930\ : std_logic;
signal \N__68927\ : std_logic;
signal \N__68924\ : std_logic;
signal \N__68919\ : std_logic;
signal \N__68914\ : std_logic;
signal \N__68911\ : std_logic;
signal \N__68910\ : std_logic;
signal \N__68907\ : std_logic;
signal \N__68904\ : std_logic;
signal \N__68901\ : std_logic;
signal \N__68898\ : std_logic;
signal \N__68895\ : std_logic;
signal \N__68890\ : std_logic;
signal \N__68887\ : std_logic;
signal \N__68884\ : std_logic;
signal \N__68881\ : std_logic;
signal \N__68878\ : std_logic;
signal \N__68875\ : std_logic;
signal \N__68872\ : std_logic;
signal \N__68871\ : std_logic;
signal \N__68866\ : std_logic;
signal \N__68863\ : std_logic;
signal \N__68862\ : std_logic;
signal \N__68861\ : std_logic;
signal \N__68858\ : std_logic;
signal \N__68855\ : std_logic;
signal \N__68852\ : std_logic;
signal \N__68845\ : std_logic;
signal \N__68842\ : std_logic;
signal \N__68839\ : std_logic;
signal \N__68836\ : std_logic;
signal \N__68833\ : std_logic;
signal \N__68830\ : std_logic;
signal \N__68829\ : std_logic;
signal \N__68826\ : std_logic;
signal \N__68823\ : std_logic;
signal \N__68818\ : std_logic;
signal \N__68815\ : std_logic;
signal \N__68812\ : std_logic;
signal \N__68809\ : std_logic;
signal \N__68806\ : std_logic;
signal \N__68803\ : std_logic;
signal \N__68800\ : std_logic;
signal \N__68799\ : std_logic;
signal \N__68794\ : std_logic;
signal \N__68793\ : std_logic;
signal \N__68792\ : std_logic;
signal \N__68789\ : std_logic;
signal \N__68786\ : std_logic;
signal \N__68783\ : std_logic;
signal \N__68776\ : std_logic;
signal \N__68773\ : std_logic;
signal \N__68770\ : std_logic;
signal \N__68769\ : std_logic;
signal \N__68766\ : std_logic;
signal \N__68763\ : std_logic;
signal \N__68760\ : std_logic;
signal \N__68757\ : std_logic;
signal \N__68754\ : std_logic;
signal \N__68751\ : std_logic;
signal \N__68746\ : std_logic;
signal \N__68743\ : std_logic;
signal \N__68740\ : std_logic;
signal \N__68737\ : std_logic;
signal \N__68734\ : std_logic;
signal \N__68731\ : std_logic;
signal \N__68728\ : std_logic;
signal \N__68727\ : std_logic;
signal \N__68722\ : std_logic;
signal \N__68721\ : std_logic;
signal \N__68720\ : std_logic;
signal \N__68717\ : std_logic;
signal \N__68714\ : std_logic;
signal \N__68711\ : std_logic;
signal \N__68704\ : std_logic;
signal \N__68701\ : std_logic;
signal \N__68698\ : std_logic;
signal \N__68697\ : std_logic;
signal \N__68694\ : std_logic;
signal \N__68691\ : std_logic;
signal \N__68688\ : std_logic;
signal \N__68685\ : std_logic;
signal \N__68682\ : std_logic;
signal \N__68679\ : std_logic;
signal \N__68674\ : std_logic;
signal \N__68671\ : std_logic;
signal \N__68668\ : std_logic;
signal \N__68665\ : std_logic;
signal \N__68662\ : std_logic;
signal \N__68659\ : std_logic;
signal \N__68658\ : std_logic;
signal \N__68653\ : std_logic;
signal \N__68650\ : std_logic;
signal \N__68649\ : std_logic;
signal \N__68648\ : std_logic;
signal \N__68645\ : std_logic;
signal \N__68642\ : std_logic;
signal \N__68639\ : std_logic;
signal \N__68636\ : std_logic;
signal \N__68631\ : std_logic;
signal \N__68626\ : std_logic;
signal \N__68623\ : std_logic;
signal \N__68620\ : std_logic;
signal \N__68617\ : std_logic;
signal \N__68614\ : std_logic;
signal \N__68611\ : std_logic;
signal \N__68608\ : std_logic;
signal \N__68607\ : std_logic;
signal \N__68602\ : std_logic;
signal \N__68601\ : std_logic;
signal \N__68598\ : std_logic;
signal \N__68595\ : std_logic;
signal \N__68594\ : std_logic;
signal \N__68591\ : std_logic;
signal \N__68588\ : std_logic;
signal \N__68585\ : std_logic;
signal \N__68582\ : std_logic;
signal \N__68577\ : std_logic;
signal \N__68572\ : std_logic;
signal \N__68569\ : std_logic;
signal \N__68566\ : std_logic;
signal \N__68563\ : std_logic;
signal \N__68560\ : std_logic;
signal \N__68557\ : std_logic;
signal \N__68554\ : std_logic;
signal \N__68551\ : std_logic;
signal \N__68550\ : std_logic;
signal \N__68549\ : std_logic;
signal \N__68546\ : std_logic;
signal \N__68543\ : std_logic;
signal \N__68540\ : std_logic;
signal \N__68537\ : std_logic;
signal \N__68534\ : std_logic;
signal \N__68531\ : std_logic;
signal \N__68528\ : std_logic;
signal \N__68523\ : std_logic;
signal \N__68518\ : std_logic;
signal \N__68515\ : std_logic;
signal \N__68512\ : std_logic;
signal \N__68509\ : std_logic;
signal \N__68506\ : std_logic;
signal \N__68503\ : std_logic;
signal \N__68500\ : std_logic;
signal \N__68497\ : std_logic;
signal \N__68496\ : std_logic;
signal \N__68493\ : std_logic;
signal \N__68490\ : std_logic;
signal \N__68487\ : std_logic;
signal \N__68484\ : std_logic;
signal \N__68479\ : std_logic;
signal \N__68476\ : std_logic;
signal \N__68473\ : std_logic;
signal \N__68470\ : std_logic;
signal \N__68467\ : std_logic;
signal \N__68464\ : std_logic;
signal \N__68461\ : std_logic;
signal \N__68460\ : std_logic;
signal \N__68459\ : std_logic;
signal \N__68456\ : std_logic;
signal \N__68453\ : std_logic;
signal \N__68450\ : std_logic;
signal \N__68445\ : std_logic;
signal \N__68440\ : std_logic;
signal \N__68437\ : std_logic;
signal \N__68436\ : std_logic;
signal \N__68435\ : std_logic;
signal \N__68434\ : std_logic;
signal \N__68429\ : std_logic;
signal \N__68428\ : std_logic;
signal \N__68427\ : std_logic;
signal \N__68426\ : std_logic;
signal \N__68423\ : std_logic;
signal \N__68422\ : std_logic;
signal \N__68419\ : std_logic;
signal \N__68418\ : std_logic;
signal \N__68415\ : std_logic;
signal \N__68412\ : std_logic;
signal \N__68411\ : std_logic;
signal \N__68408\ : std_logic;
signal \N__68407\ : std_logic;
signal \N__68404\ : std_logic;
signal \N__68403\ : std_logic;
signal \N__68402\ : std_logic;
signal \N__68401\ : std_logic;
signal \N__68400\ : std_logic;
signal \N__68399\ : std_logic;
signal \N__68398\ : std_logic;
signal \N__68397\ : std_logic;
signal \N__68396\ : std_logic;
signal \N__68395\ : std_logic;
signal \N__68394\ : std_logic;
signal \N__68393\ : std_logic;
signal \N__68392\ : std_logic;
signal \N__68391\ : std_logic;
signal \N__68390\ : std_logic;
signal \N__68387\ : std_logic;
signal \N__68384\ : std_logic;
signal \N__68379\ : std_logic;
signal \N__68374\ : std_logic;
signal \N__68365\ : std_logic;
signal \N__68364\ : std_logic;
signal \N__68361\ : std_logic;
signal \N__68360\ : std_logic;
signal \N__68357\ : std_logic;
signal \N__68356\ : std_logic;
signal \N__68353\ : std_logic;
signal \N__68352\ : std_logic;
signal \N__68349\ : std_logic;
signal \N__68348\ : std_logic;
signal \N__68345\ : std_logic;
signal \N__68344\ : std_logic;
signal \N__68341\ : std_logic;
signal \N__68340\ : std_logic;
signal \N__68337\ : std_logic;
signal \N__68336\ : std_logic;
signal \N__68333\ : std_logic;
signal \N__68332\ : std_logic;
signal \N__68329\ : std_logic;
signal \N__68326\ : std_logic;
signal \N__68323\ : std_logic;
signal \N__68320\ : std_logic;
signal \N__68317\ : std_logic;
signal \N__68314\ : std_logic;
signal \N__68311\ : std_logic;
signal \N__68306\ : std_logic;
signal \N__68303\ : std_logic;
signal \N__68300\ : std_logic;
signal \N__68283\ : std_logic;
signal \N__68266\ : std_logic;
signal \N__68257\ : std_logic;
signal \N__68250\ : std_logic;
signal \N__68247\ : std_logic;
signal \N__68244\ : std_logic;
signal \N__68231\ : std_logic;
signal \N__68226\ : std_logic;
signal \N__68223\ : std_logic;
signal \N__68218\ : std_logic;
signal \N__68215\ : std_logic;
signal \N__68214\ : std_logic;
signal \N__68211\ : std_logic;
signal \N__68208\ : std_logic;
signal \N__68203\ : std_logic;
signal \N__68200\ : std_logic;
signal \N__68197\ : std_logic;
signal \N__68194\ : std_logic;
signal \N__68191\ : std_logic;
signal \N__68188\ : std_logic;
signal \N__68187\ : std_logic;
signal \N__68184\ : std_logic;
signal \N__68181\ : std_logic;
signal \N__68180\ : std_logic;
signal \N__68179\ : std_logic;
signal \N__68174\ : std_logic;
signal \N__68171\ : std_logic;
signal \N__68168\ : std_logic;
signal \N__68165\ : std_logic;
signal \N__68162\ : std_logic;
signal \N__68159\ : std_logic;
signal \N__68156\ : std_logic;
signal \N__68151\ : std_logic;
signal \N__68146\ : std_logic;
signal \N__68143\ : std_logic;
signal \N__68140\ : std_logic;
signal \N__68137\ : std_logic;
signal \N__68136\ : std_logic;
signal \N__68133\ : std_logic;
signal \N__68130\ : std_logic;
signal \N__68125\ : std_logic;
signal \N__68122\ : std_logic;
signal \N__68119\ : std_logic;
signal \N__68116\ : std_logic;
signal \N__68113\ : std_logic;
signal \N__68110\ : std_logic;
signal \N__68107\ : std_logic;
signal \N__68106\ : std_logic;
signal \N__68101\ : std_logic;
signal \N__68100\ : std_logic;
signal \N__68099\ : std_logic;
signal \N__68096\ : std_logic;
signal \N__68091\ : std_logic;
signal \N__68086\ : std_logic;
signal \N__68083\ : std_logic;
signal \N__68080\ : std_logic;
signal \N__68077\ : std_logic;
signal \N__68076\ : std_logic;
signal \N__68073\ : std_logic;
signal \N__68070\ : std_logic;
signal \N__68065\ : std_logic;
signal \N__68062\ : std_logic;
signal \N__68059\ : std_logic;
signal \N__68056\ : std_logic;
signal \N__68053\ : std_logic;
signal \N__68050\ : std_logic;
signal \N__68049\ : std_logic;
signal \N__68048\ : std_logic;
signal \N__68047\ : std_logic;
signal \N__68042\ : std_logic;
signal \N__68037\ : std_logic;
signal \N__68034\ : std_logic;
signal \N__68031\ : std_logic;
signal \N__68028\ : std_logic;
signal \N__68025\ : std_logic;
signal \N__68020\ : std_logic;
signal \N__68017\ : std_logic;
signal \N__68014\ : std_logic;
signal \N__68013\ : std_logic;
signal \N__68010\ : std_logic;
signal \N__68007\ : std_logic;
signal \N__68004\ : std_logic;
signal \N__68001\ : std_logic;
signal \N__67996\ : std_logic;
signal \N__67993\ : std_logic;
signal \N__67990\ : std_logic;
signal \N__67987\ : std_logic;
signal \N__67984\ : std_logic;
signal \N__67981\ : std_logic;
signal \N__67978\ : std_logic;
signal \N__67977\ : std_logic;
signal \N__67974\ : std_logic;
signal \N__67971\ : std_logic;
signal \N__67970\ : std_logic;
signal \N__67965\ : std_logic;
signal \N__67964\ : std_logic;
signal \N__67961\ : std_logic;
signal \N__67958\ : std_logic;
signal \N__67955\ : std_logic;
signal \N__67952\ : std_logic;
signal \N__67949\ : std_logic;
signal \N__67946\ : std_logic;
signal \N__67943\ : std_logic;
signal \N__67936\ : std_logic;
signal \N__67933\ : std_logic;
signal \N__67930\ : std_logic;
signal \N__67929\ : std_logic;
signal \N__67926\ : std_logic;
signal \N__67923\ : std_logic;
signal \N__67918\ : std_logic;
signal \N__67915\ : std_logic;
signal \N__67912\ : std_logic;
signal \N__67909\ : std_logic;
signal \N__67906\ : std_logic;
signal \N__67903\ : std_logic;
signal \N__67900\ : std_logic;
signal \N__67899\ : std_logic;
signal \N__67898\ : std_logic;
signal \N__67895\ : std_logic;
signal \N__67892\ : std_logic;
signal \N__67889\ : std_logic;
signal \N__67886\ : std_logic;
signal \N__67885\ : std_logic;
signal \N__67880\ : std_logic;
signal \N__67877\ : std_logic;
signal \N__67874\ : std_logic;
signal \N__67867\ : std_logic;
signal \N__67864\ : std_logic;
signal \N__67861\ : std_logic;
signal \N__67858\ : std_logic;
signal \N__67855\ : std_logic;
signal \N__67852\ : std_logic;
signal \N__67849\ : std_logic;
signal \N__67846\ : std_logic;
signal \N__67843\ : std_logic;
signal \N__67842\ : std_logic;
signal \N__67839\ : std_logic;
signal \N__67836\ : std_logic;
signal \N__67833\ : std_logic;
signal \N__67830\ : std_logic;
signal \N__67825\ : std_logic;
signal \N__67822\ : std_logic;
signal \N__67819\ : std_logic;
signal \N__67816\ : std_logic;
signal \N__67813\ : std_logic;
signal \N__67810\ : std_logic;
signal \N__67809\ : std_logic;
signal \N__67806\ : std_logic;
signal \N__67803\ : std_logic;
signal \N__67798\ : std_logic;
signal \N__67795\ : std_logic;
signal \N__67792\ : std_logic;
signal \N__67789\ : std_logic;
signal \N__67786\ : std_logic;
signal \N__67783\ : std_logic;
signal \N__67780\ : std_logic;
signal \N__67779\ : std_logic;
signal \N__67776\ : std_logic;
signal \N__67773\ : std_logic;
signal \N__67768\ : std_logic;
signal \N__67765\ : std_logic;
signal \N__67762\ : std_logic;
signal \N__67759\ : std_logic;
signal \N__67758\ : std_logic;
signal \N__67755\ : std_logic;
signal \N__67752\ : std_logic;
signal \N__67747\ : std_logic;
signal \N__67744\ : std_logic;
signal \N__67741\ : std_logic;
signal \N__67738\ : std_logic;
signal \N__67735\ : std_logic;
signal \N__67732\ : std_logic;
signal \N__67729\ : std_logic;
signal \N__67728\ : std_logic;
signal \N__67725\ : std_logic;
signal \N__67722\ : std_logic;
signal \N__67717\ : std_logic;
signal \N__67714\ : std_logic;
signal \N__67711\ : std_logic;
signal \N__67708\ : std_logic;
signal \N__67705\ : std_logic;
signal \N__67702\ : std_logic;
signal \N__67699\ : std_logic;
signal \N__67696\ : std_logic;
signal \N__67695\ : std_logic;
signal \N__67692\ : std_logic;
signal \N__67689\ : std_logic;
signal \N__67686\ : std_logic;
signal \N__67683\ : std_logic;
signal \N__67678\ : std_logic;
signal \N__67677\ : std_logic;
signal \N__67674\ : std_logic;
signal \N__67673\ : std_logic;
signal \N__67670\ : std_logic;
signal \N__67667\ : std_logic;
signal \N__67664\ : std_logic;
signal \N__67661\ : std_logic;
signal \N__67654\ : std_logic;
signal \N__67651\ : std_logic;
signal \N__67650\ : std_logic;
signal \N__67647\ : std_logic;
signal \N__67644\ : std_logic;
signal \N__67641\ : std_logic;
signal \N__67638\ : std_logic;
signal \N__67633\ : std_logic;
signal \N__67630\ : std_logic;
signal \N__67627\ : std_logic;
signal \N__67624\ : std_logic;
signal \N__67621\ : std_logic;
signal \N__67618\ : std_logic;
signal \N__67617\ : std_logic;
signal \N__67612\ : std_logic;
signal \N__67611\ : std_logic;
signal \N__67610\ : std_logic;
signal \N__67607\ : std_logic;
signal \N__67604\ : std_logic;
signal \N__67601\ : std_logic;
signal \N__67596\ : std_logic;
signal \N__67591\ : std_logic;
signal \N__67588\ : std_logic;
signal \N__67585\ : std_logic;
signal \N__67582\ : std_logic;
signal \N__67581\ : std_logic;
signal \N__67578\ : std_logic;
signal \N__67575\ : std_logic;
signal \N__67570\ : std_logic;
signal \N__67567\ : std_logic;
signal \N__67564\ : std_logic;
signal \N__67561\ : std_logic;
signal \N__67558\ : std_logic;
signal \N__67555\ : std_logic;
signal \N__67554\ : std_logic;
signal \N__67549\ : std_logic;
signal \N__67548\ : std_logic;
signal \N__67547\ : std_logic;
signal \N__67544\ : std_logic;
signal \N__67541\ : std_logic;
signal \N__67538\ : std_logic;
signal \N__67535\ : std_logic;
signal \N__67530\ : std_logic;
signal \N__67525\ : std_logic;
signal \N__67522\ : std_logic;
signal \N__67519\ : std_logic;
signal \N__67516\ : std_logic;
signal \N__67513\ : std_logic;
signal \N__67510\ : std_logic;
signal \N__67507\ : std_logic;
signal \N__67504\ : std_logic;
signal \N__67503\ : std_logic;
signal \N__67500\ : std_logic;
signal \N__67497\ : std_logic;
signal \N__67492\ : std_logic;
signal \N__67489\ : std_logic;
signal \N__67486\ : std_logic;
signal \N__67485\ : std_logic;
signal \N__67482\ : std_logic;
signal \N__67479\ : std_logic;
signal \N__67474\ : std_logic;
signal \N__67471\ : std_logic;
signal \N__67468\ : std_logic;
signal \N__67467\ : std_logic;
signal \N__67466\ : std_logic;
signal \N__67465\ : std_logic;
signal \N__67464\ : std_logic;
signal \N__67463\ : std_logic;
signal \N__67462\ : std_logic;
signal \N__67461\ : std_logic;
signal \N__67460\ : std_logic;
signal \N__67459\ : std_logic;
signal \N__67458\ : std_logic;
signal \N__67457\ : std_logic;
signal \N__67456\ : std_logic;
signal \N__67455\ : std_logic;
signal \N__67452\ : std_logic;
signal \N__67449\ : std_logic;
signal \N__67446\ : std_logic;
signal \N__67443\ : std_logic;
signal \N__67442\ : std_logic;
signal \N__67439\ : std_logic;
signal \N__67436\ : std_logic;
signal \N__67433\ : std_logic;
signal \N__67430\ : std_logic;
signal \N__67427\ : std_logic;
signal \N__67426\ : std_logic;
signal \N__67425\ : std_logic;
signal \N__67422\ : std_logic;
signal \N__67421\ : std_logic;
signal \N__67418\ : std_logic;
signal \N__67417\ : std_logic;
signal \N__67414\ : std_logic;
signal \N__67413\ : std_logic;
signal \N__67410\ : std_logic;
signal \N__67409\ : std_logic;
signal \N__67406\ : std_logic;
signal \N__67405\ : std_logic;
signal \N__67404\ : std_logic;
signal \N__67401\ : std_logic;
signal \N__67398\ : std_logic;
signal \N__67397\ : std_logic;
signal \N__67396\ : std_logic;
signal \N__67395\ : std_logic;
signal \N__67392\ : std_logic;
signal \N__67389\ : std_logic;
signal \N__67386\ : std_logic;
signal \N__67381\ : std_logic;
signal \N__67372\ : std_logic;
signal \N__67355\ : std_logic;
signal \N__67352\ : std_logic;
signal \N__67351\ : std_logic;
signal \N__67348\ : std_logic;
signal \N__67345\ : std_logic;
signal \N__67342\ : std_logic;
signal \N__67337\ : std_logic;
signal \N__67334\ : std_logic;
signal \N__67331\ : std_logic;
signal \N__67328\ : std_logic;
signal \N__67323\ : std_logic;
signal \N__67320\ : std_logic;
signal \N__67315\ : std_logic;
signal \N__67312\ : std_logic;
signal \N__67309\ : std_logic;
signal \N__67306\ : std_logic;
signal \N__67303\ : std_logic;
signal \N__67300\ : std_logic;
signal \N__67297\ : std_logic;
signal \N__67296\ : std_logic;
signal \N__67293\ : std_logic;
signal \N__67290\ : std_logic;
signal \N__67287\ : std_logic;
signal \N__67284\ : std_logic;
signal \N__67279\ : std_logic;
signal \N__67272\ : std_logic;
signal \N__67269\ : std_logic;
signal \N__67262\ : std_logic;
signal \N__67259\ : std_logic;
signal \N__67254\ : std_logic;
signal \N__67243\ : std_logic;
signal \N__67240\ : std_logic;
signal \N__67237\ : std_logic;
signal \N__67234\ : std_logic;
signal \N__67227\ : std_logic;
signal \N__67224\ : std_logic;
signal \N__67221\ : std_logic;
signal \N__67216\ : std_logic;
signal \N__67213\ : std_logic;
signal \N__67210\ : std_logic;
signal \N__67207\ : std_logic;
signal \N__67204\ : std_logic;
signal \N__67203\ : std_logic;
signal \N__67200\ : std_logic;
signal \N__67197\ : std_logic;
signal \N__67192\ : std_logic;
signal \N__67189\ : std_logic;
signal \N__67186\ : std_logic;
signal \N__67183\ : std_logic;
signal \N__67180\ : std_logic;
signal \N__67177\ : std_logic;
signal \N__67174\ : std_logic;
signal \N__67171\ : std_logic;
signal \N__67168\ : std_logic;
signal \N__67165\ : std_logic;
signal \N__67162\ : std_logic;
signal \N__67161\ : std_logic;
signal \N__67158\ : std_logic;
signal \N__67155\ : std_logic;
signal \N__67150\ : std_logic;
signal \N__67147\ : std_logic;
signal \N__67144\ : std_logic;
signal \N__67141\ : std_logic;
signal \N__67138\ : std_logic;
signal \N__67135\ : std_logic;
signal \N__67132\ : std_logic;
signal \N__67129\ : std_logic;
signal \N__67126\ : std_logic;
signal \N__67123\ : std_logic;
signal \N__67120\ : std_logic;
signal \N__67117\ : std_logic;
signal \N__67116\ : std_logic;
signal \N__67113\ : std_logic;
signal \N__67110\ : std_logic;
signal \N__67105\ : std_logic;
signal \N__67102\ : std_logic;
signal \N__67099\ : std_logic;
signal \N__67096\ : std_logic;
signal \N__67093\ : std_logic;
signal \N__67090\ : std_logic;
signal \N__67087\ : std_logic;
signal \N__67084\ : std_logic;
signal \N__67081\ : std_logic;
signal \N__67078\ : std_logic;
signal \N__67077\ : std_logic;
signal \N__67074\ : std_logic;
signal \N__67071\ : std_logic;
signal \N__67066\ : std_logic;
signal \N__67063\ : std_logic;
signal \N__67060\ : std_logic;
signal \N__67057\ : std_logic;
signal \N__67054\ : std_logic;
signal \N__67051\ : std_logic;
signal \N__67048\ : std_logic;
signal \N__67045\ : std_logic;
signal \N__67042\ : std_logic;
signal \N__67039\ : std_logic;
signal \N__67036\ : std_logic;
signal \N__67033\ : std_logic;
signal \N__67032\ : std_logic;
signal \N__67029\ : std_logic;
signal \N__67026\ : std_logic;
signal \N__67021\ : std_logic;
signal \N__67018\ : std_logic;
signal \N__67015\ : std_logic;
signal \N__67012\ : std_logic;
signal \N__67009\ : std_logic;
signal \N__67006\ : std_logic;
signal \N__67003\ : std_logic;
signal \N__67000\ : std_logic;
signal \N__66997\ : std_logic;
signal \N__66994\ : std_logic;
signal \N__66991\ : std_logic;
signal \N__66988\ : std_logic;
signal \N__66985\ : std_logic;
signal \N__66982\ : std_logic;
signal \N__66979\ : std_logic;
signal \N__66976\ : std_logic;
signal \N__66973\ : std_logic;
signal \N__66970\ : std_logic;
signal \N__66967\ : std_logic;
signal \N__66964\ : std_logic;
signal \N__66961\ : std_logic;
signal \N__66958\ : std_logic;
signal \N__66955\ : std_logic;
signal \N__66952\ : std_logic;
signal \N__66949\ : std_logic;
signal \N__66946\ : std_logic;
signal \N__66943\ : std_logic;
signal \N__66940\ : std_logic;
signal \N__66937\ : std_logic;
signal \N__66934\ : std_logic;
signal \N__66931\ : std_logic;
signal \N__66930\ : std_logic;
signal \N__66929\ : std_logic;
signal \N__66928\ : std_logic;
signal \N__66927\ : std_logic;
signal \N__66926\ : std_logic;
signal \N__66925\ : std_logic;
signal \N__66924\ : std_logic;
signal \N__66923\ : std_logic;
signal \N__66922\ : std_logic;
signal \N__66921\ : std_logic;
signal \N__66920\ : std_logic;
signal \N__66917\ : std_logic;
signal \N__66914\ : std_logic;
signal \N__66913\ : std_logic;
signal \N__66910\ : std_logic;
signal \N__66907\ : std_logic;
signal \N__66904\ : std_logic;
signal \N__66901\ : std_logic;
signal \N__66898\ : std_logic;
signal \N__66895\ : std_logic;
signal \N__66892\ : std_logic;
signal \N__66891\ : std_logic;
signal \N__66890\ : std_logic;
signal \N__66889\ : std_logic;
signal \N__66888\ : std_logic;
signal \N__66885\ : std_logic;
signal \N__66884\ : std_logic;
signal \N__66881\ : std_logic;
signal \N__66880\ : std_logic;
signal \N__66877\ : std_logic;
signal \N__66876\ : std_logic;
signal \N__66875\ : std_logic;
signal \N__66870\ : std_logic;
signal \N__66861\ : std_logic;
signal \N__66852\ : std_logic;
signal \N__66849\ : std_logic;
signal \N__66846\ : std_logic;
signal \N__66843\ : std_logic;
signal \N__66840\ : std_logic;
signal \N__66837\ : std_logic;
signal \N__66834\ : std_logic;
signal \N__66831\ : std_logic;
signal \N__66830\ : std_logic;
signal \N__66829\ : std_logic;
signal \N__66828\ : std_logic;
signal \N__66825\ : std_logic;
signal \N__66824\ : std_logic;
signal \N__66823\ : std_logic;
signal \N__66822\ : std_logic;
signal \N__66819\ : std_logic;
signal \N__66816\ : std_logic;
signal \N__66813\ : std_logic;
signal \N__66808\ : std_logic;
signal \N__66805\ : std_logic;
signal \N__66796\ : std_logic;
signal \N__66789\ : std_logic;
signal \N__66786\ : std_logic;
signal \N__66783\ : std_logic;
signal \N__66782\ : std_logic;
signal \N__66779\ : std_logic;
signal \N__66776\ : std_logic;
signal \N__66773\ : std_logic;
signal \N__66770\ : std_logic;
signal \N__66767\ : std_logic;
signal \N__66764\ : std_logic;
signal \N__66761\ : std_logic;
signal \N__66760\ : std_logic;
signal \N__66757\ : std_logic;
signal \N__66750\ : std_logic;
signal \N__66747\ : std_logic;
signal \N__66744\ : std_logic;
signal \N__66741\ : std_logic;
signal \N__66738\ : std_logic;
signal \N__66735\ : std_logic;
signal \N__66732\ : std_logic;
signal \N__66729\ : std_logic;
signal \N__66726\ : std_logic;
signal \N__66723\ : std_logic;
signal \N__66720\ : std_logic;
signal \N__66717\ : std_logic;
signal \N__66714\ : std_logic;
signal \N__66711\ : std_logic;
signal \N__66708\ : std_logic;
signal \N__66705\ : std_logic;
signal \N__66698\ : std_logic;
signal \N__66695\ : std_logic;
signal \N__66688\ : std_logic;
signal \N__66685\ : std_logic;
signal \N__66676\ : std_logic;
signal \N__66673\ : std_logic;
signal \N__66668\ : std_logic;
signal \N__66663\ : std_logic;
signal \N__66658\ : std_logic;
signal \N__66649\ : std_logic;
signal \N__66646\ : std_logic;
signal \N__66643\ : std_logic;
signal \N__66640\ : std_logic;
signal \N__66639\ : std_logic;
signal \N__66638\ : std_logic;
signal \N__66635\ : std_logic;
signal \N__66632\ : std_logic;
signal \N__66631\ : std_logic;
signal \N__66630\ : std_logic;
signal \N__66629\ : std_logic;
signal \N__66626\ : std_logic;
signal \N__66625\ : std_logic;
signal \N__66622\ : std_logic;
signal \N__66619\ : std_logic;
signal \N__66616\ : std_logic;
signal \N__66613\ : std_logic;
signal \N__66612\ : std_logic;
signal \N__66609\ : std_logic;
signal \N__66608\ : std_logic;
signal \N__66605\ : std_logic;
signal \N__66604\ : std_logic;
signal \N__66601\ : std_logic;
signal \N__66600\ : std_logic;
signal \N__66599\ : std_logic;
signal \N__66598\ : std_logic;
signal \N__66595\ : std_logic;
signal \N__66592\ : std_logic;
signal \N__66589\ : std_logic;
signal \N__66586\ : std_logic;
signal \N__66583\ : std_logic;
signal \N__66580\ : std_logic;
signal \N__66577\ : std_logic;
signal \N__66576\ : std_logic;
signal \N__66575\ : std_logic;
signal \N__66574\ : std_logic;
signal \N__66571\ : std_logic;
signal \N__66568\ : std_logic;
signal \N__66565\ : std_logic;
signal \N__66562\ : std_logic;
signal \N__66559\ : std_logic;
signal \N__66556\ : std_logic;
signal \N__66549\ : std_logic;
signal \N__66542\ : std_logic;
signal \N__66539\ : std_logic;
signal \N__66538\ : std_logic;
signal \N__66535\ : std_logic;
signal \N__66534\ : std_logic;
signal \N__66531\ : std_logic;
signal \N__66528\ : std_logic;
signal \N__66525\ : std_logic;
signal \N__66522\ : std_logic;
signal \N__66521\ : std_logic;
signal \N__66520\ : std_logic;
signal \N__66519\ : std_logic;
signal \N__66518\ : std_logic;
signal \N__66517\ : std_logic;
signal \N__66516\ : std_logic;
signal \N__66515\ : std_logic;
signal \N__66512\ : std_logic;
signal \N__66509\ : std_logic;
signal \N__66506\ : std_logic;
signal \N__66503\ : std_logic;
signal \N__66496\ : std_logic;
signal \N__66493\ : std_logic;
signal \N__66486\ : std_logic;
signal \N__66483\ : std_logic;
signal \N__66478\ : std_logic;
signal \N__66475\ : std_logic;
signal \N__66472\ : std_logic;
signal \N__66469\ : std_logic;
signal \N__66468\ : std_logic;
signal \N__66465\ : std_logic;
signal \N__66464\ : std_logic;
signal \N__66461\ : std_logic;
signal \N__66458\ : std_logic;
signal \N__66455\ : std_logic;
signal \N__66448\ : std_logic;
signal \N__66445\ : std_logic;
signal \N__66442\ : std_logic;
signal \N__66435\ : std_logic;
signal \N__66432\ : std_logic;
signal \N__66429\ : std_logic;
signal \N__66416\ : std_logic;
signal \N__66411\ : std_logic;
signal \N__66408\ : std_logic;
signal \N__66393\ : std_logic;
signal \N__66388\ : std_logic;
signal \N__66385\ : std_logic;
signal \N__66382\ : std_logic;
signal \N__66379\ : std_logic;
signal \N__66376\ : std_logic;
signal \N__66373\ : std_logic;
signal \N__66370\ : std_logic;
signal \N__66367\ : std_logic;
signal \N__66364\ : std_logic;
signal \N__66361\ : std_logic;
signal \N__66360\ : std_logic;
signal \N__66359\ : std_logic;
signal \N__66356\ : std_logic;
signal \N__66353\ : std_logic;
signal \N__66350\ : std_logic;
signal \N__66349\ : std_logic;
signal \N__66348\ : std_logic;
signal \N__66347\ : std_logic;
signal \N__66346\ : std_logic;
signal \N__66345\ : std_logic;
signal \N__66344\ : std_logic;
signal \N__66343\ : std_logic;
signal \N__66340\ : std_logic;
signal \N__66337\ : std_logic;
signal \N__66334\ : std_logic;
signal \N__66331\ : std_logic;
signal \N__66328\ : std_logic;
signal \N__66327\ : std_logic;
signal \N__66324\ : std_logic;
signal \N__66321\ : std_logic;
signal \N__66318\ : std_logic;
signal \N__66315\ : std_logic;
signal \N__66312\ : std_logic;
signal \N__66307\ : std_logic;
signal \N__66304\ : std_logic;
signal \N__66301\ : std_logic;
signal \N__66298\ : std_logic;
signal \N__66295\ : std_logic;
signal \N__66294\ : std_logic;
signal \N__66293\ : std_logic;
signal \N__66290\ : std_logic;
signal \N__66287\ : std_logic;
signal \N__66286\ : std_logic;
signal \N__66283\ : std_logic;
signal \N__66280\ : std_logic;
signal \N__66277\ : std_logic;
signal \N__66268\ : std_logic;
signal \N__66265\ : std_logic;
signal \N__66262\ : std_logic;
signal \N__66261\ : std_logic;
signal \N__66260\ : std_logic;
signal \N__66259\ : std_logic;
signal \N__66256\ : std_logic;
signal \N__66253\ : std_logic;
signal \N__66250\ : std_logic;
signal \N__66247\ : std_logic;
signal \N__66244\ : std_logic;
signal \N__66235\ : std_logic;
signal \N__66232\ : std_logic;
signal \N__66229\ : std_logic;
signal \N__66226\ : std_logic;
signal \N__66221\ : std_logic;
signal \N__66220\ : std_logic;
signal \N__66219\ : std_logic;
signal \N__66218\ : std_logic;
signal \N__66217\ : std_logic;
signal \N__66214\ : std_logic;
signal \N__66211\ : std_logic;
signal \N__66208\ : std_logic;
signal \N__66201\ : std_logic;
signal \N__66198\ : std_logic;
signal \N__66193\ : std_logic;
signal \N__66192\ : std_logic;
signal \N__66189\ : std_logic;
signal \N__66188\ : std_logic;
signal \N__66185\ : std_logic;
signal \N__66184\ : std_logic;
signal \N__66181\ : std_logic;
signal \N__66180\ : std_logic;
signal \N__66177\ : std_logic;
signal \N__66174\ : std_logic;
signal \N__66169\ : std_logic;
signal \N__66166\ : std_logic;
signal \N__66163\ : std_logic;
signal \N__66160\ : std_logic;
signal \N__66143\ : std_logic;
signal \N__66140\ : std_logic;
signal \N__66137\ : std_logic;
signal \N__66132\ : std_logic;
signal \N__66127\ : std_logic;
signal \N__66118\ : std_logic;
signal \N__66115\ : std_logic;
signal \N__66112\ : std_logic;
signal \N__66109\ : std_logic;
signal \N__66106\ : std_logic;
signal \N__66103\ : std_logic;
signal \N__66100\ : std_logic;
signal \N__66099\ : std_logic;
signal \N__66098\ : std_logic;
signal \N__66095\ : std_logic;
signal \N__66094\ : std_logic;
signal \N__66093\ : std_logic;
signal \N__66092\ : std_logic;
signal \N__66091\ : std_logic;
signal \N__66090\ : std_logic;
signal \N__66087\ : std_logic;
signal \N__66086\ : std_logic;
signal \N__66083\ : std_logic;
signal \N__66080\ : std_logic;
signal \N__66077\ : std_logic;
signal \N__66074\ : std_logic;
signal \N__66071\ : std_logic;
signal \N__66070\ : std_logic;
signal \N__66067\ : std_logic;
signal \N__66064\ : std_logic;
signal \N__66063\ : std_logic;
signal \N__66060\ : std_logic;
signal \N__66057\ : std_logic;
signal \N__66056\ : std_logic;
signal \N__66053\ : std_logic;
signal \N__66050\ : std_logic;
signal \N__66047\ : std_logic;
signal \N__66044\ : std_logic;
signal \N__66041\ : std_logic;
signal \N__66040\ : std_logic;
signal \N__66037\ : std_logic;
signal \N__66036\ : std_logic;
signal \N__66033\ : std_logic;
signal \N__66032\ : std_logic;
signal \N__66031\ : std_logic;
signal \N__66030\ : std_logic;
signal \N__66029\ : std_logic;
signal \N__66028\ : std_logic;
signal \N__66025\ : std_logic;
signal \N__66022\ : std_logic;
signal \N__66019\ : std_logic;
signal \N__66016\ : std_logic;
signal \N__66013\ : std_logic;
signal \N__66012\ : std_logic;
signal \N__66005\ : std_logic;
signal \N__66002\ : std_logic;
signal \N__65999\ : std_logic;
signal \N__65996\ : std_logic;
signal \N__65993\ : std_logic;
signal \N__65990\ : std_logic;
signal \N__65987\ : std_logic;
signal \N__65984\ : std_logic;
signal \N__65983\ : std_logic;
signal \N__65980\ : std_logic;
signal \N__65979\ : std_logic;
signal \N__65976\ : std_logic;
signal \N__65975\ : std_logic;
signal \N__65972\ : std_logic;
signal \N__65969\ : std_logic;
signal \N__65966\ : std_logic;
signal \N__65963\ : std_logic;
signal \N__65958\ : std_logic;
signal \N__65955\ : std_logic;
signal \N__65952\ : std_logic;
signal \N__65941\ : std_logic;
signal \N__65938\ : std_logic;
signal \N__65935\ : std_logic;
signal \N__65928\ : std_logic;
signal \N__65917\ : std_logic;
signal \N__65914\ : std_logic;
signal \N__65911\ : std_logic;
signal \N__65908\ : std_logic;
signal \N__65905\ : std_logic;
signal \N__65902\ : std_logic;
signal \N__65897\ : std_logic;
signal \N__65890\ : std_logic;
signal \N__65887\ : std_logic;
signal \N__65884\ : std_logic;
signal \N__65877\ : std_logic;
signal \N__65872\ : std_logic;
signal \N__65863\ : std_logic;
signal \N__65860\ : std_logic;
signal \N__65857\ : std_logic;
signal \N__65854\ : std_logic;
signal \N__65851\ : std_logic;
signal \N__65848\ : std_logic;
signal \N__65845\ : std_logic;
signal \N__65844\ : std_logic;
signal \N__65843\ : std_logic;
signal \N__65840\ : std_logic;
signal \N__65839\ : std_logic;
signal \N__65836\ : std_logic;
signal \N__65833\ : std_logic;
signal \N__65832\ : std_logic;
signal \N__65831\ : std_logic;
signal \N__65830\ : std_logic;
signal \N__65829\ : std_logic;
signal \N__65828\ : std_logic;
signal \N__65825\ : std_logic;
signal \N__65822\ : std_logic;
signal \N__65819\ : std_logic;
signal \N__65816\ : std_logic;
signal \N__65813\ : std_logic;
signal \N__65810\ : std_logic;
signal \N__65809\ : std_logic;
signal \N__65808\ : std_logic;
signal \N__65807\ : std_logic;
signal \N__65804\ : std_logic;
signal \N__65801\ : std_logic;
signal \N__65798\ : std_logic;
signal \N__65795\ : std_logic;
signal \N__65792\ : std_logic;
signal \N__65791\ : std_logic;
signal \N__65786\ : std_logic;
signal \N__65783\ : std_logic;
signal \N__65780\ : std_logic;
signal \N__65777\ : std_logic;
signal \N__65776\ : std_logic;
signal \N__65773\ : std_logic;
signal \N__65770\ : std_logic;
signal \N__65767\ : std_logic;
signal \N__65764\ : std_logic;
signal \N__65761\ : std_logic;
signal \N__65756\ : std_logic;
signal \N__65753\ : std_logic;
signal \N__65746\ : std_logic;
signal \N__65743\ : std_logic;
signal \N__65740\ : std_logic;
signal \N__65739\ : std_logic;
signal \N__65738\ : std_logic;
signal \N__65737\ : std_logic;
signal \N__65736\ : std_logic;
signal \N__65735\ : std_logic;
signal \N__65734\ : std_logic;
signal \N__65731\ : std_logic;
signal \N__65728\ : std_logic;
signal \N__65725\ : std_logic;
signal \N__65718\ : std_logic;
signal \N__65715\ : std_logic;
signal \N__65710\ : std_logic;
signal \N__65707\ : std_logic;
signal \N__65704\ : std_logic;
signal \N__65701\ : std_logic;
signal \N__65698\ : std_logic;
signal \N__65697\ : std_logic;
signal \N__65694\ : std_logic;
signal \N__65691\ : std_logic;
signal \N__65688\ : std_logic;
signal \N__65683\ : std_logic;
signal \N__65680\ : std_logic;
signal \N__65675\ : std_logic;
signal \N__65670\ : std_logic;
signal \N__65667\ : std_logic;
signal \N__65662\ : std_logic;
signal \N__65653\ : std_logic;
signal \N__65648\ : std_logic;
signal \N__65645\ : std_logic;
signal \N__65636\ : std_logic;
signal \N__65629\ : std_logic;
signal \N__65626\ : std_logic;
signal \N__65623\ : std_logic;
signal \N__65620\ : std_logic;
signal \N__65617\ : std_logic;
signal \N__65614\ : std_logic;
signal \N__65611\ : std_logic;
signal \N__65610\ : std_logic;
signal \N__65609\ : std_logic;
signal \N__65606\ : std_logic;
signal \N__65603\ : std_logic;
signal \N__65602\ : std_logic;
signal \N__65601\ : std_logic;
signal \N__65600\ : std_logic;
signal \N__65597\ : std_logic;
signal \N__65596\ : std_logic;
signal \N__65595\ : std_logic;
signal \N__65592\ : std_logic;
signal \N__65589\ : std_logic;
signal \N__65586\ : std_logic;
signal \N__65583\ : std_logic;
signal \N__65582\ : std_logic;
signal \N__65581\ : std_logic;
signal \N__65580\ : std_logic;
signal \N__65577\ : std_logic;
signal \N__65574\ : std_logic;
signal \N__65571\ : std_logic;
signal \N__65570\ : std_logic;
signal \N__65567\ : std_logic;
signal \N__65562\ : std_logic;
signal \N__65559\ : std_logic;
signal \N__65556\ : std_logic;
signal \N__65553\ : std_logic;
signal \N__65550\ : std_logic;
signal \N__65547\ : std_logic;
signal \N__65546\ : std_logic;
signal \N__65543\ : std_logic;
signal \N__65540\ : std_logic;
signal \N__65537\ : std_logic;
signal \N__65534\ : std_logic;
signal \N__65531\ : std_logic;
signal \N__65524\ : std_logic;
signal \N__65521\ : std_logic;
signal \N__65518\ : std_logic;
signal \N__65515\ : std_logic;
signal \N__65512\ : std_logic;
signal \N__65511\ : std_logic;
signal \N__65510\ : std_logic;
signal \N__65509\ : std_logic;
signal \N__65508\ : std_logic;
signal \N__65507\ : std_logic;
signal \N__65504\ : std_logic;
signal \N__65499\ : std_logic;
signal \N__65496\ : std_logic;
signal \N__65493\ : std_logic;
signal \N__65492\ : std_logic;
signal \N__65483\ : std_logic;
signal \N__65480\ : std_logic;
signal \N__65477\ : std_logic;
signal \N__65468\ : std_logic;
signal \N__65467\ : std_logic;
signal \N__65464\ : std_logic;
signal \N__65459\ : std_logic;
signal \N__65456\ : std_logic;
signal \N__65453\ : std_logic;
signal \N__65448\ : std_logic;
signal \N__65445\ : std_logic;
signal \N__65442\ : std_logic;
signal \N__65439\ : std_logic;
signal \N__65438\ : std_logic;
signal \N__65437\ : std_logic;
signal \N__65432\ : std_logic;
signal \N__65427\ : std_logic;
signal \N__65418\ : std_logic;
signal \N__65413\ : std_logic;
signal \N__65404\ : std_logic;
signal \N__65401\ : std_logic;
signal \N__65398\ : std_logic;
signal \N__65395\ : std_logic;
signal \N__65392\ : std_logic;
signal \N__65389\ : std_logic;
signal \N__65388\ : std_logic;
signal \N__65387\ : std_logic;
signal \N__65386\ : std_logic;
signal \N__65385\ : std_logic;
signal \N__65384\ : std_logic;
signal \N__65381\ : std_logic;
signal \N__65378\ : std_logic;
signal \N__65375\ : std_logic;
signal \N__65374\ : std_logic;
signal \N__65371\ : std_logic;
signal \N__65368\ : std_logic;
signal \N__65365\ : std_logic;
signal \N__65362\ : std_logic;
signal \N__65361\ : std_logic;
signal \N__65356\ : std_logic;
signal \N__65353\ : std_logic;
signal \N__65352\ : std_logic;
signal \N__65349\ : std_logic;
signal \N__65348\ : std_logic;
signal \N__65343\ : std_logic;
signal \N__65342\ : std_logic;
signal \N__65341\ : std_logic;
signal \N__65338\ : std_logic;
signal \N__65335\ : std_logic;
signal \N__65330\ : std_logic;
signal \N__65327\ : std_logic;
signal \N__65324\ : std_logic;
signal \N__65321\ : std_logic;
signal \N__65320\ : std_logic;
signal \N__65317\ : std_logic;
signal \N__65314\ : std_logic;
signal \N__65313\ : std_logic;
signal \N__65310\ : std_logic;
signal \N__65301\ : std_logic;
signal \N__65296\ : std_logic;
signal \N__65293\ : std_logic;
signal \N__65288\ : std_logic;
signal \N__65285\ : std_logic;
signal \N__65284\ : std_logic;
signal \N__65281\ : std_logic;
signal \N__65274\ : std_logic;
signal \N__65271\ : std_logic;
signal \N__65268\ : std_logic;
signal \N__65265\ : std_logic;
signal \N__65264\ : std_logic;
signal \N__65261\ : std_logic;
signal \N__65258\ : std_logic;
signal \N__65251\ : std_logic;
signal \N__65248\ : std_logic;
signal \N__65245\ : std_logic;
signal \N__65242\ : std_logic;
signal \N__65239\ : std_logic;
signal \N__65236\ : std_logic;
signal \N__65227\ : std_logic;
signal \N__65224\ : std_logic;
signal \N__65221\ : std_logic;
signal \N__65218\ : std_logic;
signal \N__65215\ : std_logic;
signal \N__65212\ : std_logic;
signal \N__65209\ : std_logic;
signal \N__65206\ : std_logic;
signal \N__65203\ : std_logic;
signal \N__65202\ : std_logic;
signal \N__65201\ : std_logic;
signal \N__65198\ : std_logic;
signal \N__65195\ : std_logic;
signal \N__65194\ : std_logic;
signal \N__65193\ : std_logic;
signal \N__65192\ : std_logic;
signal \N__65189\ : std_logic;
signal \N__65188\ : std_logic;
signal \N__65185\ : std_logic;
signal \N__65182\ : std_logic;
signal \N__65179\ : std_logic;
signal \N__65178\ : std_logic;
signal \N__65175\ : std_logic;
signal \N__65172\ : std_logic;
signal \N__65171\ : std_logic;
signal \N__65170\ : std_logic;
signal \N__65169\ : std_logic;
signal \N__65166\ : std_logic;
signal \N__65163\ : std_logic;
signal \N__65156\ : std_logic;
signal \N__65153\ : std_logic;
signal \N__65152\ : std_logic;
signal \N__65149\ : std_logic;
signal \N__65146\ : std_logic;
signal \N__65143\ : std_logic;
signal \N__65140\ : std_logic;
signal \N__65139\ : std_logic;
signal \N__65136\ : std_logic;
signal \N__65135\ : std_logic;
signal \N__65132\ : std_logic;
signal \N__65129\ : std_logic;
signal \N__65126\ : std_logic;
signal \N__65123\ : std_logic;
signal \N__65120\ : std_logic;
signal \N__65119\ : std_logic;
signal \N__65118\ : std_logic;
signal \N__65109\ : std_logic;
signal \N__65106\ : std_logic;
signal \N__65103\ : std_logic;
signal \N__65100\ : std_logic;
signal \N__65095\ : std_logic;
signal \N__65090\ : std_logic;
signal \N__65087\ : std_logic;
signal \N__65082\ : std_logic;
signal \N__65077\ : std_logic;
signal \N__65072\ : std_logic;
signal \N__65065\ : std_logic;
signal \N__65062\ : std_logic;
signal \N__65061\ : std_logic;
signal \N__65058\ : std_logic;
signal \N__65055\ : std_logic;
signal \N__65050\ : std_logic;
signal \N__65047\ : std_logic;
signal \N__65038\ : std_logic;
signal \N__65035\ : std_logic;
signal \N__65032\ : std_logic;
signal \N__65029\ : std_logic;
signal \N__65026\ : std_logic;
signal \N__65023\ : std_logic;
signal \N__65020\ : std_logic;
signal \N__65017\ : std_logic;
signal \N__65016\ : std_logic;
signal \N__65015\ : std_logic;
signal \N__65014\ : std_logic;
signal \N__65013\ : std_logic;
signal \N__65012\ : std_logic;
signal \N__65011\ : std_logic;
signal \N__65010\ : std_logic;
signal \N__65009\ : std_logic;
signal \N__65008\ : std_logic;
signal \N__65007\ : std_logic;
signal \N__65006\ : std_logic;
signal \N__65005\ : std_logic;
signal \N__65004\ : std_logic;
signal \N__65001\ : std_logic;
signal \N__64998\ : std_logic;
signal \N__64995\ : std_logic;
signal \N__64992\ : std_logic;
signal \N__64989\ : std_logic;
signal \N__64986\ : std_logic;
signal \N__64983\ : std_logic;
signal \N__64980\ : std_logic;
signal \N__64977\ : std_logic;
signal \N__64974\ : std_logic;
signal \N__64971\ : std_logic;
signal \N__64968\ : std_logic;
signal \N__64965\ : std_logic;
signal \N__64964\ : std_logic;
signal \N__64961\ : std_logic;
signal \N__64960\ : std_logic;
signal \N__64957\ : std_logic;
signal \N__64956\ : std_logic;
signal \N__64955\ : std_logic;
signal \N__64948\ : std_logic;
signal \N__64947\ : std_logic;
signal \N__64940\ : std_logic;
signal \N__64933\ : std_logic;
signal \N__64922\ : std_logic;
signal \N__64921\ : std_logic;
signal \N__64918\ : std_logic;
signal \N__64915\ : std_logic;
signal \N__64914\ : std_logic;
signal \N__64911\ : std_logic;
signal \N__64910\ : std_logic;
signal \N__64907\ : std_logic;
signal \N__64904\ : std_logic;
signal \N__64901\ : std_logic;
signal \N__64900\ : std_logic;
signal \N__64899\ : std_logic;
signal \N__64892\ : std_logic;
signal \N__64889\ : std_logic;
signal \N__64888\ : std_logic;
signal \N__64887\ : std_logic;
signal \N__64884\ : std_logic;
signal \N__64881\ : std_logic;
signal \N__64878\ : std_logic;
signal \N__64875\ : std_logic;
signal \N__64872\ : std_logic;
signal \N__64869\ : std_logic;
signal \N__64864\ : std_logic;
signal \N__64863\ : std_logic;
signal \N__64862\ : std_logic;
signal \N__64859\ : std_logic;
signal \N__64856\ : std_logic;
signal \N__64851\ : std_logic;
signal \N__64848\ : std_logic;
signal \N__64845\ : std_logic;
signal \N__64844\ : std_logic;
signal \N__64837\ : std_logic;
signal \N__64832\ : std_logic;
signal \N__64829\ : std_logic;
signal \N__64826\ : std_logic;
signal \N__64823\ : std_logic;
signal \N__64820\ : std_logic;
signal \N__64817\ : std_logic;
signal \N__64810\ : std_logic;
signal \N__64807\ : std_logic;
signal \N__64804\ : std_logic;
signal \N__64801\ : std_logic;
signal \N__64798\ : std_logic;
signal \N__64787\ : std_logic;
signal \N__64782\ : std_logic;
signal \N__64779\ : std_logic;
signal \N__64776\ : std_logic;
signal \N__64771\ : std_logic;
signal \N__64766\ : std_logic;
signal \N__64759\ : std_logic;
signal \N__64758\ : std_logic;
signal \N__64755\ : std_logic;
signal \N__64754\ : std_logic;
signal \N__64753\ : std_logic;
signal \N__64750\ : std_logic;
signal \N__64749\ : std_logic;
signal \N__64748\ : std_logic;
signal \N__64747\ : std_logic;
signal \N__64744\ : std_logic;
signal \N__64741\ : std_logic;
signal \N__64738\ : std_logic;
signal \N__64735\ : std_logic;
signal \N__64734\ : std_logic;
signal \N__64731\ : std_logic;
signal \N__64728\ : std_logic;
signal \N__64727\ : std_logic;
signal \N__64726\ : std_logic;
signal \N__64723\ : std_logic;
signal \N__64720\ : std_logic;
signal \N__64717\ : std_logic;
signal \N__64714\ : std_logic;
signal \N__64713\ : std_logic;
signal \N__64712\ : std_logic;
signal \N__64709\ : std_logic;
signal \N__64706\ : std_logic;
signal \N__64703\ : std_logic;
signal \N__64700\ : std_logic;
signal \N__64697\ : std_logic;
signal \N__64694\ : std_logic;
signal \N__64693\ : std_logic;
signal \N__64690\ : std_logic;
signal \N__64683\ : std_logic;
signal \N__64680\ : std_logic;
signal \N__64677\ : std_logic;
signal \N__64674\ : std_logic;
signal \N__64671\ : std_logic;
signal \N__64666\ : std_logic;
signal \N__64663\ : std_logic;
signal \N__64660\ : std_logic;
signal \N__64657\ : std_logic;
signal \N__64648\ : std_logic;
signal \N__64647\ : std_logic;
signal \N__64646\ : std_logic;
signal \N__64645\ : std_logic;
signal \N__64644\ : std_logic;
signal \N__64643\ : std_logic;
signal \N__64642\ : std_logic;
signal \N__64641\ : std_logic;
signal \N__64640\ : std_logic;
signal \N__64639\ : std_logic;
signal \N__64638\ : std_logic;
signal \N__64633\ : std_logic;
signal \N__64632\ : std_logic;
signal \N__64625\ : std_logic;
signal \N__64622\ : std_logic;
signal \N__64619\ : std_logic;
signal \N__64616\ : std_logic;
signal \N__64613\ : std_logic;
signal \N__64612\ : std_logic;
signal \N__64609\ : std_logic;
signal \N__64606\ : std_logic;
signal \N__64603\ : std_logic;
signal \N__64600\ : std_logic;
signal \N__64599\ : std_logic;
signal \N__64596\ : std_logic;
signal \N__64593\ : std_logic;
signal \N__64592\ : std_logic;
signal \N__64589\ : std_logic;
signal \N__64588\ : std_logic;
signal \N__64585\ : std_logic;
signal \N__64582\ : std_logic;
signal \N__64579\ : std_logic;
signal \N__64576\ : std_logic;
signal \N__64573\ : std_logic;
signal \N__64570\ : std_logic;
signal \N__64565\ : std_logic;
signal \N__64556\ : std_logic;
signal \N__64549\ : std_logic;
signal \N__64538\ : std_logic;
signal \N__64533\ : std_logic;
signal \N__64528\ : std_logic;
signal \N__64519\ : std_logic;
signal \N__64516\ : std_logic;
signal \N__64507\ : std_logic;
signal \N__64504\ : std_logic;
signal \N__64501\ : std_logic;
signal \N__64498\ : std_logic;
signal \N__64497\ : std_logic;
signal \N__64496\ : std_logic;
signal \N__64493\ : std_logic;
signal \N__64490\ : std_logic;
signal \N__64489\ : std_logic;
signal \N__64488\ : std_logic;
signal \N__64485\ : std_logic;
signal \N__64482\ : std_logic;
signal \N__64479\ : std_logic;
signal \N__64478\ : std_logic;
signal \N__64475\ : std_logic;
signal \N__64472\ : std_logic;
signal \N__64471\ : std_logic;
signal \N__64470\ : std_logic;
signal \N__64467\ : std_logic;
signal \N__64466\ : std_logic;
signal \N__64461\ : std_logic;
signal \N__64458\ : std_logic;
signal \N__64455\ : std_logic;
signal \N__64454\ : std_logic;
signal \N__64453\ : std_logic;
signal \N__64452\ : std_logic;
signal \N__64451\ : std_logic;
signal \N__64450\ : std_logic;
signal \N__64447\ : std_logic;
signal \N__64444\ : std_logic;
signal \N__64441\ : std_logic;
signal \N__64440\ : std_logic;
signal \N__64439\ : std_logic;
signal \N__64438\ : std_logic;
signal \N__64437\ : std_logic;
signal \N__64434\ : std_logic;
signal \N__64431\ : std_logic;
signal \N__64426\ : std_logic;
signal \N__64423\ : std_logic;
signal \N__64420\ : std_logic;
signal \N__64417\ : std_logic;
signal \N__64414\ : std_logic;
signal \N__64411\ : std_logic;
signal \N__64408\ : std_logic;
signal \N__64403\ : std_logic;
signal \N__64400\ : std_logic;
signal \N__64397\ : std_logic;
signal \N__64396\ : std_logic;
signal \N__64393\ : std_logic;
signal \N__64392\ : std_logic;
signal \N__64389\ : std_logic;
signal \N__64388\ : std_logic;
signal \N__64385\ : std_logic;
signal \N__64384\ : std_logic;
signal \N__64383\ : std_logic;
signal \N__64382\ : std_logic;
signal \N__64381\ : std_logic;
signal \N__64378\ : std_logic;
signal \N__64375\ : std_logic;
signal \N__64368\ : std_logic;
signal \N__64365\ : std_logic;
signal \N__64362\ : std_logic;
signal \N__64359\ : std_logic;
signal \N__64356\ : std_logic;
signal \N__64349\ : std_logic;
signal \N__64336\ : std_logic;
signal \N__64335\ : std_logic;
signal \N__64332\ : std_logic;
signal \N__64331\ : std_logic;
signal \N__64328\ : std_logic;
signal \N__64327\ : std_logic;
signal \N__64324\ : std_logic;
signal \N__64323\ : std_logic;
signal \N__64320\ : std_logic;
signal \N__64315\ : std_logic;
signal \N__64308\ : std_logic;
signal \N__64303\ : std_logic;
signal \N__64298\ : std_logic;
signal \N__64281\ : std_logic;
signal \N__64278\ : std_logic;
signal \N__64275\ : std_logic;
signal \N__64268\ : std_logic;
signal \N__64261\ : std_logic;
signal \N__64258\ : std_logic;
signal \N__64255\ : std_logic;
signal \N__64252\ : std_logic;
signal \N__64249\ : std_logic;
signal \N__64246\ : std_logic;
signal \N__64243\ : std_logic;
signal \N__64242\ : std_logic;
signal \N__64241\ : std_logic;
signal \N__64240\ : std_logic;
signal \N__64239\ : std_logic;
signal \N__64238\ : std_logic;
signal \N__64237\ : std_logic;
signal \N__64236\ : std_logic;
signal \N__64235\ : std_logic;
signal \N__64234\ : std_logic;
signal \N__64233\ : std_logic;
signal \N__64232\ : std_logic;
signal \N__64231\ : std_logic;
signal \N__64230\ : std_logic;
signal \N__64227\ : std_logic;
signal \N__64224\ : std_logic;
signal \N__64221\ : std_logic;
signal \N__64220\ : std_logic;
signal \N__64219\ : std_logic;
signal \N__64216\ : std_logic;
signal \N__64215\ : std_logic;
signal \N__64212\ : std_logic;
signal \N__64211\ : std_logic;
signal \N__64208\ : std_logic;
signal \N__64207\ : std_logic;
signal \N__64204\ : std_logic;
signal \N__64201\ : std_logic;
signal \N__64200\ : std_logic;
signal \N__64197\ : std_logic;
signal \N__64196\ : std_logic;
signal \N__64193\ : std_logic;
signal \N__64192\ : std_logic;
signal \N__64189\ : std_logic;
signal \N__64186\ : std_logic;
signal \N__64183\ : std_logic;
signal \N__64182\ : std_logic;
signal \N__64179\ : std_logic;
signal \N__64178\ : std_logic;
signal \N__64175\ : std_logic;
signal \N__64172\ : std_logic;
signal \N__64169\ : std_logic;
signal \N__64166\ : std_logic;
signal \N__64149\ : std_logic;
signal \N__64146\ : std_logic;
signal \N__64133\ : std_logic;
signal \N__64132\ : std_logic;
signal \N__64129\ : std_logic;
signal \N__64126\ : std_logic;
signal \N__64123\ : std_logic;
signal \N__64120\ : std_logic;
signal \N__64117\ : std_logic;
signal \N__64112\ : std_logic;
signal \N__64111\ : std_logic;
signal \N__64108\ : std_logic;
signal \N__64105\ : std_logic;
signal \N__64102\ : std_logic;
signal \N__64101\ : std_logic;
signal \N__64098\ : std_logic;
signal \N__64095\ : std_logic;
signal \N__64092\ : std_logic;
signal \N__64091\ : std_logic;
signal \N__64090\ : std_logic;
signal \N__64081\ : std_logic;
signal \N__64078\ : std_logic;
signal \N__64075\ : std_logic;
signal \N__64072\ : std_logic;
signal \N__64067\ : std_logic;
signal \N__64064\ : std_logic;
signal \N__64061\ : std_logic;
signal \N__64054\ : std_logic;
signal \N__64051\ : std_logic;
signal \N__64048\ : std_logic;
signal \N__64043\ : std_logic;
signal \N__64038\ : std_logic;
signal \N__64031\ : std_logic;
signal \N__64026\ : std_logic;
signal \N__64023\ : std_logic;
signal \N__64020\ : std_logic;
signal \N__64017\ : std_logic;
signal \N__64014\ : std_logic;
signal \N__64009\ : std_logic;
signal \N__64000\ : std_logic;
signal \N__63997\ : std_logic;
signal \N__63994\ : std_logic;
signal \N__63991\ : std_logic;
signal \N__63988\ : std_logic;
signal \N__63985\ : std_logic;
signal \N__63982\ : std_logic;
signal \N__63981\ : std_logic;
signal \N__63980\ : std_logic;
signal \N__63979\ : std_logic;
signal \N__63976\ : std_logic;
signal \N__63975\ : std_logic;
signal \N__63974\ : std_logic;
signal \N__63971\ : std_logic;
signal \N__63968\ : std_logic;
signal \N__63967\ : std_logic;
signal \N__63964\ : std_logic;
signal \N__63963\ : std_logic;
signal \N__63962\ : std_logic;
signal \N__63959\ : std_logic;
signal \N__63956\ : std_logic;
signal \N__63955\ : std_logic;
signal \N__63952\ : std_logic;
signal \N__63951\ : std_logic;
signal \N__63950\ : std_logic;
signal \N__63949\ : std_logic;
signal \N__63948\ : std_logic;
signal \N__63947\ : std_logic;
signal \N__63946\ : std_logic;
signal \N__63943\ : std_logic;
signal \N__63940\ : std_logic;
signal \N__63937\ : std_logic;
signal \N__63936\ : std_logic;
signal \N__63933\ : std_logic;
signal \N__63930\ : std_logic;
signal \N__63929\ : std_logic;
signal \N__63926\ : std_logic;
signal \N__63921\ : std_logic;
signal \N__63918\ : std_logic;
signal \N__63915\ : std_logic;
signal \N__63912\ : std_logic;
signal \N__63909\ : std_logic;
signal \N__63906\ : std_logic;
signal \N__63903\ : std_logic;
signal \N__63900\ : std_logic;
signal \N__63897\ : std_logic;
signal \N__63896\ : std_logic;
signal \N__63895\ : std_logic;
signal \N__63894\ : std_logic;
signal \N__63893\ : std_logic;
signal \N__63892\ : std_logic;
signal \N__63891\ : std_logic;
signal \N__63890\ : std_logic;
signal \N__63889\ : std_logic;
signal \N__63888\ : std_logic;
signal \N__63885\ : std_logic;
signal \N__63882\ : std_logic;
signal \N__63879\ : std_logic;
signal \N__63876\ : std_logic;
signal \N__63875\ : std_logic;
signal \N__63872\ : std_logic;
signal \N__63869\ : std_logic;
signal \N__63866\ : std_logic;
signal \N__63863\ : std_logic;
signal \N__63862\ : std_logic;
signal \N__63859\ : std_logic;
signal \N__63856\ : std_logic;
signal \N__63853\ : std_logic;
signal \N__63846\ : std_logic;
signal \N__63839\ : std_logic;
signal \N__63836\ : std_logic;
signal \N__63833\ : std_logic;
signal \N__63830\ : std_logic;
signal \N__63827\ : std_logic;
signal \N__63824\ : std_logic;
signal \N__63821\ : std_logic;
signal \N__63818\ : std_logic;
signal \N__63815\ : std_logic;
signal \N__63812\ : std_logic;
signal \N__63805\ : std_logic;
signal \N__63802\ : std_logic;
signal \N__63799\ : std_logic;
signal \N__63794\ : std_logic;
signal \N__63791\ : std_logic;
signal \N__63788\ : std_logic;
signal \N__63785\ : std_logic;
signal \N__63780\ : std_logic;
signal \N__63777\ : std_logic;
signal \N__63772\ : std_logic;
signal \N__63763\ : std_logic;
signal \N__63754\ : std_logic;
signal \N__63751\ : std_logic;
signal \N__63746\ : std_logic;
signal \N__63739\ : std_logic;
signal \N__63734\ : std_logic;
signal \N__63731\ : std_logic;
signal \N__63720\ : std_logic;
signal \N__63715\ : std_logic;
signal \N__63706\ : std_logic;
signal \N__63703\ : std_logic;
signal \N__63700\ : std_logic;
signal \N__63697\ : std_logic;
signal \N__63694\ : std_logic;
signal \N__63691\ : std_logic;
signal \N__63688\ : std_logic;
signal \N__63687\ : std_logic;
signal \N__63686\ : std_logic;
signal \N__63683\ : std_logic;
signal \N__63682\ : std_logic;
signal \N__63679\ : std_logic;
signal \N__63676\ : std_logic;
signal \N__63673\ : std_logic;
signal \N__63670\ : std_logic;
signal \N__63669\ : std_logic;
signal \N__63668\ : std_logic;
signal \N__63665\ : std_logic;
signal \N__63662\ : std_logic;
signal \N__63659\ : std_logic;
signal \N__63656\ : std_logic;
signal \N__63655\ : std_logic;
signal \N__63652\ : std_logic;
signal \N__63649\ : std_logic;
signal \N__63648\ : std_logic;
signal \N__63647\ : std_logic;
signal \N__63644\ : std_logic;
signal \N__63641\ : std_logic;
signal \N__63636\ : std_logic;
signal \N__63635\ : std_logic;
signal \N__63634\ : std_logic;
signal \N__63633\ : std_logic;
signal \N__63632\ : std_logic;
signal \N__63631\ : std_logic;
signal \N__63630\ : std_logic;
signal \N__63627\ : std_logic;
signal \N__63626\ : std_logic;
signal \N__63625\ : std_logic;
signal \N__63624\ : std_logic;
signal \N__63623\ : std_logic;
signal \N__63622\ : std_logic;
signal \N__63619\ : std_logic;
signal \N__63616\ : std_logic;
signal \N__63613\ : std_logic;
signal \N__63610\ : std_logic;
signal \N__63609\ : std_logic;
signal \N__63608\ : std_logic;
signal \N__63607\ : std_logic;
signal \N__63600\ : std_logic;
signal \N__63599\ : std_logic;
signal \N__63596\ : std_logic;
signal \N__63595\ : std_logic;
signal \N__63592\ : std_logic;
signal \N__63591\ : std_logic;
signal \N__63588\ : std_logic;
signal \N__63587\ : std_logic;
signal \N__63584\ : std_logic;
signal \N__63581\ : std_logic;
signal \N__63578\ : std_logic;
signal \N__63575\ : std_logic;
signal \N__63572\ : std_logic;
signal \N__63569\ : std_logic;
signal \N__63566\ : std_logic;
signal \N__63565\ : std_logic;
signal \N__63562\ : std_logic;
signal \N__63561\ : std_logic;
signal \N__63558\ : std_logic;
signal \N__63553\ : std_logic;
signal \N__63550\ : std_logic;
signal \N__63547\ : std_logic;
signal \N__63544\ : std_logic;
signal \N__63541\ : std_logic;
signal \N__63538\ : std_logic;
signal \N__63535\ : std_logic;
signal \N__63518\ : std_logic;
signal \N__63515\ : std_logic;
signal \N__63510\ : std_logic;
signal \N__63507\ : std_logic;
signal \N__63504\ : std_logic;
signal \N__63493\ : std_logic;
signal \N__63488\ : std_logic;
signal \N__63485\ : std_logic;
signal \N__63482\ : std_logic;
signal \N__63479\ : std_logic;
signal \N__63472\ : std_logic;
signal \N__63469\ : std_logic;
signal \N__63464\ : std_logic;
signal \N__63457\ : std_logic;
signal \N__63454\ : std_logic;
signal \N__63451\ : std_logic;
signal \N__63448\ : std_logic;
signal \N__63443\ : std_logic;
signal \N__63438\ : std_logic;
signal \N__63433\ : std_logic;
signal \N__63424\ : std_logic;
signal \N__63421\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63415\ : std_logic;
signal \N__63412\ : std_logic;
signal \N__63409\ : std_logic;
signal \N__63406\ : std_logic;
signal \N__63405\ : std_logic;
signal \N__63402\ : std_logic;
signal \N__63401\ : std_logic;
signal \N__63400\ : std_logic;
signal \N__63399\ : std_logic;
signal \N__63396\ : std_logic;
signal \N__63393\ : std_logic;
signal \N__63390\ : std_logic;
signal \N__63389\ : std_logic;
signal \N__63386\ : std_logic;
signal \N__63385\ : std_logic;
signal \N__63384\ : std_logic;
signal \N__63383\ : std_logic;
signal \N__63382\ : std_logic;
signal \N__63379\ : std_logic;
signal \N__63378\ : std_logic;
signal \N__63377\ : std_logic;
signal \N__63374\ : std_logic;
signal \N__63371\ : std_logic;
signal \N__63368\ : std_logic;
signal \N__63365\ : std_logic;
signal \N__63362\ : std_logic;
signal \N__63361\ : std_logic;
signal \N__63360\ : std_logic;
signal \N__63359\ : std_logic;
signal \N__63358\ : std_logic;
signal \N__63355\ : std_logic;
signal \N__63352\ : std_logic;
signal \N__63349\ : std_logic;
signal \N__63346\ : std_logic;
signal \N__63343\ : std_logic;
signal \N__63340\ : std_logic;
signal \N__63337\ : std_logic;
signal \N__63336\ : std_logic;
signal \N__63329\ : std_logic;
signal \N__63326\ : std_logic;
signal \N__63323\ : std_logic;
signal \N__63320\ : std_logic;
signal \N__63319\ : std_logic;
signal \N__63316\ : std_logic;
signal \N__63315\ : std_logic;
signal \N__63312\ : std_logic;
signal \N__63311\ : std_logic;
signal \N__63308\ : std_logic;
signal \N__63305\ : std_logic;
signal \N__63302\ : std_logic;
signal \N__63299\ : std_logic;
signal \N__63296\ : std_logic;
signal \N__63293\ : std_logic;
signal \N__63290\ : std_logic;
signal \N__63287\ : std_logic;
signal \N__63286\ : std_logic;
signal \N__63285\ : std_logic;
signal \N__63284\ : std_logic;
signal \N__63281\ : std_logic;
signal \N__63280\ : std_logic;
signal \N__63279\ : std_logic;
signal \N__63274\ : std_logic;
signal \N__63271\ : std_logic;
signal \N__63268\ : std_logic;
signal \N__63255\ : std_logic;
signal \N__63252\ : std_logic;
signal \N__63247\ : std_logic;
signal \N__63238\ : std_logic;
signal \N__63237\ : std_logic;
signal \N__63234\ : std_logic;
signal \N__63233\ : std_logic;
signal \N__63230\ : std_logic;
signal \N__63229\ : std_logic;
signal \N__63226\ : std_logic;
signal \N__63221\ : std_logic;
signal \N__63218\ : std_logic;
signal \N__63215\ : std_logic;
signal \N__63210\ : std_logic;
signal \N__63207\ : std_logic;
signal \N__63200\ : std_logic;
signal \N__63187\ : std_logic;
signal \N__63184\ : std_logic;
signal \N__63181\ : std_logic;
signal \N__63180\ : std_logic;
signal \N__63177\ : std_logic;
signal \N__63174\ : std_logic;
signal \N__63167\ : std_logic;
signal \N__63162\ : std_logic;
signal \N__63159\ : std_logic;
signal \N__63148\ : std_logic;
signal \N__63145\ : std_logic;
signal \N__63142\ : std_logic;
signal \N__63139\ : std_logic;
signal \N__63136\ : std_logic;
signal \N__63135\ : std_logic;
signal \N__63134\ : std_logic;
signal \N__63133\ : std_logic;
signal \N__63132\ : std_logic;
signal \N__63131\ : std_logic;
signal \N__63128\ : std_logic;
signal \N__63127\ : std_logic;
signal \N__63124\ : std_logic;
signal \N__63121\ : std_logic;
signal \N__63118\ : std_logic;
signal \N__63115\ : std_logic;
signal \N__63114\ : std_logic;
signal \N__63113\ : std_logic;
signal \N__63112\ : std_logic;
signal \N__63111\ : std_logic;
signal \N__63110\ : std_logic;
signal \N__63109\ : std_logic;
signal \N__63106\ : std_logic;
signal \N__63103\ : std_logic;
signal \N__63100\ : std_logic;
signal \N__63099\ : std_logic;
signal \N__63098\ : std_logic;
signal \N__63097\ : std_logic;
signal \N__63096\ : std_logic;
signal \N__63095\ : std_logic;
signal \N__63094\ : std_logic;
signal \N__63093\ : std_logic;
signal \N__63084\ : std_logic;
signal \N__63081\ : std_logic;
signal \N__63078\ : std_logic;
signal \N__63075\ : std_logic;
signal \N__63072\ : std_logic;
signal \N__63069\ : std_logic;
signal \N__63066\ : std_logic;
signal \N__63065\ : std_logic;
signal \N__63062\ : std_logic;
signal \N__63059\ : std_logic;
signal \N__63056\ : std_logic;
signal \N__63053\ : std_logic;
signal \N__63052\ : std_logic;
signal \N__63049\ : std_logic;
signal \N__63048\ : std_logic;
signal \N__63045\ : std_logic;
signal \N__63044\ : std_logic;
signal \N__63041\ : std_logic;
signal \N__63038\ : std_logic;
signal \N__63035\ : std_logic;
signal \N__63032\ : std_logic;
signal \N__63031\ : std_logic;
signal \N__63028\ : std_logic;
signal \N__63019\ : std_logic;
signal \N__63016\ : std_logic;
signal \N__63013\ : std_logic;
signal \N__63010\ : std_logic;
signal \N__63003\ : std_logic;
signal \N__63000\ : std_logic;
signal \N__62999\ : std_logic;
signal \N__62986\ : std_logic;
signal \N__62983\ : std_logic;
signal \N__62978\ : std_logic;
signal \N__62975\ : std_logic;
signal \N__62974\ : std_logic;
signal \N__62971\ : std_logic;
signal \N__62968\ : std_logic;
signal \N__62963\ : std_logic;
signal \N__62960\ : std_logic;
signal \N__62959\ : std_logic;
signal \N__62954\ : std_logic;
signal \N__62951\ : std_logic;
signal \N__62948\ : std_logic;
signal \N__62945\ : std_logic;
signal \N__62942\ : std_logic;
signal \N__62939\ : std_logic;
signal \N__62938\ : std_logic;
signal \N__62935\ : std_logic;
signal \N__62930\ : std_logic;
signal \N__62925\ : std_logic;
signal \N__62922\ : std_logic;
signal \N__62919\ : std_logic;
signal \N__62916\ : std_logic;
signal \N__62913\ : std_logic;
signal \N__62906\ : std_logic;
signal \N__62903\ : std_logic;
signal \N__62900\ : std_logic;
signal \N__62895\ : std_logic;
signal \N__62892\ : std_logic;
signal \N__62887\ : std_logic;
signal \N__62882\ : std_logic;
signal \N__62879\ : std_logic;
signal \N__62872\ : std_logic;
signal \N__62869\ : std_logic;
signal \N__62866\ : std_logic;
signal \N__62861\ : std_logic;
signal \N__62854\ : std_logic;
signal \N__62851\ : std_logic;
signal \N__62848\ : std_logic;
signal \N__62845\ : std_logic;
signal \N__62842\ : std_logic;
signal \N__62839\ : std_logic;
signal \N__62836\ : std_logic;
signal \N__62833\ : std_logic;
signal \N__62830\ : std_logic;
signal \N__62827\ : std_logic;
signal \N__62824\ : std_logic;
signal \N__62821\ : std_logic;
signal \N__62818\ : std_logic;
signal \N__62815\ : std_logic;
signal \N__62812\ : std_logic;
signal \N__62809\ : std_logic;
signal \N__62806\ : std_logic;
signal \N__62803\ : std_logic;
signal \N__62800\ : std_logic;
signal \N__62797\ : std_logic;
signal \N__62794\ : std_logic;
signal \N__62791\ : std_logic;
signal \N__62788\ : std_logic;
signal \N__62785\ : std_logic;
signal \N__62782\ : std_logic;
signal \N__62779\ : std_logic;
signal \N__62776\ : std_logic;
signal \N__62773\ : std_logic;
signal \N__62770\ : std_logic;
signal \N__62767\ : std_logic;
signal \N__62764\ : std_logic;
signal \N__62761\ : std_logic;
signal \N__62758\ : std_logic;
signal \N__62755\ : std_logic;
signal \N__62752\ : std_logic;
signal \N__62749\ : std_logic;
signal \N__62746\ : std_logic;
signal \N__62743\ : std_logic;
signal \N__62740\ : std_logic;
signal \N__62737\ : std_logic;
signal \N__62734\ : std_logic;
signal \N__62731\ : std_logic;
signal \N__62728\ : std_logic;
signal \N__62725\ : std_logic;
signal \N__62722\ : std_logic;
signal \N__62721\ : std_logic;
signal \N__62718\ : std_logic;
signal \N__62715\ : std_logic;
signal \N__62714\ : std_logic;
signal \N__62711\ : std_logic;
signal \N__62708\ : std_logic;
signal \N__62705\ : std_logic;
signal \N__62698\ : std_logic;
signal \N__62697\ : std_logic;
signal \N__62694\ : std_logic;
signal \N__62691\ : std_logic;
signal \N__62688\ : std_logic;
signal \N__62687\ : std_logic;
signal \N__62684\ : std_logic;
signal \N__62681\ : std_logic;
signal \N__62678\ : std_logic;
signal \N__62671\ : std_logic;
signal \N__62668\ : std_logic;
signal \N__62667\ : std_logic;
signal \N__62664\ : std_logic;
signal \N__62661\ : std_logic;
signal \N__62660\ : std_logic;
signal \N__62655\ : std_logic;
signal \N__62652\ : std_logic;
signal \N__62647\ : std_logic;
signal \N__62644\ : std_logic;
signal \N__62641\ : std_logic;
signal \N__62638\ : std_logic;
signal \N__62635\ : std_logic;
signal \N__62632\ : std_logic;
signal \N__62629\ : std_logic;
signal \N__62626\ : std_logic;
signal \N__62623\ : std_logic;
signal \N__62620\ : std_logic;
signal \N__62617\ : std_logic;
signal \N__62614\ : std_logic;
signal \N__62611\ : std_logic;
signal \N__62608\ : std_logic;
signal \N__62605\ : std_logic;
signal \N__62602\ : std_logic;
signal \N__62599\ : std_logic;
signal \N__62596\ : std_logic;
signal \N__62593\ : std_logic;
signal \N__62590\ : std_logic;
signal \N__62587\ : std_logic;
signal \N__62584\ : std_logic;
signal \N__62581\ : std_logic;
signal \N__62578\ : std_logic;
signal \N__62575\ : std_logic;
signal \N__62572\ : std_logic;
signal \N__62569\ : std_logic;
signal \N__62566\ : std_logic;
signal \N__62565\ : std_logic;
signal \N__62564\ : std_logic;
signal \N__62561\ : std_logic;
signal \N__62556\ : std_logic;
signal \N__62551\ : std_logic;
signal \N__62548\ : std_logic;
signal \N__62547\ : std_logic;
signal \N__62544\ : std_logic;
signal \N__62541\ : std_logic;
signal \N__62536\ : std_logic;
signal \N__62535\ : std_logic;
signal \N__62534\ : std_logic;
signal \N__62531\ : std_logic;
signal \N__62528\ : std_logic;
signal \N__62525\ : std_logic;
signal \N__62518\ : std_logic;
signal \N__62517\ : std_logic;
signal \N__62516\ : std_logic;
signal \N__62513\ : std_logic;
signal \N__62510\ : std_logic;
signal \N__62507\ : std_logic;
signal \N__62504\ : std_logic;
signal \N__62501\ : std_logic;
signal \N__62494\ : std_logic;
signal \N__62491\ : std_logic;
signal \N__62490\ : std_logic;
signal \N__62487\ : std_logic;
signal \N__62484\ : std_logic;
signal \N__62483\ : std_logic;
signal \N__62480\ : std_logic;
signal \N__62477\ : std_logic;
signal \N__62474\ : std_logic;
signal \N__62467\ : std_logic;
signal \N__62464\ : std_logic;
signal \N__62461\ : std_logic;
signal \N__62460\ : std_logic;
signal \N__62459\ : std_logic;
signal \N__62456\ : std_logic;
signal \N__62453\ : std_logic;
signal \N__62450\ : std_logic;
signal \N__62443\ : std_logic;
signal \N__62440\ : std_logic;
signal \N__62437\ : std_logic;
signal \N__62436\ : std_logic;
signal \N__62435\ : std_logic;
signal \N__62432\ : std_logic;
signal \N__62429\ : std_logic;
signal \N__62426\ : std_logic;
signal \N__62419\ : std_logic;
signal \N__62416\ : std_logic;
signal \N__62415\ : std_logic;
signal \N__62412\ : std_logic;
signal \N__62411\ : std_logic;
signal \N__62408\ : std_logic;
signal \N__62405\ : std_logic;
signal \N__62402\ : std_logic;
signal \N__62395\ : std_logic;
signal \N__62392\ : std_logic;
signal \N__62389\ : std_logic;
signal \N__62388\ : std_logic;
signal \N__62387\ : std_logic;
signal \N__62384\ : std_logic;
signal \N__62381\ : std_logic;
signal \N__62378\ : std_logic;
signal \N__62371\ : std_logic;
signal \N__62368\ : std_logic;
signal \N__62367\ : std_logic;
signal \N__62366\ : std_logic;
signal \N__62363\ : std_logic;
signal \N__62360\ : std_logic;
signal \N__62357\ : std_logic;
signal \N__62350\ : std_logic;
signal \N__62347\ : std_logic;
signal \N__62344\ : std_logic;
signal \N__62341\ : std_logic;
signal \N__62340\ : std_logic;
signal \N__62339\ : std_logic;
signal \N__62336\ : std_logic;
signal \N__62333\ : std_logic;
signal \N__62330\ : std_logic;
signal \N__62323\ : std_logic;
signal \N__62320\ : std_logic;
signal \N__62317\ : std_logic;
signal \N__62314\ : std_logic;
signal \N__62311\ : std_logic;
signal \N__62308\ : std_logic;
signal \N__62307\ : std_logic;
signal \N__62304\ : std_logic;
signal \N__62301\ : std_logic;
signal \N__62300\ : std_logic;
signal \N__62297\ : std_logic;
signal \N__62294\ : std_logic;
signal \N__62291\ : std_logic;
signal \N__62284\ : std_logic;
signal \N__62283\ : std_logic;
signal \N__62280\ : std_logic;
signal \N__62279\ : std_logic;
signal \N__62276\ : std_logic;
signal \N__62273\ : std_logic;
signal \N__62270\ : std_logic;
signal \N__62267\ : std_logic;
signal \N__62264\ : std_logic;
signal \N__62261\ : std_logic;
signal \N__62254\ : std_logic;
signal \N__62251\ : std_logic;
signal \N__62250\ : std_logic;
signal \N__62247\ : std_logic;
signal \N__62244\ : std_logic;
signal \N__62243\ : std_logic;
signal \N__62238\ : std_logic;
signal \N__62235\ : std_logic;
signal \N__62230\ : std_logic;
signal \N__62227\ : std_logic;
signal \N__62226\ : std_logic;
signal \N__62223\ : std_logic;
signal \N__62220\ : std_logic;
signal \N__62215\ : std_logic;
signal \N__62214\ : std_logic;
signal \N__62211\ : std_logic;
signal \N__62208\ : std_logic;
signal \N__62203\ : std_logic;
signal \N__62202\ : std_logic;
signal \N__62199\ : std_logic;
signal \N__62196\ : std_logic;
signal \N__62191\ : std_logic;
signal \N__62190\ : std_logic;
signal \N__62187\ : std_logic;
signal \N__62184\ : std_logic;
signal \N__62179\ : std_logic;
signal \N__62176\ : std_logic;
signal \N__62175\ : std_logic;
signal \N__62172\ : std_logic;
signal \N__62169\ : std_logic;
signal \N__62166\ : std_logic;
signal \N__62165\ : std_logic;
signal \N__62160\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62152\ : std_logic;
signal \N__62149\ : std_logic;
signal \N__62146\ : std_logic;
signal \N__62143\ : std_logic;
signal \N__62142\ : std_logic;
signal \N__62139\ : std_logic;
signal \N__62136\ : std_logic;
signal \N__62131\ : std_logic;
signal \N__62130\ : std_logic;
signal \N__62127\ : std_logic;
signal \N__62124\ : std_logic;
signal \N__62119\ : std_logic;
signal \N__62118\ : std_logic;
signal \N__62117\ : std_logic;
signal \N__62116\ : std_logic;
signal \N__62115\ : std_logic;
signal \N__62114\ : std_logic;
signal \N__62113\ : std_logic;
signal \N__62112\ : std_logic;
signal \N__62111\ : std_logic;
signal \N__62110\ : std_logic;
signal \N__62109\ : std_logic;
signal \N__62108\ : std_logic;
signal \N__62107\ : std_logic;
signal \N__62106\ : std_logic;
signal \N__62105\ : std_logic;
signal \N__62104\ : std_logic;
signal \N__62071\ : std_logic;
signal \N__62068\ : std_logic;
signal \N__62065\ : std_logic;
signal \N__62064\ : std_logic;
signal \N__62061\ : std_logic;
signal \N__62060\ : std_logic;
signal \N__62057\ : std_logic;
signal \N__62054\ : std_logic;
signal \N__62051\ : std_logic;
signal \N__62048\ : std_logic;
signal \N__62045\ : std_logic;
signal \N__62040\ : std_logic;
signal \N__62035\ : std_logic;
signal \N__62032\ : std_logic;
signal \N__62029\ : std_logic;
signal \N__62028\ : std_logic;
signal \N__62027\ : std_logic;
signal \N__62026\ : std_logic;
signal \N__62025\ : std_logic;
signal \N__62024\ : std_logic;
signal \N__62023\ : std_logic;
signal \N__62022\ : std_logic;
signal \N__62021\ : std_logic;
signal \N__62020\ : std_logic;
signal \N__62019\ : std_logic;
signal \N__62018\ : std_logic;
signal \N__62017\ : std_logic;
signal \N__62016\ : std_logic;
signal \N__62015\ : std_logic;
signal \N__61998\ : std_logic;
signal \N__61987\ : std_logic;
signal \N__61986\ : std_logic;
signal \N__61985\ : std_logic;
signal \N__61982\ : std_logic;
signal \N__61981\ : std_logic;
signal \N__61978\ : std_logic;
signal \N__61977\ : std_logic;
signal \N__61976\ : std_logic;
signal \N__61975\ : std_logic;
signal \N__61974\ : std_logic;
signal \N__61973\ : std_logic;
signal \N__61972\ : std_logic;
signal \N__61971\ : std_logic;
signal \N__61970\ : std_logic;
signal \N__61969\ : std_logic;
signal \N__61968\ : std_logic;
signal \N__61967\ : std_logic;
signal \N__61966\ : std_logic;
signal \N__61961\ : std_logic;
signal \N__61956\ : std_logic;
signal \N__61943\ : std_logic;
signal \N__61934\ : std_logic;
signal \N__61923\ : std_logic;
signal \N__61912\ : std_logic;
signal \N__61911\ : std_logic;
signal \N__61910\ : std_logic;
signal \N__61909\ : std_logic;
signal \N__61908\ : std_logic;
signal \N__61907\ : std_logic;
signal \N__61906\ : std_logic;
signal \N__61905\ : std_logic;
signal \N__61904\ : std_logic;
signal \N__61903\ : std_logic;
signal \N__61902\ : std_logic;
signal \N__61901\ : std_logic;
signal \N__61900\ : std_logic;
signal \N__61899\ : std_logic;
signal \N__61898\ : std_logic;
signal \N__61897\ : std_logic;
signal \N__61896\ : std_logic;
signal \N__61895\ : std_logic;
signal \N__61894\ : std_logic;
signal \N__61893\ : std_logic;
signal \N__61892\ : std_logic;
signal \N__61891\ : std_logic;
signal \N__61890\ : std_logic;
signal \N__61889\ : std_logic;
signal \N__61888\ : std_logic;
signal \N__61887\ : std_logic;
signal \N__61886\ : std_logic;
signal \N__61885\ : std_logic;
signal \N__61884\ : std_logic;
signal \N__61883\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61869\ : std_logic;
signal \N__61856\ : std_logic;
signal \N__61839\ : std_logic;
signal \N__61834\ : std_logic;
signal \N__61827\ : std_logic;
signal \N__61822\ : std_logic;
signal \N__61815\ : std_logic;
signal \N__61798\ : std_logic;
signal \N__61795\ : std_logic;
signal \N__61792\ : std_logic;
signal \N__61789\ : std_logic;
signal \N__61786\ : std_logic;
signal \N__61783\ : std_logic;
signal \N__61780\ : std_logic;
signal \N__61777\ : std_logic;
signal \N__61776\ : std_logic;
signal \N__61775\ : std_logic;
signal \N__61772\ : std_logic;
signal \N__61767\ : std_logic;
signal \N__61762\ : std_logic;
signal \N__61759\ : std_logic;
signal \N__61758\ : std_logic;
signal \N__61755\ : std_logic;
signal \N__61754\ : std_logic;
signal \N__61751\ : std_logic;
signal \N__61748\ : std_logic;
signal \N__61743\ : std_logic;
signal \N__61738\ : std_logic;
signal \N__61735\ : std_logic;
signal \N__61732\ : std_logic;
signal \N__61731\ : std_logic;
signal \N__61730\ : std_logic;
signal \N__61727\ : std_logic;
signal \N__61722\ : std_logic;
signal \N__61717\ : std_logic;
signal \N__61716\ : std_logic;
signal \N__61713\ : std_logic;
signal \N__61712\ : std_logic;
signal \N__61709\ : std_logic;
signal \N__61706\ : std_logic;
signal \N__61703\ : std_logic;
signal \N__61700\ : std_logic;
signal \N__61697\ : std_logic;
signal \N__61692\ : std_logic;
signal \N__61687\ : std_logic;
signal \N__61686\ : std_logic;
signal \N__61685\ : std_logic;
signal \N__61680\ : std_logic;
signal \N__61677\ : std_logic;
signal \N__61674\ : std_logic;
signal \N__61671\ : std_logic;
signal \N__61668\ : std_logic;
signal \N__61665\ : std_logic;
signal \N__61660\ : std_logic;
signal \N__61657\ : std_logic;
signal \N__61656\ : std_logic;
signal \N__61655\ : std_logic;
signal \N__61650\ : std_logic;
signal \N__61647\ : std_logic;
signal \N__61642\ : std_logic;
signal \N__61639\ : std_logic;
signal \N__61636\ : std_logic;
signal \N__61633\ : std_logic;
signal \N__61630\ : std_logic;
signal \N__61629\ : std_logic;
signal \N__61626\ : std_logic;
signal \N__61623\ : std_logic;
signal \N__61622\ : std_logic;
signal \N__61619\ : std_logic;
signal \N__61616\ : std_logic;
signal \N__61613\ : std_logic;
signal \N__61610\ : std_logic;
signal \N__61605\ : std_logic;
signal \N__61600\ : std_logic;
signal \N__61597\ : std_logic;
signal \N__61596\ : std_logic;
signal \N__61593\ : std_logic;
signal \N__61592\ : std_logic;
signal \N__61589\ : std_logic;
signal \N__61586\ : std_logic;
signal \N__61583\ : std_logic;
signal \N__61580\ : std_logic;
signal \N__61575\ : std_logic;
signal \N__61570\ : std_logic;
signal \N__61567\ : std_logic;
signal \N__61564\ : std_logic;
signal \N__61561\ : std_logic;
signal \N__61558\ : std_logic;
signal \N__61555\ : std_logic;
signal \N__61552\ : std_logic;
signal \N__61551\ : std_logic;
signal \N__61550\ : std_logic;
signal \N__61547\ : std_logic;
signal \N__61542\ : std_logic;
signal \N__61539\ : std_logic;
signal \N__61536\ : std_logic;
signal \N__61531\ : std_logic;
signal \N__61530\ : std_logic;
signal \N__61529\ : std_logic;
signal \N__61526\ : std_logic;
signal \N__61521\ : std_logic;
signal \N__61516\ : std_logic;
signal \N__61513\ : std_logic;
signal \N__61510\ : std_logic;
signal \N__61507\ : std_logic;
signal \N__61504\ : std_logic;
signal \N__61501\ : std_logic;
signal \N__61498\ : std_logic;
signal \N__61495\ : std_logic;
signal \N__61492\ : std_logic;
signal \N__61489\ : std_logic;
signal \N__61486\ : std_logic;
signal \N__61483\ : std_logic;
signal \N__61480\ : std_logic;
signal \N__61479\ : std_logic;
signal \N__61478\ : std_logic;
signal \N__61477\ : std_logic;
signal \N__61476\ : std_logic;
signal \N__61475\ : std_logic;
signal \N__61472\ : std_logic;
signal \N__61471\ : std_logic;
signal \N__61470\ : std_logic;
signal \N__61469\ : std_logic;
signal \N__61466\ : std_logic;
signal \N__61463\ : std_logic;
signal \N__61462\ : std_logic;
signal \N__61461\ : std_logic;
signal \N__61460\ : std_logic;
signal \N__61459\ : std_logic;
signal \N__61458\ : std_logic;
signal \N__61455\ : std_logic;
signal \N__61454\ : std_logic;
signal \N__61451\ : std_logic;
signal \N__61450\ : std_logic;
signal \N__61449\ : std_logic;
signal \N__61446\ : std_logic;
signal \N__61437\ : std_logic;
signal \N__61426\ : std_logic;
signal \N__61421\ : std_logic;
signal \N__61418\ : std_logic;
signal \N__61415\ : std_logic;
signal \N__61412\ : std_logic;
signal \N__61405\ : std_logic;
signal \N__61390\ : std_logic;
signal \N__61389\ : std_logic;
signal \N__61388\ : std_logic;
signal \N__61387\ : std_logic;
signal \N__61386\ : std_logic;
signal \N__61383\ : std_logic;
signal \N__61382\ : std_logic;
signal \N__61381\ : std_logic;
signal \N__61380\ : std_logic;
signal \N__61379\ : std_logic;
signal \N__61378\ : std_logic;
signal \N__61377\ : std_logic;
signal \N__61376\ : std_logic;
signal \N__61375\ : std_logic;
signal \N__61374\ : std_logic;
signal \N__61373\ : std_logic;
signal \N__61372\ : std_logic;
signal \N__61371\ : std_logic;
signal \N__61368\ : std_logic;
signal \N__61365\ : std_logic;
signal \N__61356\ : std_logic;
signal \N__61347\ : std_logic;
signal \N__61336\ : std_logic;
signal \N__61331\ : std_logic;
signal \N__61318\ : std_logic;
signal \N__61315\ : std_logic;
signal \N__61312\ : std_logic;
signal \N__61309\ : std_logic;
signal \N__61306\ : std_logic;
signal \N__61303\ : std_logic;
signal \N__61300\ : std_logic;
signal \N__61297\ : std_logic;
signal \N__61294\ : std_logic;
signal \N__61291\ : std_logic;
signal \N__61288\ : std_logic;
signal \N__61285\ : std_logic;
signal \N__61282\ : std_logic;
signal \N__61279\ : std_logic;
signal \N__61276\ : std_logic;
signal \N__61273\ : std_logic;
signal \N__61270\ : std_logic;
signal \N__61267\ : std_logic;
signal \N__61264\ : std_logic;
signal \N__61261\ : std_logic;
signal \N__61258\ : std_logic;
signal \N__61255\ : std_logic;
signal \N__61252\ : std_logic;
signal \N__61249\ : std_logic;
signal \N__61246\ : std_logic;
signal \N__61243\ : std_logic;
signal \N__61240\ : std_logic;
signal \N__61237\ : std_logic;
signal \N__61236\ : std_logic;
signal \N__61233\ : std_logic;
signal \N__61230\ : std_logic;
signal \N__61227\ : std_logic;
signal \N__61224\ : std_logic;
signal \N__61221\ : std_logic;
signal \N__61218\ : std_logic;
signal \N__61213\ : std_logic;
signal \N__61210\ : std_logic;
signal \N__61207\ : std_logic;
signal \N__61204\ : std_logic;
signal \N__61201\ : std_logic;
signal \N__61200\ : std_logic;
signal \N__61197\ : std_logic;
signal \N__61194\ : std_logic;
signal \N__61189\ : std_logic;
signal \N__61186\ : std_logic;
signal \N__61183\ : std_logic;
signal \N__61180\ : std_logic;
signal \N__61177\ : std_logic;
signal \N__61174\ : std_logic;
signal \N__61171\ : std_logic;
signal \N__61168\ : std_logic;
signal \N__61165\ : std_logic;
signal \N__61162\ : std_logic;
signal \N__61159\ : std_logic;
signal \N__61156\ : std_logic;
signal \N__61153\ : std_logic;
signal \N__61150\ : std_logic;
signal \N__61147\ : std_logic;
signal \N__61144\ : std_logic;
signal \N__61141\ : std_logic;
signal \N__61138\ : std_logic;
signal \N__61135\ : std_logic;
signal \N__61132\ : std_logic;
signal \N__61129\ : std_logic;
signal \N__61126\ : std_logic;
signal \N__61123\ : std_logic;
signal \N__61120\ : std_logic;
signal \N__61117\ : std_logic;
signal \N__61114\ : std_logic;
signal \N__61111\ : std_logic;
signal \N__61108\ : std_logic;
signal \N__61105\ : std_logic;
signal \N__61102\ : std_logic;
signal \N__61099\ : std_logic;
signal \N__61096\ : std_logic;
signal \N__61093\ : std_logic;
signal \N__61090\ : std_logic;
signal \N__61087\ : std_logic;
signal \N__61084\ : std_logic;
signal \N__61081\ : std_logic;
signal \N__61078\ : std_logic;
signal \N__61075\ : std_logic;
signal \N__61072\ : std_logic;
signal \N__61069\ : std_logic;
signal \N__61066\ : std_logic;
signal \N__61063\ : std_logic;
signal \N__61060\ : std_logic;
signal \N__61057\ : std_logic;
signal \N__61054\ : std_logic;
signal \N__61051\ : std_logic;
signal \N__61048\ : std_logic;
signal \N__61045\ : std_logic;
signal \N__61042\ : std_logic;
signal \N__61039\ : std_logic;
signal \N__61036\ : std_logic;
signal \N__61033\ : std_logic;
signal \N__61030\ : std_logic;
signal \N__61027\ : std_logic;
signal \N__61024\ : std_logic;
signal \N__61021\ : std_logic;
signal \N__61018\ : std_logic;
signal \N__61015\ : std_logic;
signal \N__61012\ : std_logic;
signal \N__61009\ : std_logic;
signal \N__61006\ : std_logic;
signal \N__61003\ : std_logic;
signal \N__61000\ : std_logic;
signal \N__60997\ : std_logic;
signal \N__60994\ : std_logic;
signal \N__60991\ : std_logic;
signal \N__60988\ : std_logic;
signal \N__60985\ : std_logic;
signal \N__60982\ : std_logic;
signal \N__60979\ : std_logic;
signal \N__60976\ : std_logic;
signal \N__60973\ : std_logic;
signal \N__60970\ : std_logic;
signal \N__60967\ : std_logic;
signal \N__60966\ : std_logic;
signal \N__60963\ : std_logic;
signal \N__60960\ : std_logic;
signal \N__60959\ : std_logic;
signal \N__60958\ : std_logic;
signal \N__60957\ : std_logic;
signal \N__60956\ : std_logic;
signal \N__60955\ : std_logic;
signal \N__60954\ : std_logic;
signal \N__60953\ : std_logic;
signal \N__60952\ : std_logic;
signal \N__60951\ : std_logic;
signal \N__60946\ : std_logic;
signal \N__60943\ : std_logic;
signal \N__60940\ : std_logic;
signal \N__60939\ : std_logic;
signal \N__60938\ : std_logic;
signal \N__60935\ : std_logic;
signal \N__60934\ : std_logic;
signal \N__60931\ : std_logic;
signal \N__60930\ : std_logic;
signal \N__60927\ : std_logic;
signal \N__60926\ : std_logic;
signal \N__60923\ : std_logic;
signal \N__60922\ : std_logic;
signal \N__60919\ : std_logic;
signal \N__60918\ : std_logic;
signal \N__60915\ : std_logic;
signal \N__60914\ : std_logic;
signal \N__60911\ : std_logic;
signal \N__60904\ : std_logic;
signal \N__60903\ : std_logic;
signal \N__60902\ : std_logic;
signal \N__60899\ : std_logic;
signal \N__60886\ : std_logic;
signal \N__60869\ : std_logic;
signal \N__60866\ : std_logic;
signal \N__60863\ : std_logic;
signal \N__60862\ : std_logic;
signal \N__60859\ : std_logic;
signal \N__60858\ : std_logic;
signal \N__60857\ : std_logic;
signal \N__60856\ : std_logic;
signal \N__60853\ : std_logic;
signal \N__60848\ : std_logic;
signal \N__60843\ : std_logic;
signal \N__60840\ : std_logic;
signal \N__60839\ : std_logic;
signal \N__60836\ : std_logic;
signal \N__60833\ : std_logic;
signal \N__60830\ : std_logic;
signal \N__60829\ : std_logic;
signal \N__60828\ : std_logic;
signal \N__60825\ : std_logic;
signal \N__60822\ : std_logic;
signal \N__60817\ : std_logic;
signal \N__60814\ : std_logic;
signal \N__60811\ : std_logic;
signal \N__60806\ : std_logic;
signal \N__60803\ : std_logic;
signal \N__60800\ : std_logic;
signal \N__60797\ : std_logic;
signal \N__60796\ : std_logic;
signal \N__60793\ : std_logic;
signal \N__60786\ : std_logic;
signal \N__60783\ : std_logic;
signal \N__60774\ : std_logic;
signal \N__60771\ : std_logic;
signal \N__60768\ : std_logic;
signal \N__60765\ : std_logic;
signal \N__60762\ : std_logic;
signal \N__60757\ : std_logic;
signal \N__60748\ : std_logic;
signal \N__60745\ : std_logic;
signal \N__60742\ : std_logic;
signal \N__60739\ : std_logic;
signal \N__60736\ : std_logic;
signal \N__60733\ : std_logic;
signal \N__60730\ : std_logic;
signal \N__60727\ : std_logic;
signal \N__60724\ : std_logic;
signal \N__60721\ : std_logic;
signal \N__60718\ : std_logic;
signal \N__60715\ : std_logic;
signal \N__60712\ : std_logic;
signal \N__60709\ : std_logic;
signal \N__60706\ : std_logic;
signal \N__60703\ : std_logic;
signal \N__60700\ : std_logic;
signal \N__60697\ : std_logic;
signal \N__60694\ : std_logic;
signal \N__60691\ : std_logic;
signal \N__60688\ : std_logic;
signal \N__60685\ : std_logic;
signal \N__60682\ : std_logic;
signal \N__60679\ : std_logic;
signal \N__60676\ : std_logic;
signal \N__60673\ : std_logic;
signal \N__60670\ : std_logic;
signal \N__60667\ : std_logic;
signal \N__60664\ : std_logic;
signal \N__60661\ : std_logic;
signal \N__60658\ : std_logic;
signal \N__60655\ : std_logic;
signal \N__60652\ : std_logic;
signal \N__60649\ : std_logic;
signal \N__60646\ : std_logic;
signal \N__60643\ : std_logic;
signal \N__60640\ : std_logic;
signal \N__60637\ : std_logic;
signal \N__60634\ : std_logic;
signal \N__60631\ : std_logic;
signal \N__60628\ : std_logic;
signal \N__60625\ : std_logic;
signal \N__60622\ : std_logic;
signal \N__60619\ : std_logic;
signal \N__60616\ : std_logic;
signal \N__60613\ : std_logic;
signal \N__60610\ : std_logic;
signal \N__60607\ : std_logic;
signal \N__60604\ : std_logic;
signal \N__60601\ : std_logic;
signal \N__60598\ : std_logic;
signal \N__60595\ : std_logic;
signal \N__60592\ : std_logic;
signal \N__60589\ : std_logic;
signal \N__60586\ : std_logic;
signal \N__60583\ : std_logic;
signal \N__60580\ : std_logic;
signal \N__60577\ : std_logic;
signal \N__60574\ : std_logic;
signal \N__60571\ : std_logic;
signal \N__60568\ : std_logic;
signal \N__60565\ : std_logic;
signal \N__60562\ : std_logic;
signal \N__60559\ : std_logic;
signal \N__60556\ : std_logic;
signal \N__60553\ : std_logic;
signal \N__60550\ : std_logic;
signal \N__60547\ : std_logic;
signal \N__60544\ : std_logic;
signal \N__60541\ : std_logic;
signal \N__60538\ : std_logic;
signal \N__60535\ : std_logic;
signal \N__60532\ : std_logic;
signal \N__60529\ : std_logic;
signal \N__60526\ : std_logic;
signal \N__60523\ : std_logic;
signal \N__60520\ : std_logic;
signal \N__60517\ : std_logic;
signal \N__60514\ : std_logic;
signal \N__60511\ : std_logic;
signal \N__60508\ : std_logic;
signal \N__60505\ : std_logic;
signal \N__60502\ : std_logic;
signal \N__60499\ : std_logic;
signal \N__60496\ : std_logic;
signal \N__60493\ : std_logic;
signal \N__60490\ : std_logic;
signal \N__60487\ : std_logic;
signal \N__60484\ : std_logic;
signal \N__60481\ : std_logic;
signal \N__60478\ : std_logic;
signal \N__60475\ : std_logic;
signal \N__60472\ : std_logic;
signal \N__60469\ : std_logic;
signal \N__60466\ : std_logic;
signal \N__60463\ : std_logic;
signal \N__60460\ : std_logic;
signal \N__60457\ : std_logic;
signal \N__60454\ : std_logic;
signal \N__60451\ : std_logic;
signal \N__60448\ : std_logic;
signal \N__60447\ : std_logic;
signal \N__60444\ : std_logic;
signal \N__60443\ : std_logic;
signal \N__60442\ : std_logic;
signal \N__60441\ : std_logic;
signal \N__60438\ : std_logic;
signal \N__60433\ : std_logic;
signal \N__60426\ : std_logic;
signal \N__60421\ : std_logic;
signal \N__60418\ : std_logic;
signal \N__60415\ : std_logic;
signal \N__60412\ : std_logic;
signal \N__60411\ : std_logic;
signal \N__60408\ : std_logic;
signal \N__60405\ : std_logic;
signal \N__60402\ : std_logic;
signal \N__60399\ : std_logic;
signal \N__60398\ : std_logic;
signal \N__60395\ : std_logic;
signal \N__60392\ : std_logic;
signal \N__60389\ : std_logic;
signal \N__60382\ : std_logic;
signal \N__60381\ : std_logic;
signal \N__60376\ : std_logic;
signal \N__60375\ : std_logic;
signal \N__60372\ : std_logic;
signal \N__60369\ : std_logic;
signal \N__60366\ : std_logic;
signal \N__60363\ : std_logic;
signal \N__60358\ : std_logic;
signal \N__60355\ : std_logic;
signal \N__60354\ : std_logic;
signal \N__60351\ : std_logic;
signal \N__60348\ : std_logic;
signal \N__60345\ : std_logic;
signal \N__60342\ : std_logic;
signal \N__60341\ : std_logic;
signal \N__60336\ : std_logic;
signal \N__60333\ : std_logic;
signal \N__60328\ : std_logic;
signal \N__60327\ : std_logic;
signal \N__60322\ : std_logic;
signal \N__60321\ : std_logic;
signal \N__60318\ : std_logic;
signal \N__60315\ : std_logic;
signal \N__60310\ : std_logic;
signal \N__60309\ : std_logic;
signal \N__60304\ : std_logic;
signal \N__60303\ : std_logic;
signal \N__60300\ : std_logic;
signal \N__60297\ : std_logic;
signal \N__60292\ : std_logic;
signal \N__60289\ : std_logic;
signal \N__60286\ : std_logic;
signal \N__60285\ : std_logic;
signal \N__60282\ : std_logic;
signal \N__60279\ : std_logic;
signal \N__60274\ : std_logic;
signal \N__60271\ : std_logic;
signal \N__60270\ : std_logic;
signal \N__60267\ : std_logic;
signal \N__60264\ : std_logic;
signal \N__60259\ : std_logic;
signal \N__60258\ : std_logic;
signal \N__60255\ : std_logic;
signal \N__60252\ : std_logic;
signal \N__60251\ : std_logic;
signal \N__60248\ : std_logic;
signal \N__60245\ : std_logic;
signal \N__60242\ : std_logic;
signal \N__60239\ : std_logic;
signal \N__60234\ : std_logic;
signal \N__60229\ : std_logic;
signal \N__60226\ : std_logic;
signal \N__60223\ : std_logic;
signal \N__60222\ : std_logic;
signal \N__60219\ : std_logic;
signal \N__60216\ : std_logic;
signal \N__60215\ : std_logic;
signal \N__60212\ : std_logic;
signal \N__60209\ : std_logic;
signal \N__60206\ : std_logic;
signal \N__60199\ : std_logic;
signal \N__60196\ : std_logic;
signal \N__60193\ : std_logic;
signal \N__60190\ : std_logic;
signal \N__60189\ : std_logic;
signal \N__60186\ : std_logic;
signal \N__60183\ : std_logic;
signal \N__60178\ : std_logic;
signal \N__60175\ : std_logic;
signal \N__60174\ : std_logic;
signal \N__60171\ : std_logic;
signal \N__60168\ : std_logic;
signal \N__60163\ : std_logic;
signal \N__60160\ : std_logic;
signal \N__60157\ : std_logic;
signal \N__60154\ : std_logic;
signal \N__60151\ : std_logic;
signal \N__60148\ : std_logic;
signal \N__60147\ : std_logic;
signal \N__60144\ : std_logic;
signal \N__60141\ : std_logic;
signal \N__60140\ : std_logic;
signal \N__60137\ : std_logic;
signal \N__60132\ : std_logic;
signal \N__60127\ : std_logic;
signal \N__60124\ : std_logic;
signal \N__60123\ : std_logic;
signal \N__60120\ : std_logic;
signal \N__60117\ : std_logic;
signal \N__60112\ : std_logic;
signal \N__60111\ : std_logic;
signal \N__60110\ : std_logic;
signal \N__60107\ : std_logic;
signal \N__60102\ : std_logic;
signal \N__60097\ : std_logic;
signal \N__60094\ : std_logic;
signal \N__60093\ : std_logic;
signal \N__60092\ : std_logic;
signal \N__60089\ : std_logic;
signal \N__60084\ : std_logic;
signal \N__60079\ : std_logic;
signal \N__60076\ : std_logic;
signal \N__60073\ : std_logic;
signal \N__60070\ : std_logic;
signal \N__60069\ : std_logic;
signal \N__60068\ : std_logic;
signal \N__60065\ : std_logic;
signal \N__60060\ : std_logic;
signal \N__60055\ : std_logic;
signal \N__60052\ : std_logic;
signal \N__60049\ : std_logic;
signal \N__60046\ : std_logic;
signal \N__60043\ : std_logic;
signal \N__60040\ : std_logic;
signal \N__60037\ : std_logic;
signal \N__60034\ : std_logic;
signal \N__60031\ : std_logic;
signal \N__60028\ : std_logic;
signal \N__60025\ : std_logic;
signal \N__60022\ : std_logic;
signal \N__60019\ : std_logic;
signal \N__60016\ : std_logic;
signal \N__60013\ : std_logic;
signal \N__60010\ : std_logic;
signal \N__60007\ : std_logic;
signal \N__60006\ : std_logic;
signal \N__60005\ : std_logic;
signal \N__59998\ : std_logic;
signal \N__59995\ : std_logic;
signal \N__59992\ : std_logic;
signal \N__59989\ : std_logic;
signal \N__59986\ : std_logic;
signal \N__59983\ : std_logic;
signal \N__59980\ : std_logic;
signal \N__59977\ : std_logic;
signal \N__59974\ : std_logic;
signal \N__59973\ : std_logic;
signal \N__59972\ : std_logic;
signal \N__59965\ : std_logic;
signal \N__59962\ : std_logic;
signal \N__59959\ : std_logic;
signal \N__59956\ : std_logic;
signal \N__59953\ : std_logic;
signal \N__59950\ : std_logic;
signal \N__59947\ : std_logic;
signal \N__59944\ : std_logic;
signal \N__59941\ : std_logic;
signal \N__59938\ : std_logic;
signal \N__59935\ : std_logic;
signal \N__59932\ : std_logic;
signal \N__59929\ : std_logic;
signal \N__59926\ : std_logic;
signal \N__59923\ : std_logic;
signal \N__59920\ : std_logic;
signal \N__59917\ : std_logic;
signal \N__59914\ : std_logic;
signal \N__59911\ : std_logic;
signal \N__59908\ : std_logic;
signal \N__59905\ : std_logic;
signal \N__59902\ : std_logic;
signal \N__59899\ : std_logic;
signal \N__59896\ : std_logic;
signal \N__59893\ : std_logic;
signal \N__59890\ : std_logic;
signal \N__59887\ : std_logic;
signal \N__59884\ : std_logic;
signal \N__59881\ : std_logic;
signal \N__59878\ : std_logic;
signal \N__59875\ : std_logic;
signal \N__59872\ : std_logic;
signal \N__59869\ : std_logic;
signal \N__59866\ : std_logic;
signal \N__59863\ : std_logic;
signal \N__59860\ : std_logic;
signal \N__59857\ : std_logic;
signal \N__59854\ : std_logic;
signal \N__59851\ : std_logic;
signal \N__59848\ : std_logic;
signal \N__59845\ : std_logic;
signal \N__59842\ : std_logic;
signal \N__59839\ : std_logic;
signal \N__59836\ : std_logic;
signal \N__59833\ : std_logic;
signal \N__59830\ : std_logic;
signal \N__59827\ : std_logic;
signal \N__59824\ : std_logic;
signal \N__59821\ : std_logic;
signal \N__59818\ : std_logic;
signal \N__59815\ : std_logic;
signal \N__59812\ : std_logic;
signal \N__59809\ : std_logic;
signal \N__59806\ : std_logic;
signal \N__59803\ : std_logic;
signal \N__59800\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59794\ : std_logic;
signal \N__59791\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59787\ : std_logic;
signal \N__59786\ : std_logic;
signal \N__59783\ : std_logic;
signal \N__59778\ : std_logic;
signal \N__59773\ : std_logic;
signal \N__59770\ : std_logic;
signal \N__59767\ : std_logic;
signal \N__59764\ : std_logic;
signal \N__59761\ : std_logic;
signal \N__59758\ : std_logic;
signal \N__59755\ : std_logic;
signal \N__59752\ : std_logic;
signal \N__59749\ : std_logic;
signal \N__59746\ : std_logic;
signal \N__59743\ : std_logic;
signal \N__59740\ : std_logic;
signal \N__59737\ : std_logic;
signal \N__59734\ : std_logic;
signal \N__59731\ : std_logic;
signal \N__59728\ : std_logic;
signal \N__59725\ : std_logic;
signal \N__59722\ : std_logic;
signal \N__59719\ : std_logic;
signal \N__59716\ : std_logic;
signal \N__59713\ : std_logic;
signal \N__59710\ : std_logic;
signal \N__59707\ : std_logic;
signal \N__59704\ : std_logic;
signal \N__59701\ : std_logic;
signal \N__59698\ : std_logic;
signal \N__59695\ : std_logic;
signal \N__59692\ : std_logic;
signal \N__59689\ : std_logic;
signal \N__59686\ : std_logic;
signal \N__59683\ : std_logic;
signal \N__59680\ : std_logic;
signal \N__59677\ : std_logic;
signal \N__59674\ : std_logic;
signal \N__59671\ : std_logic;
signal \N__59668\ : std_logic;
signal \N__59665\ : std_logic;
signal \N__59662\ : std_logic;
signal \N__59659\ : std_logic;
signal \N__59656\ : std_logic;
signal \N__59653\ : std_logic;
signal \N__59650\ : std_logic;
signal \N__59647\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59641\ : std_logic;
signal \N__59638\ : std_logic;
signal \N__59635\ : std_logic;
signal \N__59632\ : std_logic;
signal \N__59629\ : std_logic;
signal \N__59626\ : std_logic;
signal \N__59623\ : std_logic;
signal \N__59620\ : std_logic;
signal \N__59617\ : std_logic;
signal \N__59614\ : std_logic;
signal \N__59611\ : std_logic;
signal \N__59608\ : std_logic;
signal \N__59605\ : std_logic;
signal \N__59602\ : std_logic;
signal \N__59599\ : std_logic;
signal \N__59596\ : std_logic;
signal \N__59593\ : std_logic;
signal \N__59590\ : std_logic;
signal \N__59587\ : std_logic;
signal \N__59584\ : std_logic;
signal \N__59581\ : std_logic;
signal \N__59578\ : std_logic;
signal \N__59575\ : std_logic;
signal \N__59572\ : std_logic;
signal \N__59569\ : std_logic;
signal \N__59566\ : std_logic;
signal \N__59563\ : std_logic;
signal \N__59560\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59551\ : std_logic;
signal \N__59548\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59542\ : std_logic;
signal \N__59539\ : std_logic;
signal \N__59536\ : std_logic;
signal \N__59533\ : std_logic;
signal \N__59530\ : std_logic;
signal \N__59527\ : std_logic;
signal \N__59524\ : std_logic;
signal \N__59521\ : std_logic;
signal \N__59518\ : std_logic;
signal \N__59515\ : std_logic;
signal \N__59512\ : std_logic;
signal \N__59509\ : std_logic;
signal \N__59506\ : std_logic;
signal \N__59503\ : std_logic;
signal \N__59500\ : std_logic;
signal \N__59497\ : std_logic;
signal \N__59494\ : std_logic;
signal \N__59491\ : std_logic;
signal \N__59488\ : std_logic;
signal \N__59485\ : std_logic;
signal \N__59482\ : std_logic;
signal \N__59481\ : std_logic;
signal \N__59476\ : std_logic;
signal \N__59473\ : std_logic;
signal \N__59470\ : std_logic;
signal \N__59467\ : std_logic;
signal \N__59466\ : std_logic;
signal \N__59465\ : std_logic;
signal \N__59462\ : std_logic;
signal \N__59459\ : std_logic;
signal \N__59456\ : std_logic;
signal \N__59449\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59443\ : std_logic;
signal \N__59442\ : std_logic;
signal \N__59441\ : std_logic;
signal \N__59440\ : std_logic;
signal \N__59437\ : std_logic;
signal \N__59434\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59430\ : std_logic;
signal \N__59429\ : std_logic;
signal \N__59428\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59425\ : std_logic;
signal \N__59424\ : std_logic;
signal \N__59423\ : std_logic;
signal \N__59420\ : std_logic;
signal \N__59419\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59417\ : std_logic;
signal \N__59416\ : std_logic;
signal \N__59415\ : std_logic;
signal \N__59412\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59402\ : std_logic;
signal \N__59391\ : std_logic;
signal \N__59388\ : std_logic;
signal \N__59381\ : std_logic;
signal \N__59374\ : std_logic;
signal \N__59359\ : std_logic;
signal \N__59358\ : std_logic;
signal \N__59355\ : std_logic;
signal \N__59352\ : std_logic;
signal \N__59351\ : std_logic;
signal \N__59350\ : std_logic;
signal \N__59345\ : std_logic;
signal \N__59342\ : std_logic;
signal \N__59339\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59331\ : std_logic;
signal \N__59326\ : std_logic;
signal \N__59325\ : std_logic;
signal \N__59322\ : std_logic;
signal \N__59319\ : std_logic;
signal \N__59316\ : std_logic;
signal \N__59315\ : std_logic;
signal \N__59312\ : std_logic;
signal \N__59309\ : std_logic;
signal \N__59308\ : std_logic;
signal \N__59307\ : std_logic;
signal \N__59306\ : std_logic;
signal \N__59305\ : std_logic;
signal \N__59304\ : std_logic;
signal \N__59301\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59299\ : std_logic;
signal \N__59298\ : std_logic;
signal \N__59297\ : std_logic;
signal \N__59296\ : std_logic;
signal \N__59295\ : std_logic;
signal \N__59294\ : std_logic;
signal \N__59293\ : std_logic;
signal \N__59292\ : std_logic;
signal \N__59287\ : std_logic;
signal \N__59280\ : std_logic;
signal \N__59269\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59259\ : std_logic;
signal \N__59252\ : std_logic;
signal \N__59239\ : std_logic;
signal \N__59236\ : std_logic;
signal \N__59233\ : std_logic;
signal \N__59230\ : std_logic;
signal \N__59227\ : std_logic;
signal \N__59224\ : std_logic;
signal \N__59221\ : std_logic;
signal \N__59218\ : std_logic;
signal \N__59215\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59209\ : std_logic;
signal \N__59206\ : std_logic;
signal \N__59203\ : std_logic;
signal \N__59200\ : std_logic;
signal \N__59197\ : std_logic;
signal \N__59196\ : std_logic;
signal \N__59191\ : std_logic;
signal \N__59188\ : std_logic;
signal \N__59185\ : std_logic;
signal \N__59182\ : std_logic;
signal \N__59181\ : std_logic;
signal \N__59180\ : std_logic;
signal \N__59177\ : std_logic;
signal \N__59174\ : std_logic;
signal \N__59171\ : std_logic;
signal \N__59164\ : std_logic;
signal \N__59161\ : std_logic;
signal \N__59158\ : std_logic;
signal \N__59155\ : std_logic;
signal \N__59152\ : std_logic;
signal \N__59151\ : std_logic;
signal \N__59150\ : std_logic;
signal \N__59147\ : std_logic;
signal \N__59144\ : std_logic;
signal \N__59141\ : std_logic;
signal \N__59134\ : std_logic;
signal \N__59131\ : std_logic;
signal \N__59128\ : std_logic;
signal \N__59125\ : std_logic;
signal \N__59122\ : std_logic;
signal \N__59119\ : std_logic;
signal \N__59116\ : std_logic;
signal \N__59113\ : std_logic;
signal \N__59110\ : std_logic;
signal \N__59107\ : std_logic;
signal \N__59104\ : std_logic;
signal \N__59101\ : std_logic;
signal \N__59098\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59092\ : std_logic;
signal \N__59089\ : std_logic;
signal \N__59086\ : std_logic;
signal \N__59083\ : std_logic;
signal \N__59080\ : std_logic;
signal \N__59077\ : std_logic;
signal \N__59074\ : std_logic;
signal \N__59071\ : std_logic;
signal \N__59068\ : std_logic;
signal \N__59065\ : std_logic;
signal \N__59062\ : std_logic;
signal \N__59059\ : std_logic;
signal \N__59056\ : std_logic;
signal \N__59053\ : std_logic;
signal \N__59050\ : std_logic;
signal \N__59047\ : std_logic;
signal \N__59044\ : std_logic;
signal \N__59041\ : std_logic;
signal \N__59038\ : std_logic;
signal \N__59035\ : std_logic;
signal \N__59032\ : std_logic;
signal \N__59029\ : std_logic;
signal \N__59026\ : std_logic;
signal \N__59023\ : std_logic;
signal \N__59020\ : std_logic;
signal \N__59017\ : std_logic;
signal \N__59014\ : std_logic;
signal \N__59011\ : std_logic;
signal \N__59008\ : std_logic;
signal \N__59005\ : std_logic;
signal \N__59002\ : std_logic;
signal \N__58999\ : std_logic;
signal \N__58996\ : std_logic;
signal \N__58993\ : std_logic;
signal \N__58990\ : std_logic;
signal \N__58987\ : std_logic;
signal \N__58984\ : std_logic;
signal \N__58983\ : std_logic;
signal \N__58980\ : std_logic;
signal \N__58977\ : std_logic;
signal \N__58972\ : std_logic;
signal \N__58969\ : std_logic;
signal \N__58966\ : std_logic;
signal \N__58963\ : std_logic;
signal \N__58960\ : std_logic;
signal \N__58957\ : std_logic;
signal \N__58954\ : std_logic;
signal \N__58951\ : std_logic;
signal \N__58948\ : std_logic;
signal \N__58945\ : std_logic;
signal \N__58942\ : std_logic;
signal \N__58939\ : std_logic;
signal \N__58936\ : std_logic;
signal \N__58933\ : std_logic;
signal \N__58930\ : std_logic;
signal \N__58927\ : std_logic;
signal \N__58924\ : std_logic;
signal \N__58921\ : std_logic;
signal \N__58918\ : std_logic;
signal \N__58915\ : std_logic;
signal \N__58912\ : std_logic;
signal \N__58911\ : std_logic;
signal \N__58910\ : std_logic;
signal \N__58909\ : std_logic;
signal \N__58908\ : std_logic;
signal \N__58907\ : std_logic;
signal \N__58906\ : std_logic;
signal \N__58905\ : std_logic;
signal \N__58904\ : std_logic;
signal \N__58903\ : std_logic;
signal \N__58902\ : std_logic;
signal \N__58901\ : std_logic;
signal \N__58900\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58895\ : std_logic;
signal \N__58892\ : std_logic;
signal \N__58891\ : std_logic;
signal \N__58888\ : std_logic;
signal \N__58887\ : std_logic;
signal \N__58884\ : std_logic;
signal \N__58881\ : std_logic;
signal \N__58878\ : std_logic;
signal \N__58875\ : std_logic;
signal \N__58874\ : std_logic;
signal \N__58871\ : std_logic;
signal \N__58870\ : std_logic;
signal \N__58867\ : std_logic;
signal \N__58866\ : std_logic;
signal \N__58865\ : std_logic;
signal \N__58864\ : std_logic;
signal \N__58861\ : std_logic;
signal \N__58860\ : std_logic;
signal \N__58857\ : std_logic;
signal \N__58856\ : std_logic;
signal \N__58853\ : std_logic;
signal \N__58852\ : std_logic;
signal \N__58849\ : std_logic;
signal \N__58846\ : std_logic;
signal \N__58845\ : std_logic;
signal \N__58842\ : std_logic;
signal \N__58829\ : std_logic;
signal \N__58826\ : std_logic;
signal \N__58823\ : std_logic;
signal \N__58820\ : std_logic;
signal \N__58817\ : std_logic;
signal \N__58814\ : std_logic;
signal \N__58811\ : std_logic;
signal \N__58810\ : std_logic;
signal \N__58807\ : std_logic;
signal \N__58804\ : std_logic;
signal \N__58801\ : std_logic;
signal \N__58784\ : std_logic;
signal \N__58781\ : std_logic;
signal \N__58780\ : std_logic;
signal \N__58777\ : std_logic;
signal \N__58772\ : std_logic;
signal \N__58765\ : std_logic;
signal \N__58762\ : std_logic;
signal \N__58759\ : std_logic;
signal \N__58756\ : std_logic;
signal \N__58755\ : std_logic;
signal \N__58752\ : std_logic;
signal \N__58747\ : std_logic;
signal \N__58740\ : std_logic;
signal \N__58737\ : std_logic;
signal \N__58734\ : std_logic;
signal \N__58731\ : std_logic;
signal \N__58722\ : std_logic;
signal \N__58719\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58707\ : std_logic;
signal \N__58698\ : std_logic;
signal \N__58695\ : std_logic;
signal \N__58692\ : std_logic;
signal \N__58687\ : std_logic;
signal \N__58684\ : std_logic;
signal \N__58681\ : std_logic;
signal \N__58678\ : std_logic;
signal \N__58675\ : std_logic;
signal \N__58672\ : std_logic;
signal \N__58669\ : std_logic;
signal \N__58666\ : std_logic;
signal \N__58663\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58657\ : std_logic;
signal \N__58654\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58648\ : std_logic;
signal \N__58645\ : std_logic;
signal \N__58642\ : std_logic;
signal \N__58639\ : std_logic;
signal \N__58636\ : std_logic;
signal \N__58633\ : std_logic;
signal \N__58630\ : std_logic;
signal \N__58627\ : std_logic;
signal \N__58624\ : std_logic;
signal \N__58621\ : std_logic;
signal \N__58618\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58612\ : std_logic;
signal \N__58609\ : std_logic;
signal \N__58606\ : std_logic;
signal \N__58603\ : std_logic;
signal \N__58600\ : std_logic;
signal \N__58597\ : std_logic;
signal \N__58594\ : std_logic;
signal \N__58591\ : std_logic;
signal \N__58588\ : std_logic;
signal \N__58585\ : std_logic;
signal \N__58582\ : std_logic;
signal \N__58579\ : std_logic;
signal \N__58576\ : std_logic;
signal \N__58573\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58567\ : std_logic;
signal \N__58564\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58558\ : std_logic;
signal \N__58555\ : std_logic;
signal \N__58552\ : std_logic;
signal \N__58549\ : std_logic;
signal \N__58546\ : std_logic;
signal \N__58543\ : std_logic;
signal \N__58540\ : std_logic;
signal \N__58537\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58531\ : std_logic;
signal \N__58528\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58522\ : std_logic;
signal \N__58519\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58513\ : std_logic;
signal \N__58512\ : std_logic;
signal \N__58509\ : std_logic;
signal \N__58506\ : std_logic;
signal \N__58503\ : std_logic;
signal \N__58500\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58494\ : std_logic;
signal \N__58489\ : std_logic;
signal \N__58488\ : std_logic;
signal \N__58487\ : std_logic;
signal \N__58482\ : std_logic;
signal \N__58479\ : std_logic;
signal \N__58476\ : std_logic;
signal \N__58473\ : std_logic;
signal \N__58470\ : std_logic;
signal \N__58467\ : std_logic;
signal \N__58464\ : std_logic;
signal \N__58459\ : std_logic;
signal \N__58456\ : std_logic;
signal \N__58453\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58451\ : std_logic;
signal \N__58450\ : std_logic;
signal \N__58447\ : std_logic;
signal \N__58446\ : std_logic;
signal \N__58443\ : std_logic;
signal \N__58442\ : std_logic;
signal \N__58439\ : std_logic;
signal \N__58438\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58434\ : std_logic;
signal \N__58433\ : std_logic;
signal \N__58430\ : std_logic;
signal \N__58415\ : std_logic;
signal \N__58412\ : std_logic;
signal \N__58405\ : std_logic;
signal \N__58404\ : std_logic;
signal \N__58403\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58399\ : std_logic;
signal \N__58396\ : std_logic;
signal \N__58395\ : std_logic;
signal \N__58392\ : std_logic;
signal \N__58381\ : std_logic;
signal \N__58378\ : std_logic;
signal \N__58375\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58369\ : std_logic;
signal \N__58368\ : std_logic;
signal \N__58367\ : std_logic;
signal \N__58364\ : std_logic;
signal \N__58361\ : std_logic;
signal \N__58358\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58350\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58344\ : std_logic;
signal \N__58339\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58333\ : std_logic;
signal \N__58330\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58324\ : std_logic;
signal \N__58321\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58315\ : std_logic;
signal \N__58312\ : std_logic;
signal \N__58309\ : std_logic;
signal \N__58306\ : std_logic;
signal \N__58303\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58297\ : std_logic;
signal \N__58294\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58288\ : std_logic;
signal \N__58285\ : std_logic;
signal \N__58282\ : std_logic;
signal \N__58279\ : std_logic;
signal \N__58278\ : std_logic;
signal \N__58275\ : std_logic;
signal \N__58272\ : std_logic;
signal \N__58269\ : std_logic;
signal \N__58266\ : std_logic;
signal \N__58263\ : std_logic;
signal \N__58260\ : std_logic;
signal \N__58255\ : std_logic;
signal \N__58252\ : std_logic;
signal \N__58249\ : std_logic;
signal \N__58246\ : std_logic;
signal \N__58243\ : std_logic;
signal \N__58240\ : std_logic;
signal \N__58239\ : std_logic;
signal \N__58238\ : std_logic;
signal \N__58235\ : std_logic;
signal \N__58232\ : std_logic;
signal \N__58229\ : std_logic;
signal \N__58222\ : std_logic;
signal \N__58219\ : std_logic;
signal \N__58216\ : std_logic;
signal \N__58213\ : std_logic;
signal \N__58212\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58203\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58197\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58191\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58183\ : std_logic;
signal \N__58180\ : std_logic;
signal \N__58177\ : std_logic;
signal \N__58174\ : std_logic;
signal \N__58171\ : std_logic;
signal \N__58170\ : std_logic;
signal \N__58169\ : std_logic;
signal \N__58164\ : std_logic;
signal \N__58161\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58150\ : std_logic;
signal \N__58147\ : std_logic;
signal \N__58144\ : std_logic;
signal \N__58141\ : std_logic;
signal \N__58140\ : std_logic;
signal \N__58137\ : std_logic;
signal \N__58134\ : std_logic;
signal \N__58129\ : std_logic;
signal \N__58126\ : std_logic;
signal \N__58123\ : std_logic;
signal \N__58120\ : std_logic;
signal \N__58117\ : std_logic;
signal \N__58114\ : std_logic;
signal \N__58111\ : std_logic;
signal \N__58110\ : std_logic;
signal \N__58109\ : std_logic;
signal \N__58106\ : std_logic;
signal \N__58101\ : std_logic;
signal \N__58098\ : std_logic;
signal \N__58095\ : std_logic;
signal \N__58092\ : std_logic;
signal \N__58089\ : std_logic;
signal \N__58084\ : std_logic;
signal \N__58081\ : std_logic;
signal \N__58080\ : std_logic;
signal \N__58077\ : std_logic;
signal \N__58074\ : std_logic;
signal \N__58071\ : std_logic;
signal \N__58068\ : std_logic;
signal \N__58065\ : std_logic;
signal \N__58062\ : std_logic;
signal \N__58057\ : std_logic;
signal \N__58054\ : std_logic;
signal \N__58051\ : std_logic;
signal \N__58048\ : std_logic;
signal \N__58045\ : std_logic;
signal \N__58042\ : std_logic;
signal \N__58041\ : std_logic;
signal \N__58040\ : std_logic;
signal \N__58035\ : std_logic;
signal \N__58032\ : std_logic;
signal \N__58029\ : std_logic;
signal \N__58026\ : std_logic;
signal \N__58021\ : std_logic;
signal \N__58018\ : std_logic;
signal \N__58015\ : std_logic;
signal \N__58012\ : std_logic;
signal \N__58011\ : std_logic;
signal \N__58008\ : std_logic;
signal \N__58005\ : std_logic;
signal \N__58002\ : std_logic;
signal \N__57999\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57991\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57987\ : std_logic;
signal \N__57986\ : std_logic;
signal \N__57981\ : std_logic;
signal \N__57978\ : std_logic;
signal \N__57973\ : std_logic;
signal \N__57970\ : std_logic;
signal \N__57967\ : std_logic;
signal \N__57964\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57954\ : std_logic;
signal \N__57951\ : std_logic;
signal \N__57948\ : std_logic;
signal \N__57945\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57939\ : std_logic;
signal \N__57938\ : std_logic;
signal \N__57935\ : std_logic;
signal \N__57932\ : std_logic;
signal \N__57929\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57919\ : std_logic;
signal \N__57916\ : std_logic;
signal \N__57913\ : std_logic;
signal \N__57910\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57906\ : std_logic;
signal \N__57903\ : std_logic;
signal \N__57898\ : std_logic;
signal \N__57895\ : std_logic;
signal \N__57892\ : std_logic;
signal \N__57889\ : std_logic;
signal \N__57888\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57884\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57871\ : std_logic;
signal \N__57868\ : std_logic;
signal \N__57865\ : std_logic;
signal \N__57862\ : std_logic;
signal \N__57859\ : std_logic;
signal \N__57856\ : std_logic;
signal \N__57853\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57838\ : std_logic;
signal \N__57835\ : std_logic;
signal \N__57832\ : std_logic;
signal \N__57829\ : std_logic;
signal \N__57826\ : std_logic;
signal \N__57823\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57817\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57810\ : std_logic;
signal \N__57807\ : std_logic;
signal \N__57802\ : std_logic;
signal \N__57799\ : std_logic;
signal \N__57796\ : std_logic;
signal \N__57793\ : std_logic;
signal \N__57790\ : std_logic;
signal \N__57787\ : std_logic;
signal \N__57786\ : std_logic;
signal \N__57785\ : std_logic;
signal \N__57782\ : std_logic;
signal \N__57779\ : std_logic;
signal \N__57776\ : std_logic;
signal \N__57773\ : std_logic;
signal \N__57770\ : std_logic;
signal \N__57767\ : std_logic;
signal \N__57762\ : std_logic;
signal \N__57759\ : std_logic;
signal \N__57754\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57748\ : std_logic;
signal \N__57745\ : std_logic;
signal \N__57744\ : std_logic;
signal \N__57741\ : std_logic;
signal \N__57738\ : std_logic;
signal \N__57733\ : std_logic;
signal \N__57730\ : std_logic;
signal \N__57727\ : std_logic;
signal \N__57724\ : std_logic;
signal \N__57721\ : std_logic;
signal \N__57718\ : std_logic;
signal \N__57717\ : std_logic;
signal \N__57716\ : std_logic;
signal \N__57713\ : std_logic;
signal \N__57710\ : std_logic;
signal \N__57707\ : std_logic;
signal \N__57704\ : std_logic;
signal \N__57699\ : std_logic;
signal \N__57696\ : std_logic;
signal \N__57693\ : std_logic;
signal \N__57688\ : std_logic;
signal \N__57685\ : std_logic;
signal \N__57684\ : std_logic;
signal \N__57681\ : std_logic;
signal \N__57678\ : std_logic;
signal \N__57675\ : std_logic;
signal \N__57672\ : std_logic;
signal \N__57669\ : std_logic;
signal \N__57666\ : std_logic;
signal \N__57661\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57649\ : std_logic;
signal \N__57646\ : std_logic;
signal \N__57643\ : std_logic;
signal \N__57640\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57636\ : std_logic;
signal \N__57635\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57629\ : std_logic;
signal \N__57626\ : std_logic;
signal \N__57623\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57612\ : std_logic;
signal \N__57609\ : std_logic;
signal \N__57604\ : std_logic;
signal \N__57601\ : std_logic;
signal \N__57600\ : std_logic;
signal \N__57597\ : std_logic;
signal \N__57594\ : std_logic;
signal \N__57591\ : std_logic;
signal \N__57588\ : std_logic;
signal \N__57585\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57577\ : std_logic;
signal \N__57574\ : std_logic;
signal \N__57571\ : std_logic;
signal \N__57568\ : std_logic;
signal \N__57565\ : std_logic;
signal \N__57562\ : std_logic;
signal \N__57561\ : std_logic;
signal \N__57558\ : std_logic;
signal \N__57555\ : std_logic;
signal \N__57552\ : std_logic;
signal \N__57551\ : std_logic;
signal \N__57548\ : std_logic;
signal \N__57545\ : std_logic;
signal \N__57542\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57529\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57525\ : std_logic;
signal \N__57522\ : std_logic;
signal \N__57519\ : std_logic;
signal \N__57514\ : std_logic;
signal \N__57511\ : std_logic;
signal \N__57508\ : std_logic;
signal \N__57505\ : std_logic;
signal \N__57502\ : std_logic;
signal \N__57499\ : std_logic;
signal \N__57496\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57492\ : std_logic;
signal \N__57491\ : std_logic;
signal \N__57488\ : std_logic;
signal \N__57485\ : std_logic;
signal \N__57482\ : std_logic;
signal \N__57479\ : std_logic;
signal \N__57474\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57466\ : std_logic;
signal \N__57463\ : std_logic;
signal \N__57460\ : std_logic;
signal \N__57457\ : std_logic;
signal \N__57456\ : std_logic;
signal \N__57453\ : std_logic;
signal \N__57450\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57439\ : std_logic;
signal \N__57436\ : std_logic;
signal \N__57433\ : std_logic;
signal \N__57430\ : std_logic;
signal \N__57427\ : std_logic;
signal \N__57424\ : std_logic;
signal \N__57421\ : std_logic;
signal \N__57420\ : std_logic;
signal \N__57419\ : std_logic;
signal \N__57416\ : std_logic;
signal \N__57411\ : std_logic;
signal \N__57408\ : std_logic;
signal \N__57405\ : std_logic;
signal \N__57402\ : std_logic;
signal \N__57399\ : std_logic;
signal \N__57396\ : std_logic;
signal \N__57393\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57385\ : std_logic;
signal \N__57384\ : std_logic;
signal \N__57381\ : std_logic;
signal \N__57378\ : std_logic;
signal \N__57375\ : std_logic;
signal \N__57372\ : std_logic;
signal \N__57367\ : std_logic;
signal \N__57364\ : std_logic;
signal \N__57361\ : std_logic;
signal \N__57358\ : std_logic;
signal \N__57355\ : std_logic;
signal \N__57352\ : std_logic;
signal \N__57349\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57343\ : std_logic;
signal \N__57340\ : std_logic;
signal \N__57337\ : std_logic;
signal \N__57334\ : std_logic;
signal \N__57333\ : std_logic;
signal \N__57330\ : std_logic;
signal \N__57327\ : std_logic;
signal \N__57324\ : std_logic;
signal \N__57321\ : std_logic;
signal \N__57316\ : std_logic;
signal \N__57313\ : std_logic;
signal \N__57310\ : std_logic;
signal \N__57307\ : std_logic;
signal \N__57304\ : std_logic;
signal \N__57301\ : std_logic;
signal \N__57298\ : std_logic;
signal \N__57297\ : std_logic;
signal \N__57294\ : std_logic;
signal \N__57291\ : std_logic;
signal \N__57288\ : std_logic;
signal \N__57285\ : std_logic;
signal \N__57280\ : std_logic;
signal \N__57277\ : std_logic;
signal \N__57276\ : std_logic;
signal \N__57273\ : std_logic;
signal \N__57270\ : std_logic;
signal \N__57267\ : std_logic;
signal \N__57264\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57253\ : std_logic;
signal \N__57250\ : std_logic;
signal \N__57247\ : std_logic;
signal \N__57244\ : std_logic;
signal \N__57241\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57235\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57229\ : std_logic;
signal \N__57226\ : std_logic;
signal \N__57223\ : std_logic;
signal \N__57220\ : std_logic;
signal \N__57219\ : std_logic;
signal \N__57216\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57210\ : std_logic;
signal \N__57207\ : std_logic;
signal \N__57202\ : std_logic;
signal \N__57199\ : std_logic;
signal \N__57196\ : std_logic;
signal \N__57195\ : std_logic;
signal \N__57192\ : std_logic;
signal \N__57189\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57183\ : std_logic;
signal \N__57178\ : std_logic;
signal \N__57175\ : std_logic;
signal \N__57172\ : std_logic;
signal \N__57169\ : std_logic;
signal \N__57166\ : std_logic;
signal \N__57163\ : std_logic;
signal \N__57160\ : std_logic;
signal \N__57157\ : std_logic;
signal \N__57154\ : std_logic;
signal \N__57153\ : std_logic;
signal \N__57150\ : std_logic;
signal \N__57147\ : std_logic;
signal \N__57144\ : std_logic;
signal \N__57141\ : std_logic;
signal \N__57136\ : std_logic;
signal \N__57133\ : std_logic;
signal \N__57130\ : std_logic;
signal \N__57127\ : std_logic;
signal \N__57124\ : std_logic;
signal \N__57121\ : std_logic;
signal \N__57118\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57114\ : std_logic;
signal \N__57111\ : std_logic;
signal \N__57108\ : std_logic;
signal \N__57103\ : std_logic;
signal \N__57100\ : std_logic;
signal \N__57097\ : std_logic;
signal \N__57094\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57088\ : std_logic;
signal \N__57085\ : std_logic;
signal \N__57082\ : std_logic;
signal \N__57079\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57070\ : std_logic;
signal \N__57067\ : std_logic;
signal \N__57064\ : std_logic;
signal \N__57061\ : std_logic;
signal \N__57058\ : std_logic;
signal \N__57055\ : std_logic;
signal \N__57052\ : std_logic;
signal \N__57049\ : std_logic;
signal \N__57046\ : std_logic;
signal \N__57043\ : std_logic;
signal \N__57040\ : std_logic;
signal \N__57037\ : std_logic;
signal \N__57034\ : std_logic;
signal \N__57031\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57025\ : std_logic;
signal \N__57022\ : std_logic;
signal \N__57019\ : std_logic;
signal \N__57016\ : std_logic;
signal \N__57013\ : std_logic;
signal \N__57010\ : std_logic;
signal \N__57007\ : std_logic;
signal \N__57004\ : std_logic;
signal \N__57001\ : std_logic;
signal \N__56998\ : std_logic;
signal \N__56995\ : std_logic;
signal \N__56992\ : std_logic;
signal \N__56989\ : std_logic;
signal \N__56986\ : std_logic;
signal \N__56983\ : std_logic;
signal \N__56980\ : std_logic;
signal \N__56977\ : std_logic;
signal \N__56974\ : std_logic;
signal \N__56971\ : std_logic;
signal \N__56968\ : std_logic;
signal \N__56965\ : std_logic;
signal \N__56962\ : std_logic;
signal \N__56959\ : std_logic;
signal \N__56956\ : std_logic;
signal \N__56953\ : std_logic;
signal \N__56950\ : std_logic;
signal \N__56947\ : std_logic;
signal \N__56944\ : std_logic;
signal \N__56941\ : std_logic;
signal \N__56938\ : std_logic;
signal \N__56935\ : std_logic;
signal \N__56932\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56926\ : std_logic;
signal \N__56923\ : std_logic;
signal \N__56920\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56913\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56907\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56896\ : std_logic;
signal \N__56893\ : std_logic;
signal \N__56890\ : std_logic;
signal \N__56887\ : std_logic;
signal \N__56884\ : std_logic;
signal \N__56881\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56872\ : std_logic;
signal \N__56869\ : std_logic;
signal \N__56866\ : std_logic;
signal \N__56863\ : std_logic;
signal \N__56860\ : std_logic;
signal \N__56857\ : std_logic;
signal \N__56854\ : std_logic;
signal \N__56851\ : std_logic;
signal \N__56848\ : std_logic;
signal \N__56845\ : std_logic;
signal \N__56842\ : std_logic;
signal \N__56839\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56833\ : std_logic;
signal \N__56830\ : std_logic;
signal \N__56827\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56821\ : std_logic;
signal \N__56820\ : std_logic;
signal \N__56819\ : std_logic;
signal \N__56818\ : std_logic;
signal \N__56817\ : std_logic;
signal \N__56814\ : std_logic;
signal \N__56813\ : std_logic;
signal \N__56812\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56810\ : std_logic;
signal \N__56809\ : std_logic;
signal \N__56808\ : std_logic;
signal \N__56807\ : std_logic;
signal \N__56806\ : std_logic;
signal \N__56805\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56803\ : std_logic;
signal \N__56802\ : std_logic;
signal \N__56801\ : std_logic;
signal \N__56794\ : std_logic;
signal \N__56785\ : std_logic;
signal \N__56784\ : std_logic;
signal \N__56783\ : std_logic;
signal \N__56782\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56780\ : std_logic;
signal \N__56779\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56775\ : std_logic;
signal \N__56766\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56752\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56740\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56724\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56704\ : std_logic;
signal \N__56701\ : std_logic;
signal \N__56698\ : std_logic;
signal \N__56695\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56689\ : std_logic;
signal \N__56686\ : std_logic;
signal \N__56683\ : std_logic;
signal \N__56680\ : std_logic;
signal \N__56677\ : std_logic;
signal \N__56676\ : std_logic;
signal \N__56671\ : std_logic;
signal \N__56668\ : std_logic;
signal \N__56665\ : std_logic;
signal \N__56662\ : std_logic;
signal \N__56659\ : std_logic;
signal \N__56656\ : std_logic;
signal \N__56653\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56647\ : std_logic;
signal \N__56644\ : std_logic;
signal \N__56641\ : std_logic;
signal \N__56638\ : std_logic;
signal \N__56635\ : std_logic;
signal \N__56632\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56623\ : std_logic;
signal \N__56620\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56614\ : std_logic;
signal \N__56611\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56605\ : std_logic;
signal \N__56602\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56596\ : std_logic;
signal \N__56593\ : std_logic;
signal \N__56590\ : std_logic;
signal \N__56587\ : std_logic;
signal \N__56584\ : std_logic;
signal \N__56581\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56575\ : std_logic;
signal \N__56572\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56566\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56551\ : std_logic;
signal \N__56548\ : std_logic;
signal \N__56545\ : std_logic;
signal \N__56542\ : std_logic;
signal \N__56539\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56533\ : std_logic;
signal \N__56530\ : std_logic;
signal \N__56527\ : std_logic;
signal \N__56524\ : std_logic;
signal \N__56521\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56503\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56497\ : std_logic;
signal \N__56494\ : std_logic;
signal \N__56493\ : std_logic;
signal \N__56492\ : std_logic;
signal \N__56485\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56482\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56479\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56477\ : std_logic;
signal \N__56476\ : std_logic;
signal \N__56473\ : std_logic;
signal \N__56464\ : std_logic;
signal \N__56463\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56461\ : std_logic;
signal \N__56460\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56458\ : std_logic;
signal \N__56457\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56454\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56450\ : std_logic;
signal \N__56449\ : std_logic;
signal \N__56448\ : std_logic;
signal \N__56447\ : std_logic;
signal \N__56444\ : std_logic;
signal \N__56443\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56433\ : std_logic;
signal \N__56428\ : std_logic;
signal \N__56425\ : std_logic;
signal \N__56412\ : std_logic;
signal \N__56399\ : std_logic;
signal \N__56390\ : std_logic;
signal \N__56383\ : std_logic;
signal \N__56368\ : std_logic;
signal \N__56367\ : std_logic;
signal \N__56366\ : std_logic;
signal \N__56365\ : std_logic;
signal \N__56364\ : std_logic;
signal \N__56363\ : std_logic;
signal \N__56362\ : std_logic;
signal \N__56361\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56352\ : std_logic;
signal \N__56349\ : std_logic;
signal \N__56346\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56344\ : std_logic;
signal \N__56343\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56332\ : std_logic;
signal \N__56331\ : std_logic;
signal \N__56330\ : std_logic;
signal \N__56329\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56310\ : std_logic;
signal \N__56309\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56307\ : std_logic;
signal \N__56306\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56303\ : std_logic;
signal \N__56302\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56300\ : std_logic;
signal \N__56299\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56294\ : std_logic;
signal \N__56285\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56251\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56218\ : std_logic;
signal \N__56215\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56211\ : std_logic;
signal \N__56208\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56206\ : std_logic;
signal \N__56205\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56198\ : std_logic;
signal \N__56197\ : std_logic;
signal \N__56194\ : std_logic;
signal \N__56191\ : std_logic;
signal \N__56190\ : std_logic;
signal \N__56189\ : std_logic;
signal \N__56186\ : std_logic;
signal \N__56183\ : std_logic;
signal \N__56182\ : std_logic;
signal \N__56179\ : std_logic;
signal \N__56176\ : std_logic;
signal \N__56173\ : std_logic;
signal \N__56170\ : std_logic;
signal \N__56167\ : std_logic;
signal \N__56164\ : std_logic;
signal \N__56161\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56157\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56151\ : std_logic;
signal \N__56150\ : std_logic;
signal \N__56149\ : std_logic;
signal \N__56148\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56142\ : std_logic;
signal \N__56139\ : std_logic;
signal \N__56136\ : std_logic;
signal \N__56131\ : std_logic;
signal \N__56128\ : std_logic;
signal \N__56125\ : std_logic;
signal \N__56122\ : std_logic;
signal \N__56121\ : std_logic;
signal \N__56116\ : std_logic;
signal \N__56113\ : std_logic;
signal \N__56110\ : std_logic;
signal \N__56107\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56102\ : std_logic;
signal \N__56099\ : std_logic;
signal \N__56098\ : std_logic;
signal \N__56095\ : std_logic;
signal \N__56094\ : std_logic;
signal \N__56091\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56083\ : std_logic;
signal \N__56076\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56042\ : std_logic;
signal \N__56039\ : std_logic;
signal \N__56038\ : std_logic;
signal \N__56035\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56020\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56014\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56004\ : std_logic;
signal \N__55995\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55981\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55972\ : std_logic;
signal \N__55969\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55947\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55945\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55939\ : std_logic;
signal \N__55936\ : std_logic;
signal \N__55933\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55925\ : std_logic;
signal \N__55922\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55918\ : std_logic;
signal \N__55917\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55915\ : std_logic;
signal \N__55912\ : std_logic;
signal \N__55909\ : std_logic;
signal \N__55906\ : std_logic;
signal \N__55903\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55897\ : std_logic;
signal \N__55894\ : std_logic;
signal \N__55891\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55879\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55874\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55866\ : std_logic;
signal \N__55863\ : std_logic;
signal \N__55860\ : std_logic;
signal \N__55849\ : std_logic;
signal \N__55846\ : std_logic;
signal \N__55843\ : std_logic;
signal \N__55840\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55831\ : std_logic;
signal \N__55828\ : std_logic;
signal \N__55827\ : std_logic;
signal \N__55824\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55806\ : std_logic;
signal \N__55803\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55797\ : std_logic;
signal \N__55794\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55774\ : std_logic;
signal \N__55769\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55753\ : std_logic;
signal \N__55750\ : std_logic;
signal \N__55747\ : std_logic;
signal \N__55744\ : std_logic;
signal \N__55741\ : std_logic;
signal \N__55738\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55736\ : std_logic;
signal \N__55733\ : std_logic;
signal \N__55730\ : std_logic;
signal \N__55729\ : std_logic;
signal \N__55726\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55723\ : std_logic;
signal \N__55722\ : std_logic;
signal \N__55719\ : std_logic;
signal \N__55718\ : std_logic;
signal \N__55717\ : std_logic;
signal \N__55714\ : std_logic;
signal \N__55711\ : std_logic;
signal \N__55708\ : std_logic;
signal \N__55705\ : std_logic;
signal \N__55702\ : std_logic;
signal \N__55699\ : std_logic;
signal \N__55698\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55691\ : std_logic;
signal \N__55688\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55679\ : std_logic;
signal \N__55676\ : std_logic;
signal \N__55673\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55664\ : std_logic;
signal \N__55663\ : std_logic;
signal \N__55660\ : std_logic;
signal \N__55659\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55642\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55624\ : std_logic;
signal \N__55621\ : std_logic;
signal \N__55620\ : std_logic;
signal \N__55619\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55617\ : std_logic;
signal \N__55616\ : std_logic;
signal \N__55615\ : std_logic;
signal \N__55612\ : std_logic;
signal \N__55605\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55595\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55586\ : std_logic;
signal \N__55583\ : std_logic;
signal \N__55582\ : std_logic;
signal \N__55579\ : std_logic;
signal \N__55576\ : std_logic;
signal \N__55573\ : std_logic;
signal \N__55570\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55557\ : std_logic;
signal \N__55554\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55519\ : std_logic;
signal \N__55516\ : std_logic;
signal \N__55513\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55511\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55495\ : std_logic;
signal \N__55494\ : std_logic;
signal \N__55493\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55491\ : std_logic;
signal \N__55490\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55488\ : std_logic;
signal \N__55487\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55481\ : std_logic;
signal \N__55472\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55449\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55446\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55416\ : std_logic;
signal \N__55407\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55395\ : std_logic;
signal \N__55390\ : std_logic;
signal \N__55387\ : std_logic;
signal \N__55384\ : std_logic;
signal \N__55381\ : std_logic;
signal \N__55378\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55374\ : std_logic;
signal \N__55371\ : std_logic;
signal \N__55370\ : std_logic;
signal \N__55367\ : std_logic;
signal \N__55366\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55364\ : std_logic;
signal \N__55363\ : std_logic;
signal \N__55360\ : std_logic;
signal \N__55357\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55349\ : std_logic;
signal \N__55348\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55342\ : std_logic;
signal \N__55341\ : std_logic;
signal \N__55338\ : std_logic;
signal \N__55337\ : std_logic;
signal \N__55334\ : std_logic;
signal \N__55331\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55325\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55316\ : std_logic;
signal \N__55313\ : std_logic;
signal \N__55310\ : std_logic;
signal \N__55307\ : std_logic;
signal \N__55306\ : std_logic;
signal \N__55303\ : std_logic;
signal \N__55300\ : std_logic;
signal \N__55297\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55286\ : std_logic;
signal \N__55283\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55275\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55269\ : std_logic;
signal \N__55268\ : std_logic;
signal \N__55267\ : std_logic;
signal \N__55266\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55260\ : std_logic;
signal \N__55253\ : std_logic;
signal \N__55242\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55233\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55216\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55210\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55204\ : std_logic;
signal \N__55189\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55181\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55176\ : std_logic;
signal \N__55173\ : std_logic;
signal \N__55170\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55155\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55150\ : std_logic;
signal \N__55147\ : std_logic;
signal \N__55144\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55138\ : std_logic;
signal \N__55135\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55122\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55106\ : std_logic;
signal \N__55103\ : std_logic;
signal \N__55100\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55094\ : std_logic;
signal \N__55093\ : std_logic;
signal \N__55090\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55084\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55074\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55070\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55060\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55048\ : std_logic;
signal \N__55045\ : std_logic;
signal \N__55042\ : std_logic;
signal \N__55039\ : std_logic;
signal \N__55036\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55032\ : std_logic;
signal \N__55027\ : std_logic;
signal \N__55024\ : std_logic;
signal \N__55021\ : std_logic;
signal \N__55018\ : std_logic;
signal \N__55015\ : std_logic;
signal \N__55012\ : std_logic;
signal \N__55009\ : std_logic;
signal \N__55006\ : std_logic;
signal \N__55005\ : std_logic;
signal \N__55002\ : std_logic;
signal \N__55001\ : std_logic;
signal \N__54998\ : std_logic;
signal \N__54997\ : std_logic;
signal \N__54996\ : std_logic;
signal \N__54993\ : std_logic;
signal \N__54990\ : std_logic;
signal \N__54989\ : std_logic;
signal \N__54988\ : std_logic;
signal \N__54987\ : std_logic;
signal \N__54984\ : std_logic;
signal \N__54981\ : std_logic;
signal \N__54978\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54970\ : std_logic;
signal \N__54969\ : std_logic;
signal \N__54966\ : std_logic;
signal \N__54963\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54952\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54946\ : std_logic;
signal \N__54945\ : std_logic;
signal \N__54942\ : std_logic;
signal \N__54941\ : std_logic;
signal \N__54940\ : std_logic;
signal \N__54935\ : std_logic;
signal \N__54932\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54926\ : std_logic;
signal \N__54923\ : std_logic;
signal \N__54918\ : std_logic;
signal \N__54915\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54902\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54886\ : std_logic;
signal \N__54883\ : std_logic;
signal \N__54880\ : std_logic;
signal \N__54873\ : std_logic;
signal \N__54862\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54856\ : std_logic;
signal \N__54853\ : std_logic;
signal \N__54850\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54844\ : std_logic;
signal \N__54841\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54826\ : std_logic;
signal \N__54823\ : std_logic;
signal \N__54820\ : std_logic;
signal \N__54817\ : std_logic;
signal \N__54814\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54805\ : std_logic;
signal \N__54804\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54802\ : std_logic;
signal \N__54801\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54799\ : std_logic;
signal \N__54798\ : std_logic;
signal \N__54797\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54793\ : std_logic;
signal \N__54790\ : std_logic;
signal \N__54787\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54781\ : std_logic;
signal \N__54778\ : std_logic;
signal \N__54775\ : std_logic;
signal \N__54774\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54772\ : std_logic;
signal \N__54771\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54769\ : std_logic;
signal \N__54768\ : std_logic;
signal \N__54765\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54761\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54742\ : std_logic;
signal \N__54739\ : std_logic;
signal \N__54736\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54730\ : std_logic;
signal \N__54727\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54721\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54715\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54713\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54705\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54699\ : std_logic;
signal \N__54696\ : std_logic;
signal \N__54681\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54675\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54665\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54650\ : std_logic;
signal \N__54637\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54629\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54577\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54565\ : std_logic;
signal \N__54562\ : std_logic;
signal \N__54559\ : std_logic;
signal \N__54556\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54547\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54530\ : std_logic;
signal \N__54527\ : std_logic;
signal \N__54526\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54521\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54513\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54500\ : std_logic;
signal \N__54499\ : std_logic;
signal \N__54498\ : std_logic;
signal \N__54497\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54491\ : std_logic;
signal \N__54488\ : std_logic;
signal \N__54485\ : std_logic;
signal \N__54482\ : std_logic;
signal \N__54481\ : std_logic;
signal \N__54480\ : std_logic;
signal \N__54477\ : std_logic;
signal \N__54474\ : std_logic;
signal \N__54473\ : std_logic;
signal \N__54470\ : std_logic;
signal \N__54469\ : std_logic;
signal \N__54466\ : std_logic;
signal \N__54463\ : std_logic;
signal \N__54460\ : std_logic;
signal \N__54457\ : std_logic;
signal \N__54454\ : std_logic;
signal \N__54451\ : std_logic;
signal \N__54450\ : std_logic;
signal \N__54449\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54445\ : std_logic;
signal \N__54442\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54437\ : std_logic;
signal \N__54434\ : std_logic;
signal \N__54433\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54411\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54397\ : std_logic;
signal \N__54390\ : std_logic;
signal \N__54387\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54383\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54365\ : std_logic;
signal \N__54362\ : std_logic;
signal \N__54355\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54349\ : std_logic;
signal \N__54344\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54333\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54317\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54300\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54286\ : std_logic;
signal \N__54283\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54268\ : std_logic;
signal \N__54265\ : std_logic;
signal \N__54264\ : std_logic;
signal \N__54261\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54257\ : std_logic;
signal \N__54256\ : std_logic;
signal \N__54255\ : std_logic;
signal \N__54254\ : std_logic;
signal \N__54253\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54251\ : std_logic;
signal \N__54250\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54248\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54242\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54233\ : std_logic;
signal \N__54232\ : std_logic;
signal \N__54229\ : std_logic;
signal \N__54228\ : std_logic;
signal \N__54225\ : std_logic;
signal \N__54224\ : std_logic;
signal \N__54221\ : std_logic;
signal \N__54220\ : std_logic;
signal \N__54217\ : std_logic;
signal \N__54214\ : std_logic;
signal \N__54211\ : std_logic;
signal \N__54208\ : std_logic;
signal \N__54207\ : std_logic;
signal \N__54202\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54196\ : std_logic;
signal \N__54195\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54193\ : std_logic;
signal \N__54190\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54166\ : std_logic;
signal \N__54163\ : std_logic;
signal \N__54160\ : std_logic;
signal \N__54157\ : std_logic;
signal \N__54156\ : std_logic;
signal \N__54153\ : std_logic;
signal \N__54148\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54137\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54132\ : std_logic;
signal \N__54129\ : std_logic;
signal \N__54126\ : std_logic;
signal \N__54123\ : std_logic;
signal \N__54120\ : std_logic;
signal \N__54111\ : std_logic;
signal \N__54108\ : std_logic;
signal \N__54105\ : std_logic;
signal \N__54100\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54084\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54080\ : std_logic;
signal \N__54077\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54055\ : std_logic;
signal \N__54046\ : std_logic;
signal \N__54043\ : std_logic;
signal \N__54038\ : std_logic;
signal \N__54033\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54016\ : std_logic;
signal \N__54013\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54004\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__54000\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53992\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53971\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53955\ : std_logic;
signal \N__53952\ : std_logic;
signal \N__53949\ : std_logic;
signal \N__53946\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53941\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53937\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53915\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53907\ : std_logic;
signal \N__53904\ : std_logic;
signal \N__53903\ : std_logic;
signal \N__53900\ : std_logic;
signal \N__53897\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53887\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53883\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53876\ : std_logic;
signal \N__53873\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53867\ : std_logic;
signal \N__53854\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53836\ : std_logic;
signal \N__53833\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53826\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53802\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53775\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53743\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53734\ : std_logic;
signal \N__53731\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53725\ : std_logic;
signal \N__53724\ : std_logic;
signal \N__53723\ : std_logic;
signal \N__53722\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53716\ : std_logic;
signal \N__53715\ : std_logic;
signal \N__53712\ : std_logic;
signal \N__53711\ : std_logic;
signal \N__53708\ : std_logic;
signal \N__53707\ : std_logic;
signal \N__53706\ : std_logic;
signal \N__53705\ : std_logic;
signal \N__53702\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53693\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53687\ : std_logic;
signal \N__53684\ : std_logic;
signal \N__53681\ : std_logic;
signal \N__53680\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53665\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53661\ : std_logic;
signal \N__53658\ : std_logic;
signal \N__53657\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53651\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53644\ : std_logic;
signal \N__53641\ : std_logic;
signal \N__53638\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53625\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53611\ : std_logic;
signal \N__53610\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53608\ : std_logic;
signal \N__53607\ : std_logic;
signal \N__53604\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53592\ : std_logic;
signal \N__53589\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53582\ : std_logic;
signal \N__53575\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53569\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53567\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53563\ : std_logic;
signal \N__53560\ : std_logic;
signal \N__53559\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53544\ : std_logic;
signal \N__53541\ : std_logic;
signal \N__53534\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53516\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53508\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53488\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53478\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53471\ : std_logic;
signal \N__53470\ : std_logic;
signal \N__53469\ : std_logic;
signal \N__53468\ : std_logic;
signal \N__53467\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53465\ : std_logic;
signal \N__53464\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53452\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53434\ : std_logic;
signal \N__53431\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53429\ : std_logic;
signal \N__53428\ : std_logic;
signal \N__53427\ : std_logic;
signal \N__53426\ : std_logic;
signal \N__53423\ : std_logic;
signal \N__53420\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53382\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53378\ : std_logic;
signal \N__53377\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53373\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53369\ : std_logic;
signal \N__53364\ : std_logic;
signal \N__53359\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53353\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53347\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53323\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53317\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53297\ : std_logic;
signal \N__53288\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53284\ : std_logic;
signal \N__53281\ : std_logic;
signal \N__53278\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53262\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53251\ : std_logic;
signal \N__53248\ : std_logic;
signal \N__53245\ : std_logic;
signal \N__53242\ : std_logic;
signal \N__53239\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53227\ : std_logic;
signal \N__53224\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53215\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53210\ : std_logic;
signal \N__53207\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53203\ : std_logic;
signal \N__53202\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53198\ : std_logic;
signal \N__53197\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53191\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53186\ : std_logic;
signal \N__53183\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53171\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53169\ : std_logic;
signal \N__53166\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53158\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53151\ : std_logic;
signal \N__53148\ : std_logic;
signal \N__53147\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53072\ : std_logic;
signal \N__53069\ : std_logic;
signal \N__53066\ : std_logic;
signal \N__53059\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52945\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52929\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52912\ : std_logic;
signal \N__52909\ : std_logic;
signal \N__52906\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52867\ : std_logic;
signal \N__52864\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52843\ : std_logic;
signal \N__52842\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52828\ : std_logic;
signal \N__52825\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52819\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52804\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52789\ : std_logic;
signal \N__52786\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52773\ : std_logic;
signal \N__52772\ : std_logic;
signal \N__52767\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52756\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52750\ : std_logic;
signal \N__52747\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52729\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52687\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52681\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52657\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52645\ : std_logic;
signal \N__52642\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52582\ : std_logic;
signal \N__52579\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52569\ : std_logic;
signal \N__52566\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52537\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52516\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52510\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52501\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52492\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52363\ : std_logic;
signal \N__52360\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52354\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52341\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52333\ : std_logic;
signal \N__52330\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52324\ : std_logic;
signal \N__52321\ : std_logic;
signal \N__52318\ : std_logic;
signal \N__52315\ : std_logic;
signal \N__52312\ : std_logic;
signal \N__52309\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52273\ : std_logic;
signal \N__52270\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52252\ : std_logic;
signal \N__52249\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52219\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52204\ : std_logic;
signal \N__52201\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52180\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52129\ : std_logic;
signal \N__52126\ : std_logic;
signal \N__52123\ : std_logic;
signal \N__52120\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52056\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51988\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51949\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51925\ : std_logic;
signal \N__51922\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51877\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51850\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51844\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51835\ : std_logic;
signal \N__51832\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51799\ : std_logic;
signal \N__51796\ : std_logic;
signal \N__51793\ : std_logic;
signal \N__51790\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51745\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51736\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51709\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51694\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51628\ : std_logic;
signal \N__51625\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51511\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51385\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51376\ : std_logic;
signal \N__51373\ : std_logic;
signal \N__51370\ : std_logic;
signal \N__51367\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51337\ : std_logic;
signal \N__51334\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51325\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51274\ : std_logic;
signal \N__51271\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51160\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51146\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51140\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51116\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51061\ : std_logic;
signal \N__51058\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51035\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51018\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51008\ : std_logic;
signal \N__51005\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50959\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50926\ : std_logic;
signal \N__50923\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50890\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50862\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50842\ : std_logic;
signal \N__50839\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50812\ : std_logic;
signal \N__50809\ : std_logic;
signal \N__50806\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50671\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50503\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49258\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48028\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45325\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal pin3_clk_16mhz_pad_gb_input : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_6_20_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17336\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8176\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8175\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8174\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8173\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8172\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17349\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8177\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17448\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8490\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2338\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2438\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2538\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2638\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2738\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2838\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2938\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3038\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17458\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3138\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252\ : std_logic;
signal \bfn_7_23_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17478\ : std_logic;
signal \bfn_7_24_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2341\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2344\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2441\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2444\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2541\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2544\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2641\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2644\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2741\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2744\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2841\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2844\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2941\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2944\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3041\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17468\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3044\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3141\ : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3144\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \foc.u_Park_Transform.n17107\ : std_logic;
signal \foc.u_Park_Transform.n17108\ : std_logic;
signal \foc.u_Park_Transform.n17109\ : std_logic;
signal \foc.u_Park_Transform.n17110\ : std_logic;
signal \foc.u_Park_Transform.n17111\ : std_logic;
signal \foc.u_Park_Transform.n17112\ : std_logic;
signal \foc.u_Park_Transform.n17113\ : std_logic;
signal \foc.u_Park_Transform.n17114\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \foc.u_Park_Transform.n17115\ : std_logic;
signal \foc.u_Park_Transform.n17116\ : std_logic;
signal \foc.u_Park_Transform.n779_adj_2070\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n81\ : std_logic;
signal \foc.u_Park_Transform.n17118\ : std_logic;
signal \foc.u_Park_Transform.n130\ : std_logic;
signal \foc.u_Park_Transform.n17119\ : std_logic;
signal \foc.u_Park_Transform.n179\ : std_logic;
signal \foc.u_Park_Transform.n17120\ : std_logic;
signal \foc.u_Park_Transform.n228_adj_2063\ : std_logic;
signal \foc.u_Park_Transform.n17121\ : std_logic;
signal \foc.u_Park_Transform.n277_adj_2060\ : std_logic;
signal \foc.u_Park_Transform.n17122\ : std_logic;
signal \foc.u_Park_Transform.n326_adj_2056\ : std_logic;
signal \foc.u_Park_Transform.n17123\ : std_logic;
signal \foc.u_Park_Transform.n375_adj_2055\ : std_logic;
signal \foc.u_Park_Transform.n17124\ : std_logic;
signal \foc.u_Park_Transform.n17125\ : std_logic;
signal \foc.u_Park_Transform.n424_adj_2052\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n473_adj_2050\ : std_logic;
signal \foc.u_Park_Transform.n17126\ : std_logic;
signal \foc.u_Park_Transform.n17127\ : std_logic;
signal \foc.u_Park_Transform.n17128\ : std_logic;
signal \foc.u_Park_Transform.n522_adj_2046\ : std_logic;
signal \foc.u_Park_Transform.n17129\ : std_logic;
signal \foc.u_Park_Transform.n775_adj_2047\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n16935\ : std_logic;
signal \foc.u_Park_Transform.n16936\ : std_logic;
signal \foc.u_Park_Transform.n16937\ : std_logic;
signal \foc.u_Park_Transform.n16938\ : std_logic;
signal \foc.u_Park_Transform.n16939\ : std_logic;
signal \foc.u_Park_Transform.n16940\ : std_logic;
signal \foc.u_Park_Transform.n16941\ : std_logic;
signal \foc.u_Park_Transform.n16942\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n16943\ : std_logic;
signal \foc.u_Park_Transform.n16944\ : std_logic;
signal \foc.u_Park_Transform.n16945\ : std_logic;
signal \foc.u_Park_Transform.n16946\ : std_logic;
signal \foc.u_Park_Transform.n775\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15467\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2834\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15471\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2335\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2435\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2535\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2635\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2735\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2835\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2935\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17438\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3035\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3135\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7897\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7896\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7895\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7894\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7893\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7892\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7891\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17343\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2347\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7473\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2447\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2547\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2647\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2747\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2847\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2947\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3047\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17488\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3147\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17489\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \foc.u_Park_Transform.n17146\ : std_logic;
signal \foc.u_Park_Transform.n17147\ : std_logic;
signal \foc.u_Park_Transform.n17148\ : std_logic;
signal \foc.u_Park_Transform.n17149\ : std_logic;
signal \foc.u_Park_Transform.n17150\ : std_logic;
signal \foc.u_Park_Transform.n17151\ : std_logic;
signal \foc.u_Park_Transform.n17152\ : std_logic;
signal \foc.u_Park_Transform.n17153\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \foc.u_Park_Transform.n17154\ : std_logic;
signal \foc.u_Park_Transform.n17155\ : std_logic;
signal \foc.u_Park_Transform.n17156\ : std_logic;
signal \foc.u_Park_Transform.n17157\ : std_logic;
signal \foc.u_Park_Transform.n17158\ : std_logic;
signal \foc.u_Park_Transform.n17159\ : std_logic;
signal \foc.u_Park_Transform.n767\ : std_logic;
signal \foc.u_Park_Transform.n75\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n78\ : std_logic;
signal \foc.u_Park_Transform.n124\ : std_logic;
signal \foc.u_Park_Transform.n17131\ : std_logic;
signal \foc.u_Park_Transform.n127\ : std_logic;
signal \foc.u_Park_Transform.n173\ : std_logic;
signal \foc.u_Park_Transform.n17132\ : std_logic;
signal \foc.u_Park_Transform.n176\ : std_logic;
signal \foc.u_Park_Transform.n222\ : std_logic;
signal \foc.u_Park_Transform.n17133\ : std_logic;
signal \foc.u_Park_Transform.n225\ : std_logic;
signal \foc.u_Park_Transform.n271\ : std_logic;
signal \foc.u_Park_Transform.n17134\ : std_logic;
signal \foc.u_Park_Transform.n274\ : std_logic;
signal \foc.u_Park_Transform.n320\ : std_logic;
signal \foc.u_Park_Transform.n17135\ : std_logic;
signal \foc.u_Park_Transform.n323\ : std_logic;
signal \foc.u_Park_Transform.n369\ : std_logic;
signal \foc.u_Park_Transform.n17136\ : std_logic;
signal \foc.u_Park_Transform.n372\ : std_logic;
signal \foc.u_Park_Transform.n418_adj_2024\ : std_logic;
signal \foc.u_Park_Transform.n17137\ : std_logic;
signal \foc.u_Park_Transform.n17138\ : std_logic;
signal \foc.u_Park_Transform.n421_adj_2039\ : std_logic;
signal \foc.u_Park_Transform.n467_adj_2019\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n470_adj_2038\ : std_logic;
signal \foc.u_Park_Transform.n516_adj_2018\ : std_logic;
signal \foc.u_Park_Transform.n17139\ : std_logic;
signal \foc.u_Park_Transform.n519_adj_2035\ : std_logic;
signal \foc.u_Park_Transform.n565\ : std_logic;
signal \foc.u_Park_Transform.n17140\ : std_logic;
signal \foc.u_Park_Transform.n568_adj_2034\ : std_logic;
signal \foc.u_Park_Transform.n614_adj_2017\ : std_logic;
signal \foc.u_Park_Transform.n17141\ : std_logic;
signal \foc.u_Park_Transform.n663_adj_2016\ : std_logic;
signal \foc.u_Park_Transform.n17142\ : std_logic;
signal \foc.u_Park_Transform.n712_adj_2015\ : std_logic;
signal \foc.u_Park_Transform.n17143\ : std_logic;
signal \foc.u_Park_Transform.n617_adj_2031\ : std_logic;
signal \foc.u_Park_Transform.n17144\ : std_logic;
signal \foc.u_Park_Transform.n771_adj_2032\ : std_logic;
signal \foc.u_Park_Transform.n773\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \foc.u_Park_Transform.n18160\ : std_logic;
signal \foc.u_Park_Transform.n18161\ : std_logic;
signal \foc.u_Park_Transform.n18162\ : std_logic;
signal \foc.u_Park_Transform.n18163\ : std_logic;
signal \foc.u_Park_Transform.n18164\ : std_logic;
signal \foc.u_Park_Transform.n18165\ : std_logic;
signal \foc.u_Park_Transform.n787\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n87\ : std_logic;
signal \foc.u_Park_Transform.n16915\ : std_logic;
signal \foc.u_Park_Transform.n136\ : std_logic;
signal \foc.u_Park_Transform.n16916\ : std_logic;
signal \foc.u_Park_Transform.n185\ : std_logic;
signal \foc.u_Park_Transform.n16917\ : std_logic;
signal \foc.u_Park_Transform.n234\ : std_logic;
signal \foc.u_Park_Transform.n16918\ : std_logic;
signal \foc.u_Park_Transform.n283\ : std_logic;
signal \foc.u_Park_Transform.n16919\ : std_logic;
signal \foc.u_Park_Transform.n16920\ : std_logic;
signal \foc.u_Park_Transform.n16921\ : std_logic;
signal \foc.u_Park_Transform.n16922\ : std_logic;
signal \foc.u_Park_Transform.n332\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n783_adj_2167\ : std_logic;
signal \foc.u_Park_Transform.n81_adj_2120\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \foc.u_Park_Transform.n84_adj_2118\ : std_logic;
signal \foc.u_Park_Transform.n130_adj_2105\ : std_logic;
signal \foc.u_Park_Transform.n16924\ : std_logic;
signal \foc.u_Park_Transform.n133\ : std_logic;
signal \foc.u_Park_Transform.n179_adj_2076\ : std_logic;
signal \foc.u_Park_Transform.n16925\ : std_logic;
signal \foc.u_Park_Transform.n182\ : std_logic;
signal \foc.u_Park_Transform.n228\ : std_logic;
signal \foc.u_Park_Transform.n16926\ : std_logic;
signal \foc.u_Park_Transform.n231\ : std_logic;
signal \foc.u_Park_Transform.n277\ : std_logic;
signal \foc.u_Park_Transform.n16927\ : std_logic;
signal \foc.u_Park_Transform.n280\ : std_logic;
signal \foc.u_Park_Transform.n326\ : std_logic;
signal \foc.u_Park_Transform.n16928\ : std_logic;
signal \foc.u_Park_Transform.n329\ : std_logic;
signal \foc.u_Park_Transform.n375\ : std_logic;
signal \foc.u_Park_Transform.n16929\ : std_logic;
signal \foc.u_Park_Transform.n378\ : std_logic;
signal \foc.u_Park_Transform.n424\ : std_logic;
signal \foc.u_Park_Transform.n16930\ : std_logic;
signal \foc.u_Park_Transform.n16931\ : std_logic;
signal \foc.u_Park_Transform.n473\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \foc.u_Park_Transform.n619\ : std_logic;
signal \foc.u_Park_Transform.n522\ : std_logic;
signal \foc.u_Park_Transform.n16932\ : std_logic;
signal \foc.u_Park_Transform.n777\ : std_logic;
signal \foc.u_Park_Transform.n427\ : std_logic;
signal \foc.u_Park_Transform.n16933\ : std_logic;
signal \foc.u_Park_Transform.n779\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17392\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2332\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2432\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2532\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2632\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2732\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2832\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2932\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17428\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3032\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2828\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3132\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2420\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2520\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2620\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2720\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2820\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2920\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3020\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3120\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17401\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7554\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7472\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7553\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7471\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7552\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7470\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7551\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7469\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7550\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7468\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7549\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7467\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7548\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7466\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17357\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7547\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\ : std_logic;
signal \bfn_10_26_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7465\ : std_logic;
signal \foc.u_Park_Transform.n84\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \foc.u_Park_Transform.n133_adj_2101\ : std_logic;
signal \foc.u_Park_Transform.n17098\ : std_logic;
signal \foc.u_Park_Transform.n182_adj_2094\ : std_logic;
signal \foc.u_Park_Transform.n17099\ : std_logic;
signal \foc.u_Park_Transform.n231_adj_2089\ : std_logic;
signal \foc.u_Park_Transform.n17100\ : std_logic;
signal \foc.u_Park_Transform.n280_adj_2087\ : std_logic;
signal \foc.u_Park_Transform.n17101\ : std_logic;
signal \foc.u_Park_Transform.n329_adj_2080\ : std_logic;
signal \foc.u_Park_Transform.n17102\ : std_logic;
signal \foc.u_Park_Transform.n378_adj_2078\ : std_logic;
signal \foc.u_Park_Transform.n17103\ : std_logic;
signal \foc.u_Park_Transform.n427_adj_2069\ : std_logic;
signal \foc.u_Park_Transform.n17104\ : std_logic;
signal \foc.u_Park_Transform.n17105\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \foc.u_Park_Transform.n783\ : std_logic;
signal \foc.u_Park_Transform.n622\ : std_logic;
signal \foc.u_Park_Transform.n781\ : std_logic;
signal \foc.u_Park_Transform.n87_adj_2138\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n136_adj_2127\ : std_logic;
signal \foc.u_Park_Transform.n17980\ : std_logic;
signal \foc.u_Park_Transform.n185_adj_2126\ : std_logic;
signal \foc.u_Park_Transform.n17981\ : std_logic;
signal \foc.u_Park_Transform.n234_adj_2125\ : std_logic;
signal \foc.u_Park_Transform.n17982\ : std_logic;
signal \foc.u_Park_Transform.n283_adj_2122\ : std_logic;
signal \foc.u_Park_Transform.n17983\ : std_logic;
signal \foc.u_Park_Transform.n332_adj_2110\ : std_logic;
signal \foc.u_Park_Transform.n17984\ : std_logic;
signal \foc.u_Park_Transform.n17985\ : std_logic;
signal \foc.u_Park_Transform.n787_adj_2149\ : std_logic;
signal \foc.u_Park_Transform.n625\ : std_logic;
signal \n21486_cascade_\ : std_logic;
signal n139 : std_logic;
signal \foc.u_Park_Transform.n90\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946\ : std_logic;
signal \foc.Look_Up_Table_out1_1_6\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947\ : std_logic;
signal \foc.Look_Up_Table_out1_1_7\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948\ : std_logic;
signal \foc.Look_Up_Table_out1_1_8\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949\ : std_logic;
signal \foc.Look_Up_Table_out1_1_9\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15951\ : std_logic;
signal \foc.Look_Up_Table_out1_1_10\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \foc.Look_Up_Table_out1_1_11\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15956\ : std_logic;
signal \foc.Look_Up_Table_out1_1_12\ : std_logic;
signal \foc.u_Park_Transform.n785\ : std_logic;
signal \foc.u_Park_Transform.n616\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n78_adj_2145\ : std_logic;
signal \foc.u_Park_Transform.n16948\ : std_logic;
signal \foc.u_Park_Transform.n127_adj_2119\ : std_logic;
signal \foc.u_Park_Transform.n16949\ : std_logic;
signal \foc.u_Park_Transform.n176_adj_2104\ : std_logic;
signal \foc.u_Park_Transform.n16950\ : std_logic;
signal \foc.u_Park_Transform.n225_adj_2075\ : std_logic;
signal \foc.u_Park_Transform.n16951\ : std_logic;
signal \foc.u_Park_Transform.n274_adj_2058\ : std_logic;
signal \foc.u_Park_Transform.n16952\ : std_logic;
signal \foc.u_Park_Transform.n323_adj_2057\ : std_logic;
signal \foc.u_Park_Transform.n16953\ : std_logic;
signal \foc.u_Park_Transform.n372_adj_2042\ : std_logic;
signal \foc.u_Park_Transform.n16954\ : std_logic;
signal \foc.u_Park_Transform.n16955\ : std_logic;
signal \foc.u_Park_Transform.n421\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n470\ : std_logic;
signal \foc.u_Park_Transform.n16956\ : std_logic;
signal \foc.u_Park_Transform.n519\ : std_logic;
signal \foc.u_Park_Transform.n16957\ : std_logic;
signal \foc.u_Park_Transform.n568\ : std_logic;
signal \foc.u_Park_Transform.n16958\ : std_logic;
signal \foc.u_Park_Transform.n16959\ : std_logic;
signal \foc.u_Park_Transform.n16960\ : std_logic;
signal \foc.u_Park_Transform.n769\ : std_logic;
signal \foc.u_Park_Transform.n617\ : std_logic;
signal \foc.u_Park_Transform.n16961\ : std_logic;
signal \foc.u_Park_Transform.n771\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17358\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17359\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17360\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17361\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17362\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2807\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17365\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3008\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3108\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3211\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_34\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_35\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_36\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3223\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_37\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3227\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_38\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_39\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17497\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_40\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3239\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_41\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3243\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_42\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3247\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_43\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3251\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_44\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3255\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_45\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3259\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_46\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3263\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17504\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_47\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2329\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2429\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2529\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2629\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2729\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2829\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2929\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3029\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17419\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3129\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3235\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2825\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2423\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2426\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2523\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2526\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2623\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2626\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2723\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2726\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2823\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2826\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2923\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2926\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3023\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3026\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3123\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17410\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3126\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3231\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_CO\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \foc.u_Park_Transform.n72\ : std_logic;
signal \foc.u_Park_Transform.n17161\ : std_logic;
signal \foc.u_Park_Transform.n121\ : std_logic;
signal \foc.u_Park_Transform.n17162\ : std_logic;
signal \foc.u_Park_Transform.n170\ : std_logic;
signal \foc.u_Park_Transform.n17163\ : std_logic;
signal \foc.u_Park_Transform.n219\ : std_logic;
signal \foc.u_Park_Transform.n17164\ : std_logic;
signal \foc.u_Park_Transform.n268\ : std_logic;
signal \foc.u_Park_Transform.n17165\ : std_logic;
signal \foc.u_Park_Transform.n317\ : std_logic;
signal \foc.u_Park_Transform.n17166\ : std_logic;
signal \foc.u_Park_Transform.n366\ : std_logic;
signal \foc.u_Park_Transform.n17167\ : std_logic;
signal \foc.u_Park_Transform.n17168\ : std_logic;
signal \foc.u_Park_Transform.n415_adj_2008\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \foc.u_Park_Transform.n464_adj_2005\ : std_logic;
signal \foc.u_Park_Transform.n17169\ : std_logic;
signal \foc.u_Park_Transform.n513_adj_2002\ : std_logic;
signal \foc.u_Park_Transform.n17170\ : std_logic;
signal \foc.u_Park_Transform.n562_adj_2000\ : std_logic;
signal \foc.u_Park_Transform.n17171\ : std_logic;
signal \foc.u_Park_Transform.n611\ : std_logic;
signal \foc.u_Park_Transform.n17172\ : std_logic;
signal \foc.u_Park_Transform.n660\ : std_logic;
signal \foc.u_Park_Transform.n17173\ : std_logic;
signal \foc.u_Park_Transform.n709\ : std_logic;
signal \foc.u_Park_Transform.n17174\ : std_logic;
signal \foc.u_Park_Transform.n763\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n69\ : std_logic;
signal \foc.u_Park_Transform.n17176\ : std_logic;
signal \foc.u_Park_Transform.n118\ : std_logic;
signal \foc.u_Park_Transform.n17177\ : std_logic;
signal \foc.u_Park_Transform.n167\ : std_logic;
signal \foc.u_Park_Transform.n17178\ : std_logic;
signal \foc.u_Park_Transform.n216\ : std_logic;
signal \foc.u_Park_Transform.n17179\ : std_logic;
signal \foc.u_Park_Transform.n265\ : std_logic;
signal \foc.u_Park_Transform.n17180\ : std_logic;
signal \foc.u_Park_Transform.n314\ : std_logic;
signal \foc.u_Park_Transform.n17181\ : std_logic;
signal \foc.u_Park_Transform.n363\ : std_logic;
signal \foc.u_Park_Transform.n17182\ : std_logic;
signal \foc.u_Park_Transform.n17183\ : std_logic;
signal \foc.u_Park_Transform.n412\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n461\ : std_logic;
signal \foc.u_Park_Transform.n17184\ : std_logic;
signal \foc.u_Park_Transform.n510_adj_2004\ : std_logic;
signal \foc.u_Park_Transform.n17185\ : std_logic;
signal \foc.u_Park_Transform.n559_adj_2001\ : std_logic;
signal \foc.u_Park_Transform.n17186\ : std_logic;
signal \foc.u_Park_Transform.n608\ : std_logic;
signal \foc.u_Park_Transform.n17187\ : std_logic;
signal \foc.u_Park_Transform.n657\ : std_logic;
signal \foc.u_Park_Transform.n17188\ : std_logic;
signal \foc.u_Park_Transform.n706\ : std_logic;
signal \foc.u_Park_Transform.n17189\ : std_logic;
signal \foc.u_Park_Transform.n759_adj_2166\ : std_logic;
signal \foc.Look_Up_Table_out1_1_3\ : std_logic;
signal \foc.Look_Up_Table_out1_1_5\ : std_logic;
signal \foc.Look_Up_Table_out1_1_4\ : std_logic;
signal \n4_cascade_\ : std_logic;
signal \foc.u_Park_Transform.n237\ : std_logic;
signal \foc.u_Park_Transform.n188\ : std_logic;
signal \foc.u_Park_Transform.n613\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n75_adj_2123\ : std_logic;
signal \foc.u_Park_Transform.n16963\ : std_logic;
signal \foc.u_Park_Transform.n124_adj_2090\ : std_logic;
signal \foc.u_Park_Transform.n16964\ : std_logic;
signal \foc.u_Park_Transform.n173_adj_2061\ : std_logic;
signal \foc.u_Park_Transform.n16965\ : std_logic;
signal \foc.u_Park_Transform.n222_adj_2049\ : std_logic;
signal \foc.u_Park_Transform.n16966\ : std_logic;
signal \foc.u_Park_Transform.n271_adj_2043\ : std_logic;
signal \foc.u_Park_Transform.n16967\ : std_logic;
signal \foc.u_Park_Transform.n320_adj_2036\ : std_logic;
signal \foc.u_Park_Transform.n16968\ : std_logic;
signal \foc.u_Park_Transform.n369_adj_2026\ : std_logic;
signal \foc.u_Park_Transform.n16969\ : std_logic;
signal \foc.u_Park_Transform.n16970\ : std_logic;
signal \foc.u_Park_Transform.n418\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n467\ : std_logic;
signal \foc.u_Park_Transform.n16971\ : std_logic;
signal \foc.u_Park_Transform.n516\ : std_logic;
signal \foc.u_Park_Transform.n16972\ : std_logic;
signal \foc.u_Park_Transform.n565_adj_2020\ : std_logic;
signal \foc.u_Park_Transform.n16973\ : std_logic;
signal \foc.u_Park_Transform.n614\ : std_logic;
signal \foc.u_Park_Transform.n16974\ : std_logic;
signal \foc.u_Park_Transform.n663\ : std_logic;
signal \foc.u_Park_Transform.n16975\ : std_logic;
signal \foc.u_Park_Transform.n765\ : std_logic;
signal \foc.u_Park_Transform.n712\ : std_logic;
signal \foc.u_Park_Transform.n16976\ : std_logic;
signal \foc.u_Park_Transform.n767_adj_2041\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \foc.u_Park_Transform.n16900\ : std_logic;
signal \foc.u_Park_Transform.n16901\ : std_logic;
signal \foc.u_Park_Transform.n16902\ : std_logic;
signal \foc.u_Park_Transform.n16903\ : std_logic;
signal \foc.u_Park_Transform.n16904\ : std_logic;
signal \foc.u_Park_Transform.n16905\ : std_logic;
signal \foc.u_Park_Transform.n16906\ : std_logic;
signal \foc.u_Park_Transform.n16907\ : std_logic;
signal \foc.u_Park_Transform.n766_adj_2053\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \foc.u_Park_Transform.n770\ : std_logic;
signal \foc.u_Park_Transform.n767_adj_2041_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n16908\ : std_logic;
signal \foc.u_Park_Transform.n774\ : std_logic;
signal \foc.u_Park_Transform.n771_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n16909\ : std_logic;
signal \foc.u_Park_Transform.n778\ : std_logic;
signal \foc.u_Park_Transform.n775_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n16910\ : std_logic;
signal \foc.u_Park_Transform.n782\ : std_logic;
signal \foc.u_Park_Transform.n779_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n16911\ : std_logic;
signal \foc.u_Park_Transform.n786\ : std_logic;
signal \foc.u_Park_Transform.n783_adj_2167_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n16912\ : std_logic;
signal \foc.u_Park_Transform.n787_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n16913\ : std_logic;
signal \foc.u_Park_Transform.n16914\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2417\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2517\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2617\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2717\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2817\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2917\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3017\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17383\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3117\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3219\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_CO\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17656\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17657\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17658\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17659\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17660\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17661\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17662\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17663\ : std_logic;
signal \bfn_12_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17664\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17665\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17666\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17667\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n775\ : std_logic;
signal \bfn_12_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n78_adj_617\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18107\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n127_adj_615\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18108\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n176_adj_613\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18109\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n225_adj_611\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18110\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n274_adj_609\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18111\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n323_adj_607\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18112\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n372\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18113\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18114\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n421\ : std_logic;
signal \bfn_12_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n470\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18115\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n519\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18116\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n568\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18117\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18118\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18119\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n617\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18120\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \foc.u_Park_Transform.n17083\ : std_logic;
signal \foc.u_Park_Transform.n17084\ : std_logic;
signal \foc.u_Park_Transform.n17085\ : std_logic;
signal \foc.u_Park_Transform.n17086\ : std_logic;
signal \foc.u_Park_Transform.n17087\ : std_logic;
signal \foc.u_Park_Transform.n758_adj_2168\ : std_logic;
signal \foc.u_Park_Transform.n17088\ : std_logic;
signal \foc.u_Park_Transform.n759_adj_2166_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n762\ : std_logic;
signal \foc.u_Park_Transform.n17089\ : std_logic;
signal \foc.u_Park_Transform.n17090\ : std_logic;
signal \foc.u_Park_Transform.n766\ : std_logic;
signal \foc.u_Park_Transform.n763_THRU_CO\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \foc.u_Park_Transform.n770_adj_2030\ : std_logic;
signal \foc.u_Park_Transform.n767_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n17091\ : std_logic;
signal \foc.u_Park_Transform.n774_adj_2045\ : std_logic;
signal \foc.u_Park_Transform.n771_adj_2032_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n17092\ : std_logic;
signal \foc.u_Park_Transform.n778_adj_2068\ : std_logic;
signal \foc.u_Park_Transform.n775_adj_2047_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n17093\ : std_logic;
signal \foc.u_Park_Transform.n782_adj_2109\ : std_logic;
signal \foc.u_Park_Transform.n779_adj_2070_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n17094\ : std_logic;
signal \foc.u_Park_Transform.n786_adj_2152\ : std_logic;
signal \foc.u_Park_Transform.n783_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n17095\ : std_logic;
signal \foc.u_Park_Transform.n790\ : std_logic;
signal \foc.u_Park_Transform.n787_adj_2149_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n17096\ : std_logic;
signal \foc.u_Park_Transform.n17097\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n66\ : std_logic;
signal \foc.u_Park_Transform.n17191\ : std_logic;
signal \foc.u_Park_Transform.n115\ : std_logic;
signal \foc.u_Park_Transform.n17192\ : std_logic;
signal \foc.u_Park_Transform.n164\ : std_logic;
signal \foc.u_Park_Transform.n17193\ : std_logic;
signal \foc.u_Park_Transform.n213\ : std_logic;
signal \foc.u_Park_Transform.n17194\ : std_logic;
signal \foc.u_Park_Transform.n262_adj_1996\ : std_logic;
signal \foc.u_Park_Transform.n17195\ : std_logic;
signal \foc.u_Park_Transform.n311\ : std_logic;
signal \foc.u_Park_Transform.n17196\ : std_logic;
signal \foc.u_Park_Transform.n360\ : std_logic;
signal \foc.u_Park_Transform.n17197\ : std_logic;
signal \foc.u_Park_Transform.n17198\ : std_logic;
signal \foc.u_Park_Transform.n409\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n458\ : std_logic;
signal \foc.u_Park_Transform.n17199\ : std_logic;
signal \foc.u_Park_Transform.n507_adj_2165\ : std_logic;
signal \foc.u_Park_Transform.n17200\ : std_logic;
signal \foc.u_Park_Transform.n556_adj_2164\ : std_logic;
signal \foc.u_Park_Transform.n17201\ : std_logic;
signal \foc.u_Park_Transform.n605_adj_2163\ : std_logic;
signal \foc.u_Park_Transform.n17202\ : std_logic;
signal \foc.u_Park_Transform.n654_adj_2162\ : std_logic;
signal \foc.u_Park_Transform.n17203\ : std_logic;
signal \foc.u_Park_Transform.n703_adj_2160\ : std_logic;
signal \foc.u_Park_Transform.n754_adj_2159\ : std_logic;
signal \foc.u_Park_Transform.n17204\ : std_logic;
signal \foc.u_Park_Transform.n755_adj_2161\ : std_logic;
signal \foc.u_Park_Transform.n755_adj_2161_THRU_CO\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \foc.u_Park_Transform.n16993\ : std_logic;
signal \foc.u_Park_Transform.n16994\ : std_logic;
signal \foc.u_Park_Transform.n16995\ : std_logic;
signal \foc.u_Park_Transform.n16996\ : std_logic;
signal \foc.u_Park_Transform.n16997\ : std_logic;
signal \foc.u_Park_Transform.n16998\ : std_logic;
signal \foc.u_Park_Transform.n16999\ : std_logic;
signal \foc.u_Park_Transform.n17000\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \foc.u_Park_Transform.n17001\ : std_logic;
signal \foc.u_Park_Transform.n17002\ : std_logic;
signal \foc.u_Park_Transform.n17003\ : std_logic;
signal \foc.u_Park_Transform.n17004\ : std_logic;
signal \foc.u_Park_Transform.n17005\ : std_logic;
signal \foc.u_Park_Transform.n757\ : std_logic;
signal \foc.u_Park_Transform.n758\ : std_logic;
signal \foc.u_Park_Transform.n17006\ : std_logic;
signal \foc.u_Park_Transform.n759\ : std_logic;
signal \foc.u_Park_Transform.n759_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n610\ : std_logic;
signal \foc.u_Park_Transform.n69_adj_2059\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n72_adj_2062\ : std_logic;
signal \foc.u_Park_Transform.n118_adj_2037\ : std_logic;
signal \foc.u_Park_Transform.n16978\ : std_logic;
signal \foc.u_Park_Transform.n121_adj_2051\ : std_logic;
signal \foc.u_Park_Transform.n167_adj_2029\ : std_logic;
signal \foc.u_Park_Transform.n16979\ : std_logic;
signal \foc.u_Park_Transform.n170_adj_2048\ : std_logic;
signal \foc.u_Park_Transform.n216_adj_2025\ : std_logic;
signal \foc.u_Park_Transform.n16980\ : std_logic;
signal \foc.u_Park_Transform.n219_adj_2040\ : std_logic;
signal \foc.u_Park_Transform.n265_adj_2023\ : std_logic;
signal \foc.u_Park_Transform.n16981\ : std_logic;
signal \foc.u_Park_Transform.n268_adj_2027\ : std_logic;
signal \foc.u_Park_Transform.n314_adj_2010\ : std_logic;
signal \foc.u_Park_Transform.n16982\ : std_logic;
signal \foc.u_Park_Transform.n317_adj_2021\ : std_logic;
signal \foc.u_Park_Transform.n363_adj_1998\ : std_logic;
signal \foc.u_Park_Transform.n16983\ : std_logic;
signal \foc.u_Park_Transform.n366_adj_2013\ : std_logic;
signal \foc.u_Park_Transform.n412_adj_1995\ : std_logic;
signal \foc.u_Park_Transform.n16984\ : std_logic;
signal \foc.u_Park_Transform.n16985\ : std_logic;
signal \foc.u_Park_Transform.n415\ : std_logic;
signal \foc.u_Park_Transform.n461_adj_2007\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n464\ : std_logic;
signal \foc.u_Park_Transform.n510\ : std_logic;
signal \foc.u_Park_Transform.n16986\ : std_logic;
signal \foc.u_Park_Transform.n513\ : std_logic;
signal \foc.u_Park_Transform.n559\ : std_logic;
signal \foc.u_Park_Transform.n16987\ : std_logic;
signal \foc.u_Park_Transform.n562\ : std_logic;
signal \foc.u_Park_Transform.n608_adj_2067\ : std_logic;
signal \foc.u_Park_Transform.n16988\ : std_logic;
signal \foc.u_Park_Transform.n611_adj_2107\ : std_logic;
signal \foc.u_Park_Transform.n657_adj_2064\ : std_logic;
signal \foc.u_Park_Transform.n16989\ : std_logic;
signal \foc.u_Park_Transform.n660_adj_2091\ : std_logic;
signal \foc.u_Park_Transform.n607\ : std_logic;
signal \foc.u_Park_Transform.n706_adj_2044\ : std_logic;
signal \foc.u_Park_Transform.n16990\ : std_logic;
signal \foc.u_Park_Transform.n761\ : std_logic;
signal \foc.u_Park_Transform.n709_adj_2066\ : std_logic;
signal \foc.u_Park_Transform.n762_adj_2065\ : std_logic;
signal \foc.u_Park_Transform.n16991\ : std_logic;
signal \foc.u_Park_Transform.n763_adj_2054\ : std_logic;
signal \foc.u_Park_Transform.n763_adj_2054_THRU_CO\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2411\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2414\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2511\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2514\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2611\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2614\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2711\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2714\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2811\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2814\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2911\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2914\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3011\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3014\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3111\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17374\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3114\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3215\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216\ : std_logic;
signal \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_CO\ : std_logic;
signal \foc.Look_Up_Table_out1_1_0\ : std_logic;
signal n794 : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n81_adj_750\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n130_adj_748\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17856\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n179_adj_746\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17857\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n228_adj_742\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17858\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n277_adj_741\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17859\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n326\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17860\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n375\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17861\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n424\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17862\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17863\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n473\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n522\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17864\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17865\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17957\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17958\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17959\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17960\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17961\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17962\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17963\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17964\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n770_adj_597\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17965\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n774\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17966\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n778_adj_737\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17967\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17968\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17969\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17970\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17971\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17972\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n75_adj_618\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18092\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n124_adj_616\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18093\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n173_adj_614\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18094\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n222_adj_612\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18095\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n271_adj_610\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18096\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n320_adj_608\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18097\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n369_adj_606\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18098\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18099\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n418_adj_605\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n467_adj_604\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18100\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n516_adj_603\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18101\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n565_adj_602\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18102\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n614_adj_601\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18103\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n663_adj_600\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18104\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n712_adj_599\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n766_adj_619\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18105\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_CO\ : std_logic;
signal \foc.dCurrent_4\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \foc.dCurrent_5\ : std_logic;
signal \foc.u_Park_Transform.n17277\ : std_logic;
signal \foc.dCurrent_6\ : std_logic;
signal \foc.u_Park_Transform.n17278\ : std_logic;
signal \foc.dCurrent_7\ : std_logic;
signal \foc.u_Park_Transform.n17279\ : std_logic;
signal \foc.dCurrent_8\ : std_logic;
signal \foc.u_Park_Transform.n17280\ : std_logic;
signal \foc.dCurrent_9\ : std_logic;
signal \foc.u_Park_Transform.n17281\ : std_logic;
signal \foc.dCurrent_10\ : std_logic;
signal \foc.u_Park_Transform.n17282\ : std_logic;
signal \foc.dCurrent_11\ : std_logic;
signal \foc.u_Park_Transform.n17283\ : std_logic;
signal \foc.u_Park_Transform.n17284\ : std_logic;
signal \foc.dCurrent_12\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \foc.dCurrent_13\ : std_logic;
signal \foc.u_Park_Transform.n17285\ : std_logic;
signal \foc.dCurrent_14\ : std_logic;
signal \foc.u_Park_Transform.n17286\ : std_logic;
signal \foc.dCurrent_15\ : std_logic;
signal \foc.u_Park_Transform.n17287\ : std_logic;
signal \foc.dCurrent_16\ : std_logic;
signal \foc.u_Park_Transform.n17288\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_15\ : std_logic;
signal \foc.dCurrent_17\ : std_logic;
signal \foc.u_Park_Transform.n17289\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_16\ : std_logic;
signal \foc.dCurrent_18\ : std_logic;
signal \foc.u_Park_Transform.n17290\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_17\ : std_logic;
signal \foc.dCurrent_19\ : std_logic;
signal \foc.u_Park_Transform.n17291\ : std_logic;
signal \foc.u_Park_Transform.n17292\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_18\ : std_logic;
signal \foc.dCurrent_20\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_19\ : std_logic;
signal \foc.dCurrent_21\ : std_logic;
signal \foc.u_Park_Transform.n17293\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_20\ : std_logic;
signal \foc.dCurrent_22\ : std_logic;
signal \foc.u_Park_Transform.n17294\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_21\ : std_logic;
signal \foc.dCurrent_23\ : std_logic;
signal \foc.u_Park_Transform.n17295\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_22\ : std_logic;
signal \foc.dCurrent_24\ : std_logic;
signal \foc.u_Park_Transform.n17296\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_23\ : std_logic;
signal \foc.dCurrent_25\ : std_logic;
signal \foc.u_Park_Transform.n17297\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_24\ : std_logic;
signal \foc.u_Park_Transform.n17298\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_25\ : std_logic;
signal \foc.u_Park_Transform.n17299\ : std_logic;
signal \foc.u_Park_Transform.n17300\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_26\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_27\ : std_logic;
signal \foc.u_Park_Transform.n17301\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_28\ : std_logic;
signal \foc.u_Park_Transform.n17302\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_29\ : std_logic;
signal \foc.u_Park_Transform.n17303\ : std_logic;
signal \foc.dCurrent_31_cascade_\ : std_logic;
signal \foc.dCurrent_29\ : std_logic;
signal \foc.dCurrent_28\ : std_logic;
signal \foc.dCurrent_30\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n17221\ : std_logic;
signal \foc.u_Park_Transform.n17222\ : std_logic;
signal \foc.u_Park_Transform.n17223\ : std_logic;
signal \foc.u_Park_Transform.n17224\ : std_logic;
signal \foc.u_Park_Transform.n17225\ : std_logic;
signal \foc.u_Park_Transform.n17226\ : std_logic;
signal \foc.u_Park_Transform.n17227\ : std_logic;
signal \foc.u_Park_Transform.n17228\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n17229\ : std_logic;
signal \foc.u_Park_Transform.n17230\ : std_logic;
signal \foc.u_Park_Transform.n17231\ : std_logic;
signal \foc.u_Park_Transform.n17232\ : std_logic;
signal \foc.u_Park_Transform.n17233\ : std_logic;
signal \foc.u_Park_Transform.n746\ : std_logic;
signal \foc.u_Park_Transform.n17234\ : std_logic;
signal \foc.u_Park_Transform.n747\ : std_logic;
signal \foc.u_Park_Transform.n747_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n604\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \foc.u_Park_Transform.n66_adj_2033\ : std_logic;
signal \foc.u_Park_Transform.n17008\ : std_logic;
signal \foc.u_Park_Transform.n115_adj_2028\ : std_logic;
signal \foc.u_Park_Transform.n17009\ : std_logic;
signal \foc.u_Park_Transform.n164_adj_2014\ : std_logic;
signal \foc.u_Park_Transform.n17010\ : std_logic;
signal \foc.u_Park_Transform.n213_adj_1999\ : std_logic;
signal \foc.u_Park_Transform.n17011\ : std_logic;
signal \foc.u_Park_Transform.n262\ : std_logic;
signal \foc.u_Park_Transform.n17012\ : std_logic;
signal \foc.u_Park_Transform.n311_adj_2022\ : std_logic;
signal \foc.u_Park_Transform.n17013\ : std_logic;
signal \foc.u_Park_Transform.n360_adj_2009\ : std_logic;
signal \foc.u_Park_Transform.n17014\ : std_logic;
signal \foc.u_Park_Transform.n17015\ : std_logic;
signal \foc.u_Park_Transform.n409_adj_1997\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \foc.u_Park_Transform.n458_adj_2093\ : std_logic;
signal \foc.u_Park_Transform.n17016\ : std_logic;
signal \foc.u_Park_Transform.n507\ : std_logic;
signal \foc.u_Park_Transform.n17017\ : std_logic;
signal \foc.u_Park_Transform.n556\ : std_logic;
signal \foc.u_Park_Transform.n17018\ : std_logic;
signal \foc.u_Park_Transform.n605\ : std_logic;
signal \foc.u_Park_Transform.n17019\ : std_logic;
signal \foc.u_Park_Transform.n654\ : std_logic;
signal \foc.u_Park_Transform.n17020\ : std_logic;
signal \foc.u_Park_Transform.n753\ : std_logic;
signal \foc.u_Park_Transform.n703\ : std_logic;
signal \foc.u_Park_Transform.n754\ : std_logic;
signal \foc.u_Park_Transform.n17021\ : std_logic;
signal \foc.u_Park_Transform.n755\ : std_logic;
signal \foc.u_Park_Transform.n755_THRU_CO\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n17068\ : std_logic;
signal \foc.u_Park_Transform.n17069\ : std_logic;
signal \foc.u_Park_Transform.n17070\ : std_logic;
signal \foc.u_Park_Transform.n17071\ : std_logic;
signal \foc.u_Park_Transform.n17072\ : std_logic;
signal \foc.u_Park_Transform.n17073\ : std_logic;
signal \foc.u_Park_Transform.n17074\ : std_logic;
signal \foc.u_Park_Transform.n17075\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n17076\ : std_logic;
signal \foc.u_Park_Transform.n17077\ : std_logic;
signal \foc.u_Park_Transform.n17078\ : std_logic;
signal \foc.u_Park_Transform.n17079\ : std_logic;
signal \foc.u_Park_Transform.n17080\ : std_logic;
signal \foc.u_Park_Transform.n738_adj_2003\ : std_logic;
signal \foc.u_Park_Transform.n17081\ : std_logic;
signal \foc.u_Park_Transform.n739_adj_2006\ : std_logic;
signal \foc.u_Park_Transform.n739_adj_2006_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_2\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_3\ : std_logic;
signal \foc.u_Park_Transform.n15748\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_4\ : std_logic;
signal \foc.u_Park_Transform.n15749\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_5\ : std_logic;
signal \foc.u_Park_Transform.n15750\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_6\ : std_logic;
signal \foc.u_Park_Transform.n15751\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_7\ : std_logic;
signal \foc.u_Park_Transform.n15752\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_8\ : std_logic;
signal \foc.u_Park_Transform.n15753\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_9\ : std_logic;
signal \foc.u_Park_Transform.n15754\ : std_logic;
signal \foc.u_Park_Transform.n15755\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_10\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_11\ : std_logic;
signal \foc.u_Park_Transform.n15756\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_12\ : std_logic;
signal \foc.u_Park_Transform.n15757\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_13\ : std_logic;
signal \foc.u_Park_Transform.n15758\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_14\ : std_logic;
signal \foc.u_Park_Transform.n15759\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_15\ : std_logic;
signal \foc.u_Park_Transform.n15760\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_16\ : std_logic;
signal \foc.u_Park_Transform.n15761\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_17\ : std_logic;
signal \foc.u_Park_Transform.n15762\ : std_logic;
signal \foc.u_Park_Transform.n15763\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_18\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_19\ : std_logic;
signal \foc.u_Park_Transform.n15764\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_20\ : std_logic;
signal \foc.u_Park_Transform.n15765\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_21\ : std_logic;
signal \foc.u_Park_Transform.n15766\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_22\ : std_logic;
signal \foc.u_Park_Transform.n15767\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_23\ : std_logic;
signal \foc.u_Park_Transform.n15768\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_24\ : std_logic;
signal \foc.u_Park_Transform.n15769\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_25\ : std_logic;
signal \foc.u_Park_Transform.n15770\ : std_logic;
signal \foc.u_Park_Transform.n15771\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_26\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_27\ : std_logic;
signal \foc.u_Park_Transform.n15772\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_28\ : std_logic;
signal \foc.u_Park_Transform.n15773\ : std_logic;
signal \foc.u_Park_Transform.Product4_mul_temp_29\ : std_logic;
signal \foc.u_Park_Transform.n15774\ : std_logic;
signal \foc.qCurrent_21\ : std_logic;
signal \foc.qCurrent_29\ : std_logic;
signal \foc.qCurrent_23\ : std_logic;
signal \foc.qCurrent_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n84_adj_749\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n133_adj_747\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17727\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n182_adj_745\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17728\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n231_adj_744\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17729\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n280_adj_743\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17730\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n329_adj_740\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17731\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n378_adj_739\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17732\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17733\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17734\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n782_adj_735\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_CO\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18047\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18048\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18049\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18050\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18051\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18052\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18053\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18054\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18055\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18056\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18057\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18058\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18059\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n754_adj_667\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18060\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_CO\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n63_adj_682\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18032\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n112_adj_681\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18033\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n161_adj_680\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18034\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n210_adj_679\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18035\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n259_adj_678\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18036\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n308_adj_677\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18037\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n357_adj_676\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18038\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18039\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n406_adj_675\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n455_adj_674\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18040\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n504_adj_673\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18041\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n553_adj_672\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18042\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n602_adj_671\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18043\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n651_adj_670\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18044\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n700_adj_669\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n750_adj_683\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18045\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_CO\ : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15775\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15776\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15777\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15778\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15779\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15780\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15781\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15782\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n24\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15783\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15784\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15785\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15786\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15787\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15788\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15789\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15790\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n16\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15_adj_518\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15791\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n14_adj_517\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15792\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15793\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n12_adj_516\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15794\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15795\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15796\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15797\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15798\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n8\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15799\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15800\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15801\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n4_adj_515\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15802\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15803\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15804\ : std_logic;
signal \foc.dCurrent_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n7\ : std_logic;
signal \foc.dCurrent_3\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_2\ : std_logic;
signal \foc.u_Park_Transform.n17251\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_3\ : std_logic;
signal \foc.u_Park_Transform.n17252\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_4\ : std_logic;
signal \foc.u_Park_Transform.n17253\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_5\ : std_logic;
signal \foc.u_Park_Transform.n17254\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_6\ : std_logic;
signal \foc.u_Park_Transform.n17255\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_7\ : std_logic;
signal \foc.u_Park_Transform.n17256\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_8\ : std_logic;
signal \foc.u_Park_Transform.n17257\ : std_logic;
signal \foc.u_Park_Transform.n17258\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_9\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_10\ : std_logic;
signal \foc.u_Park_Transform.n17259\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_11\ : std_logic;
signal \foc.u_Park_Transform.n17260\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_12\ : std_logic;
signal \foc.u_Park_Transform.n17261\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_13\ : std_logic;
signal \foc.u_Park_Transform.n17262\ : std_logic;
signal \foc.u_Park_Transform.dCurrent_2\ : std_logic;
signal \foc.u_Park_Transform.Product1_mul_temp_14\ : std_logic;
signal \foc.u_Park_Transform.n17263\ : std_logic;
signal \foc.u_Park_Transform.n737\ : std_logic;
signal \foc.u_Park_Transform.n738\ : std_logic;
signal \foc.u_Park_Transform.n17264\ : std_logic;
signal \foc.u_Park_Transform.n739\ : std_logic;
signal \foc.u_Park_Transform.n739_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n54_adj_2095\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n57_adj_2116\ : std_logic;
signal \foc.u_Park_Transform.n103_adj_2092\ : std_logic;
signal \foc.u_Park_Transform.n17236\ : std_logic;
signal \foc.u_Park_Transform.n106_adj_2115\ : std_logic;
signal \foc.u_Park_Transform.n152_adj_2088\ : std_logic;
signal \foc.u_Park_Transform.n17237\ : std_logic;
signal \foc.u_Park_Transform.n155_adj_2114\ : std_logic;
signal \foc.u_Park_Transform.n201_adj_2085\ : std_logic;
signal \foc.u_Park_Transform.n17238\ : std_logic;
signal \foc.u_Park_Transform.n204_adj_2113\ : std_logic;
signal \foc.u_Park_Transform.n250_adj_2084\ : std_logic;
signal \foc.u_Park_Transform.n17239\ : std_logic;
signal \foc.u_Park_Transform.n253_adj_2112\ : std_logic;
signal \foc.u_Park_Transform.n299_adj_2083\ : std_logic;
signal \foc.u_Park_Transform.n17240\ : std_logic;
signal \foc.u_Park_Transform.n302_adj_2111\ : std_logic;
signal \foc.u_Park_Transform.n348_adj_2082\ : std_logic;
signal \foc.u_Park_Transform.n17241\ : std_logic;
signal \foc.u_Park_Transform.n351_adj_2108\ : std_logic;
signal \foc.u_Park_Transform.n397_adj_2081\ : std_logic;
signal \foc.u_Park_Transform.n17242\ : std_logic;
signal \foc.u_Park_Transform.n17243\ : std_logic;
signal \foc.u_Park_Transform.n400_adj_2106\ : std_logic;
signal \foc.u_Park_Transform.n446_adj_2079\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n449_adj_2103\ : std_logic;
signal \foc.u_Park_Transform.n495_adj_2077\ : std_logic;
signal \foc.u_Park_Transform.n17244\ : std_logic;
signal \foc.u_Park_Transform.n498_adj_2102\ : std_logic;
signal \foc.u_Park_Transform.n544_adj_2074\ : std_logic;
signal \foc.u_Park_Transform.n17245\ : std_logic;
signal \foc.u_Park_Transform.n547_adj_2100\ : std_logic;
signal \foc.u_Park_Transform.n593_adj_2073\ : std_logic;
signal \foc.u_Park_Transform.n17246\ : std_logic;
signal \foc.u_Park_Transform.n596_adj_2099\ : std_logic;
signal \foc.u_Park_Transform.n642_adj_2072\ : std_logic;
signal \foc.u_Park_Transform.n17247\ : std_logic;
signal \foc.u_Park_Transform.n645_adj_2098\ : std_logic;
signal \foc.u_Park_Transform.n691_adj_2071\ : std_logic;
signal \foc.u_Park_Transform.n17248\ : std_logic;
signal \foc.u_Park_Transform.n694_adj_2097\ : std_logic;
signal \foc.u_Park_Transform.n742\ : std_logic;
signal \foc.u_Park_Transform.n17249\ : std_logic;
signal \foc.u_Park_Transform.n743\ : std_logic;
signal \foc.u_Park_Transform.n743_THRU_CO\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \foc.u_Park_Transform.n63\ : std_logic;
signal \foc.u_Park_Transform.n17023\ : std_logic;
signal \foc.u_Park_Transform.n112\ : std_logic;
signal \foc.u_Park_Transform.n17024\ : std_logic;
signal \foc.u_Park_Transform.n161\ : std_logic;
signal \foc.u_Park_Transform.n17025\ : std_logic;
signal \foc.u_Park_Transform.n210\ : std_logic;
signal \foc.u_Park_Transform.n17026\ : std_logic;
signal \foc.u_Park_Transform.n259\ : std_logic;
signal \foc.u_Park_Transform.n17027\ : std_logic;
signal \foc.u_Park_Transform.n308\ : std_logic;
signal \foc.u_Park_Transform.n17028\ : std_logic;
signal \foc.u_Park_Transform.n357\ : std_logic;
signal \foc.u_Park_Transform.n17029\ : std_logic;
signal \foc.u_Park_Transform.n17030\ : std_logic;
signal \foc.u_Park_Transform.n406\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \foc.u_Park_Transform.n455\ : std_logic;
signal \foc.u_Park_Transform.n17031\ : std_logic;
signal \foc.u_Park_Transform.n504\ : std_logic;
signal \foc.u_Park_Transform.n17032\ : std_logic;
signal \foc.u_Park_Transform.n553\ : std_logic;
signal \foc.u_Park_Transform.n17033\ : std_logic;
signal \foc.u_Park_Transform.n602\ : std_logic;
signal \foc.u_Park_Transform.n17034\ : std_logic;
signal \foc.u_Park_Transform.n651\ : std_logic;
signal \foc.u_Park_Transform.n17035\ : std_logic;
signal \foc.u_Park_Transform.n700\ : std_logic;
signal \foc.u_Park_Transform.n750_adj_2117\ : std_logic;
signal \foc.u_Park_Transform.n17036\ : std_logic;
signal \foc.u_Park_Transform.n751\ : std_logic;
signal \foc.u_Park_Transform.n751_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n54\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \foc.u_Park_Transform.n103\ : std_logic;
signal \foc.u_Park_Transform.n17053\ : std_logic;
signal \foc.u_Park_Transform.n152\ : std_logic;
signal \foc.u_Park_Transform.n17054\ : std_logic;
signal \foc.u_Park_Transform.n201\ : std_logic;
signal \foc.u_Park_Transform.n17055\ : std_logic;
signal \foc.u_Park_Transform.n250\ : std_logic;
signal \foc.u_Park_Transform.n17056\ : std_logic;
signal \foc.u_Park_Transform.n299\ : std_logic;
signal \foc.u_Park_Transform.n17057\ : std_logic;
signal \foc.u_Park_Transform.n348\ : std_logic;
signal \foc.u_Park_Transform.n17058\ : std_logic;
signal \foc.u_Park_Transform.n397\ : std_logic;
signal \foc.u_Park_Transform.n17059\ : std_logic;
signal \foc.u_Park_Transform.n17060\ : std_logic;
signal \foc.u_Park_Transform.n446\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \foc.u_Park_Transform.n495\ : std_logic;
signal \foc.u_Park_Transform.n17061\ : std_logic;
signal \foc.u_Park_Transform.n544\ : std_logic;
signal \foc.u_Park_Transform.n17062\ : std_logic;
signal \foc.u_Park_Transform.n593\ : std_logic;
signal \foc.u_Park_Transform.n17063\ : std_logic;
signal \foc.u_Park_Transform.n642\ : std_logic;
signal \foc.u_Park_Transform.n17064\ : std_logic;
signal \foc.u_Park_Transform.n691\ : std_logic;
signal \foc.u_Park_Transform.n17065\ : std_logic;
signal \foc.u_Park_Transform.n742_adj_2086\ : std_logic;
signal \foc.u_Park_Transform.n17066\ : std_logic;
signal \foc.u_Park_Transform.n743_adj_2096\ : std_logic;
signal \foc.u_Park_Transform.n743_adj_2096_THRU_CO\ : std_logic;
signal \foc.qCurrent_6\ : std_logic;
signal \foc.u_Park_Transform.n741\ : std_logic;
signal \Look_Up_Table_out1_1_14\ : std_logic;
signal \Look_Up_Table_out1_1_15\ : std_logic;
signal \foc.qCurrent_8\ : std_logic;
signal \foc.Look_Up_Table_out1_1_1\ : std_logic;
signal \foc.u_Park_Transform.n592\ : std_logic;
signal \foc.qCurrent_3\ : std_logic;
signal \foc.qCurrent_18\ : std_logic;
signal \foc.qCurrent_19\ : std_logic;
signal \foc.qCurrent_13\ : std_logic;
signal \foc.qCurrent_16\ : std_logic;
signal \foc.qCurrent_14\ : std_logic;
signal \foc.qCurrent_4\ : std_logic;
signal \foc.qCurrent_11\ : std_logic;
signal \foc.qCurrent_15\ : std_logic;
signal \foc.qCurrent_22\ : std_logic;
signal \foc.qCurrent_17\ : std_logic;
signal \foc.qCurrent_24\ : std_logic;
signal \foc.qCurrent_27\ : std_logic;
signal \foc.qCurrent_26\ : std_logic;
signal \foc.qCurrent_12\ : std_logic;
signal \foc.qCurrent_28\ : std_logic;
signal \foc.qCurrent_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_757_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_758\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19841_cascade_\ : std_logic;
signal \foc.qCurrent_31\ : std_logic;
signal \foc.qCurrent_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n87_adj_730\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n136_adj_728\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17973\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n185_adj_726\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17974\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n234_adj_724\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17975\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n283_adj_723\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17976\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17977\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n786_adj_719\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17978\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n90_adj_729\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n7_adj_760_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_adj_732\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n26_adj_759\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n790_adj_733\ : std_logic;
signal n794_adj_2425 : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n66_adj_666\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n115_adj_665\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18062\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n164_adj_664\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18063\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n213_adj_663\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18064\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n262_adj_662\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18065\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n311_adj_661\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18066\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n360_adj_660\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18067\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n409_adj_659\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18068\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18069\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n458_adj_658\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n507_adj_657\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18070\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n556_adj_656\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18071\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n605_adj_655\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18072\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n654_adj_654\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18073\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n703_adj_653\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18074\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n758_adj_651\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18075\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n69_adj_650\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n72_adj_634\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n118_adj_649\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18077\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n121_adj_633\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n167_adj_648\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18078\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n170_adj_632\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n216_adj_647\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18079\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n219_adj_631\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n265_adj_646\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18080\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n268_adj_630\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n314_adj_645\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18081\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n317_adj_629\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n363_adj_644\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18082\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n366_adj_628\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n412_adj_643\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18083\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18084\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n415_adj_627\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n461_adj_642\ : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n464_adj_626\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n510_adj_641\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18085\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n513_adj_625\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n559_adj_640\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18086\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n562_adj_624\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n608_adj_639\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18087\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n611_adj_623\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n657_adj_638\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18088\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n660_adj_622\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n706_adj_637\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18089\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n709_adj_621\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n762_adj_635\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18090\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_24\ : std_logic;
signal \foc.dCurrent_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n6\ : std_logic;
signal \foc.u_Park_Transform.n601\ : std_logic;
signal \foc.u_Park_Transform.n60_adj_2140\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \foc.u_Park_Transform.n63_adj_2158\ : std_logic;
signal \foc.u_Park_Transform.n109_adj_2139\ : std_logic;
signal \foc.u_Park_Transform.n17206\ : std_logic;
signal \foc.u_Park_Transform.n112_adj_2157\ : std_logic;
signal \foc.u_Park_Transform.n158_adj_2137\ : std_logic;
signal \foc.u_Park_Transform.n17207\ : std_logic;
signal \foc.u_Park_Transform.n161_adj_2156\ : std_logic;
signal \foc.u_Park_Transform.n207_adj_2136\ : std_logic;
signal \foc.u_Park_Transform.n17208\ : std_logic;
signal \foc.u_Park_Transform.n210_adj_2155\ : std_logic;
signal \foc.u_Park_Transform.n256_adj_2135\ : std_logic;
signal \foc.u_Park_Transform.n17209\ : std_logic;
signal \foc.u_Park_Transform.n259_adj_2154\ : std_logic;
signal \foc.u_Park_Transform.n305_adj_2134\ : std_logic;
signal \foc.u_Park_Transform.n17210\ : std_logic;
signal \foc.u_Park_Transform.n308_adj_2153\ : std_logic;
signal \foc.u_Park_Transform.n354_adj_2133\ : std_logic;
signal \foc.u_Park_Transform.n17211\ : std_logic;
signal \foc.u_Park_Transform.n357_adj_2151\ : std_logic;
signal \foc.u_Park_Transform.n403_adj_2132\ : std_logic;
signal \foc.u_Park_Transform.n17212\ : std_logic;
signal \foc.u_Park_Transform.n17213\ : std_logic;
signal \foc.u_Park_Transform.n406_adj_2150\ : std_logic;
signal \foc.u_Park_Transform.n452_adj_2131\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \foc.u_Park_Transform.n455_adj_2148\ : std_logic;
signal \foc.u_Park_Transform.n501_adj_2130\ : std_logic;
signal \foc.u_Park_Transform.n17214\ : std_logic;
signal \foc.u_Park_Transform.n504_adj_2147\ : std_logic;
signal \foc.u_Park_Transform.n550_adj_2129\ : std_logic;
signal \foc.u_Park_Transform.n17215\ : std_logic;
signal \foc.u_Park_Transform.n553_adj_2146\ : std_logic;
signal \foc.u_Park_Transform.n599_adj_2128\ : std_logic;
signal \foc.u_Park_Transform.n17216\ : std_logic;
signal \foc.u_Park_Transform.n602_adj_2144\ : std_logic;
signal \foc.u_Park_Transform.n648_adj_2124\ : std_logic;
signal \foc.u_Park_Transform.n17217\ : std_logic;
signal \foc.u_Park_Transform.n651_adj_2143\ : std_logic;
signal \foc.u_Park_Transform.n697_adj_2121\ : std_logic;
signal \foc.u_Park_Transform.n17218\ : std_logic;
signal \foc.u_Park_Transform.n749\ : std_logic;
signal \foc.u_Park_Transform.n700_adj_2141\ : std_logic;
signal \foc.u_Park_Transform.n750\ : std_logic;
signal \foc.u_Park_Transform.n17219\ : std_logic;
signal \foc.u_Park_Transform.n751_adj_2142\ : std_logic;
signal \foc.u_Park_Transform.n751_adj_2142_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n598\ : std_logic;
signal \foc.u_Park_Transform.n57\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \foc.u_Park_Transform.n60\ : std_logic;
signal \foc.u_Park_Transform.n106\ : std_logic;
signal \foc.u_Park_Transform.n17038\ : std_logic;
signal \foc.u_Park_Transform.n109\ : std_logic;
signal \foc.u_Park_Transform.n155\ : std_logic;
signal \foc.u_Park_Transform.n17039\ : std_logic;
signal \foc.u_Park_Transform.n158\ : std_logic;
signal \foc.u_Park_Transform.n204\ : std_logic;
signal \foc.u_Park_Transform.n17040\ : std_logic;
signal \foc.u_Park_Transform.n207\ : std_logic;
signal \foc.u_Park_Transform.n253\ : std_logic;
signal \foc.u_Park_Transform.n17041\ : std_logic;
signal \foc.u_Park_Transform.n256\ : std_logic;
signal \foc.u_Park_Transform.n302\ : std_logic;
signal \foc.u_Park_Transform.n17042\ : std_logic;
signal \foc.u_Park_Transform.n305\ : std_logic;
signal \foc.u_Park_Transform.n351\ : std_logic;
signal \foc.u_Park_Transform.n17043\ : std_logic;
signal \foc.u_Park_Transform.n354\ : std_logic;
signal \foc.u_Park_Transform.n400\ : std_logic;
signal \foc.u_Park_Transform.n17044\ : std_logic;
signal \foc.u_Park_Transform.n17045\ : std_logic;
signal \foc.u_Park_Transform.n403\ : std_logic;
signal \foc.u_Park_Transform.n449\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \foc.u_Park_Transform.n452\ : std_logic;
signal \foc.u_Park_Transform.n498\ : std_logic;
signal \foc.u_Park_Transform.n17046\ : std_logic;
signal \foc.u_Park_Transform.n501\ : std_logic;
signal \foc.u_Park_Transform.n547\ : std_logic;
signal \foc.u_Park_Transform.n17047\ : std_logic;
signal \foc.u_Park_Transform.n550\ : std_logic;
signal \foc.u_Park_Transform.n596\ : std_logic;
signal \foc.u_Park_Transform.n17048\ : std_logic;
signal \foc.u_Park_Transform.n599\ : std_logic;
signal \foc.u_Park_Transform.n645\ : std_logic;
signal \foc.u_Park_Transform.n17049\ : std_logic;
signal \foc.u_Park_Transform.n648\ : std_logic;
signal \foc.u_Park_Transform.n694\ : std_logic;
signal \foc.u_Park_Transform.n17050\ : std_logic;
signal \foc.u_Park_Transform.n745\ : std_logic;
signal \foc.u_Park_Transform.n697\ : std_logic;
signal \foc.u_Park_Transform.n746_adj_2011\ : std_logic;
signal \foc.u_Park_Transform.n17051\ : std_logic;
signal \foc.u_Park_Transform.n747_adj_2012\ : std_logic;
signal \foc.u_Park_Transform.n747_adj_2012_THRU_CO\ : std_logic;
signal \foc.u_Park_Transform.n6_cascade_\ : std_logic;
signal \foc.Look_Up_Table_out1_1_2\ : std_logic;
signal \foc.u_Park_Transform.n595\ : std_logic;
signal n4 : std_logic;
signal \foc.qCurrent_10\ : std_logic;
signal \foc.qCurrent_7\ : std_logic;
signal \foc.qCurrent_5\ : std_logic;
signal \foc.qCurrent_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n30\ : std_logic;
signal \foc.u_DQ_Current_Control.n31\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15720\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15721\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n27_adj_753\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15722\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15723\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15724\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15725\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15726\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15727\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n22\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_adj_752\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15728\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15729\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15730\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_751\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15731\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15732\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15733\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15734\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15735\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n14\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15736\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15737\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15738\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15739\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15740\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15741\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15742\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15743\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n6\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15744\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n4\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15745\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15746\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15747\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n188_adj_725\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_22\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17987\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17988\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17989\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17990\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17991\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17992\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17993\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17994\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17995\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17996\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17997\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17998\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n17999\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n738_adj_718\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18000\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n739\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_CO\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n60_adj_698\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18017\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n109_adj_697\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18018\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n158_adj_696\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18019\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n207_adj_695\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18020\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n256_adj_694\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18021\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n305_adj_693\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18022\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n354_adj_692\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18023\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18024\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n403_adj_691\ : std_logic;
signal \bfn_16_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n452_adj_690\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18025\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n501_adj_689\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18026\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n550_adj_688\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18027\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n599_adj_687\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18028\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n648_adj_686\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18029\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n697_adj_685\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n746_adj_699\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18030\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n54\ : std_logic;
signal \bfn_16_27_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n57_adj_714\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n103\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18002\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n106_adj_713\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n152\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18003\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n155_adj_712\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n201\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18004\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n204_adj_711\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n250\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18005\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n253_adj_710\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n299\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18006\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n302_adj_709\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n348\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18007\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n351_adj_708\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n397\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18008\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18009\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n400_adj_707\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n446\ : std_logic;
signal \bfn_16_28_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n449_adj_706\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n495\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18010\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n498_adj_705\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n544\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18011\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n547_adj_704\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n593\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18012\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n596_adj_703\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n642\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18013\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n645_adj_702\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n691_adj_717\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18014\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n694_adj_701\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n742_adj_715\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18015\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_CO\ : std_logic;
signal \bfn_17_5_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18135\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18136\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18137\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18138\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18139\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18140\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18141\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18142\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n87_adj_400\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n90\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n136_adj_399\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18167\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n185_adj_398\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18168\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n234_adj_397\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18169\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n283\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18170\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n332\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18171\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18172\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n787\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n188\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n138_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n139\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n237\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n4\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n4_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19269_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19273\ : std_logic;
signal n142_adj_2419 : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19273_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19269\ : std_logic;
signal \foc.u_Park_Transform.n7_cascade_\ : std_logic;
signal \foc.u_Park_Transform.n791\ : std_logic;
signal \foc.u_Park_Transform.n4_cascade_\ : std_logic;
signal \Look_Up_Table_out1_1_13\ : std_logic;
signal \foc.u_Park_Transform.n14\ : std_logic;
signal \n628_cascade_\ : std_logic;
signal \foc.u_Park_Transform.n12\ : std_logic;
signal n142 : std_logic;
signal n628 : std_logic;
signal \foc.u_Park_Transform.n18_cascade_\ : std_logic;
signal \foc.u_Park_Transform.n19845\ : std_logic;
signal \foc.u_Park_Transform.n26\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n66_adj_433\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17781\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17782\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17783\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17784\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17785\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17786\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17787\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17788\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17789\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17790\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17791\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17792\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17793\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17794\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n755\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n63_adj_384\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17766\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n112\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17767\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n161\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17768\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n210\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17769\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n259\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17770\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n308_adj_368\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17771\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n357_adj_366\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17772\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17773\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n406_adj_363\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n455_adj_350\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17774\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n504\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17775\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n553\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17776\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n602\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17777\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n651_adj_474\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17778\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n700_adj_455\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17779\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n751\ : std_logic;
signal \n142_adj_2422_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n14_adj_756\ : std_logic;
signal \Amp25_out1_14\ : std_logic;
signal n142_adj_2422 : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n6_adj_763\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n139_adj_727\ : std_logic;
signal \n141_adj_2421_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19450_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19743\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19741_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20180_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19827_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19812\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18\ : std_logic;
signal \Error_sub_temp_30_adj_2385\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n737\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n741\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18369\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n745\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18370\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n749\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18371\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n753\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18372\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n757\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18373\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n761\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18374\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n765\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18375\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18376\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n769\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n773\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18377\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n777\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18378\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n781\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18379\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n785\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18380\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n789\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18381\ : std_logic;
signal n793_adj_2424 : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18382\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n795\ : std_logic;
signal \bfn_18_5_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n84\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17266\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n133\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17267\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n182\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17268\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n231\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17269\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n280\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17270\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n329\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17271\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n378\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17272\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17273\ : std_logic;
signal \bfn_18_6_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17274\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n427\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17275\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_22\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17942\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17943\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17944\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17945\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17946\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17947\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17948\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17949\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17950\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n777\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17951\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n781\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17952\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n785\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17953\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n789\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17954\ : std_logic;
signal n793 : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17955\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n795\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n84_adj_389\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17882\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17883\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17884\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17885\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17886\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17887\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17888\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17889\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17890\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17891\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17892\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17893\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17894\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17895\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n779\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n81_adj_457\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17867\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n130_adj_453\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17868\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n179_adj_452\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17869\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n228_adj_450\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17870\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n277_adj_448\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17871\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n326_adj_443\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17872\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n375_adj_438\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17873\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17874\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n424_adj_435\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n473_adj_431\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17875\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n522_adj_430\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17876\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n571\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17877\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n620\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17878\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n669\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17879\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n718\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17880\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n775\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n78_adj_480\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17841\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n127_adj_479\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17842\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n176_adj_478\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17843\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n225_adj_477\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17844\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n274_adj_476\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17845\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n323_adj_475\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17846\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n372_adj_473\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17847\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17848\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n421_adj_465\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n470_adj_463\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17849\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n519_adj_461\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17850\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n568_adj_460\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17851\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n617_adj_459\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17852\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n666\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17853\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n715\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17854\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n75\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17826\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n124_adj_507\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17827\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n173_adj_506\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17828\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n222_adj_505\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17829\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n271_adj_503\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17830\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n320_adj_502\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17831\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n369_adj_501\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17832\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17833\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n418_adj_500\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n467_adj_499\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17834\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n516_adj_498\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17835\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n565_adj_497\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17836\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n614_adj_496\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17837\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n663_adj_494\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17838\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n712_adj_493\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17839\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n767\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n60\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17751\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n109_adj_383\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17752\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n158_adj_375\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17753\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n207\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17754\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n256\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17755\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n305\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17756\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n354_adj_367\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17757\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17758\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n403_adj_365\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n452_adj_362\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17759\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n501\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17760\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n550\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17761\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n599\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17762\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n648_adj_347\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17763\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n697\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17764\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n747\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20108\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20092_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19914_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20102\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20086_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19890\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20858_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20174\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_1\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15883\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15884\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15885\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_4\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15886\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15887\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15888\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15889\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15890\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_8\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15891\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15892\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15893\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15894\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15895\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_14\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15896\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15897\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15898\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_16\ : std_logic;
signal \bfn_18_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15899\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15900\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15901\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15902\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15903\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15904\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15905\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15906\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_24\ : std_logic;
signal \bfn_18_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15907\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15908\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15909\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15910\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15911\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15912\ : std_logic;
signal \bfn_18_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n93\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18354\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n142\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18355\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n191\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18356\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n240\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18357\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n289\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18358\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n338\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18359\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n387\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18360\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18361\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n436\ : std_logic;
signal \bfn_18_27_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n485\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18362\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n534\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18363\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n583\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18364\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n632\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18365\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n681\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18366\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n730\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18367\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n791\ : std_logic;
signal \bfn_19_5_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17641\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17642\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17643\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17644\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17645\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17646\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17647\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17648\ : std_logic;
signal \bfn_19_6_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17649\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17650\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17651\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17652\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17653\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n769\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17654\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n771\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n75_adj_510\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17626\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n124\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17627\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n173\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17628\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n222\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17629\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n271\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17630\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n320\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17631\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n369\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17632\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17633\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n418\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n467\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17634\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n516\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17635\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n565\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17636\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n614\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17637\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n663\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17638\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n765\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n712\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17639\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382\ : std_logic;
signal \bfn_19_9_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n93\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17927\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n142_adj_414\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17928\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n191\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17929\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n240\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17930\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n289\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17931\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n338\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17932\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n387\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17933\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17934\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n436\ : std_logic;
signal \bfn_19_10_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n485\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17935\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n534\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17936\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n583\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17937\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n632\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17938\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n681\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17939\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n730\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17940\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416\ : std_logic;
signal \bfn_19_11_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n90_adj_420\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17912\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n139_adj_419\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17913\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n188_adj_418\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17914\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n237_adj_417\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17915\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n286\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17916\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n335\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17917\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n384\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17918\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17919\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n433\ : std_logic;
signal \bfn_19_12_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n482\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17920\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n531\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17921\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n580\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17922\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n629\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17923\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n678\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17924\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n727\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17925\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421\ : std_logic;
signal \bfn_19_13_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n72\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17811\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n121\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17812\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n170\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17813\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n219\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17814\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n268_adj_437\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17815\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n317_adj_428\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17816\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n366_adj_426\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17817\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17818\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n415\ : std_logic;
signal \bfn_19_14_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n464_adj_423\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17819\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n513_adj_412\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17820\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n562_adj_378\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17821\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n611_adj_373\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17822\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n660_adj_372\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17823\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n709\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17824\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n763\ : std_logic;
signal \bfn_19_15_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n69\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n115\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17796\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n118\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n164\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17797\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n167\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n213\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17798\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n216\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n262_adj_425\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17799\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n265\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n311_adj_422\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17800\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n314_adj_401\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n360\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17801\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n363_adj_380\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n409\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17802\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17803\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n412\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n458\ : std_logic;
signal \bfn_19_16_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n461\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n507\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17804\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n510\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n556_adj_370\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17805\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n559_adj_358\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n605_adj_462\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17806\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n608_adj_377\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n654_adj_456\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17807\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n657_adj_360\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n703_adj_359\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17808\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n706_adj_371\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17809\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354\ : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17711\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17712\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n746\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17713\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n750\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17714\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n754\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17715\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n758\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17716\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n762\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17717\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17718\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n766\ : std_logic;
signal \bfn_19_18_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n770\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17719\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n774\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17720\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n778\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17721\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17722\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n786\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17723\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n790_adj_415\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17724\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n794_adj_413\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17725\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17726\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_CO\ : std_logic;
signal \bfn_19_19_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20870\ : std_logic;
signal \foc.preSatVoltage_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n738\ : std_logic;
signal \bfn_19_21_0_\ : std_logic;
signal \Error_sub_temp_31_adj_2384\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18144\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n8356\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18145\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18146\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18147\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18148\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18149\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18150\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18151\ : std_logic;
signal \bfn_19_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18152\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18153\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18154\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18155\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18156\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n790\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18157\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n794\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18158\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18159\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n796\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \bfn_19_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n60\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18189\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18190\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18191\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18192\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18193\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18194\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18195\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18196\ : std_logic;
signal \bfn_19_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18197\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18198\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18199\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18200\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18201\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n746\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18202\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n747\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_CO\ : std_logic;
signal \bfn_19_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n90\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18339\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n139\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18340\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n188\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18341\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n237\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18342\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n286\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18343\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n335\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18344\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n384\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18345\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18346\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n433\ : std_logic;
signal \bfn_19_27_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n482\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18347\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n531\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18348\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n580\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18349\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n629\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18350\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n678\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18351\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n727\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n786\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18352\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n787\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_CO\ : std_logic;
signal \bfn_19_28_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n87\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18324\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n136\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18325\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n185\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18326\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n234\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18327\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n283\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18328\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n332\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18329\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n381\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18330\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18331\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n430\ : std_logic;
signal \bfn_19_29_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n479\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18332\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n528\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18333\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n577\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18334\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n626\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18335\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n675\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18336\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n724\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n782\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18337\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n783\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n78\ : std_logic;
signal \bfn_20_5_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n81\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n127\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18122\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n130\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n176\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18123\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n179\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n225\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18124\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n228\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n274\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18125\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n277\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n323\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18126\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n326\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n372\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18127\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n375\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n421\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18128\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18129\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n424\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n470\ : std_logic;
signal \bfn_20_6_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n473\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n519\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18130\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n568\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18131\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n617\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18132\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n773\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n522\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n18133\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357\ : std_logic;
signal \bfn_20_7_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n72_adj_508\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17611\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n121_adj_504\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17612\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n170_adj_490\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17613\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n219_adj_472\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17614\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n268\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17615\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n317\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17616\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n366\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17617\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17618\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n415_adj_449\ : std_logic;
signal \bfn_20_8_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n464\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17619\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n513\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17620\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n562\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17621\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n611\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17622\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n660\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17623\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n709_adj_512\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n761\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17624\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386\ : std_logic;
signal \bfn_20_9_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17581\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17582\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17583\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17584\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17585\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17586\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17587\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17588\ : std_logic;
signal \bfn_20_10_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17589\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17590\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17591\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17592\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17593\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n753\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17594\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404\ : std_logic;
signal \bfn_20_11_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n87\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n133_adj_388\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17897\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n136\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n182_adj_451\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17898\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n185\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n231_adj_387\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17899\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n234\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n280_adj_379\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17900\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n283_adj_514\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n329_adj_439\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17901\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n332_adj_513\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n378_adj_436\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17902\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n381\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n427_adj_432\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17903\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17904\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n430\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n476\ : std_logic;
signal \bfn_20_12_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n479\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n525\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17905\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n528\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n574\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17906\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n577\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n623\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17907\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n626\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n672\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17908\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n675\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n721\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17909\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n724\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n782\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17910\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n783\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_CO\ : std_logic;
signal \Error_sub_temp_30\ : std_logic;
signal \bfn_20_14_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17505\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17506\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17507\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17508\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n754_adj_405\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17509\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17510\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n762_adj_402\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17511\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17512\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n766_adj_385\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_CO\ : std_logic;
signal \bfn_20_15_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n770_adj_381\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17513\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n774_adj_374\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17514\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n778_adj_356\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17515\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n782_adj_351\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17516\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n786_adj_348\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17517\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n790\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17518\ : std_logic;
signal n794_adj_2420 : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n791\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17519\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17520\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n796\ : std_logic;
signal \bfn_20_16_0_\ : std_logic;
signal \foc.preSatVoltage_19\ : std_logic;
signal \foc.qVoltage_10\ : std_logic;
signal \foc.preSatVoltage_22\ : std_logic;
signal \foc.qVoltage_13\ : std_logic;
signal \foc.qVoltage_3\ : std_logic;
signal \foc.preSatVoltage_13\ : std_logic;
signal \foc.qVoltage_4_cascade_\ : std_logic;
signal \foc.preSatVoltage_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17\ : std_logic;
signal \foc.qVoltage_8_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n8265\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19884\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20586_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20590\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20614\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20602_cascade_\ : std_logic;
signal \foc.qVoltage_7\ : std_logic;
signal \Error_sub_temp_31\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20664_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20650_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n58_cascade_\ : std_logic;
signal \Saturate_out1_31__N_266_adj_2417_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20620\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20608\ : std_logic;
signal \Saturate_out1_31__N_267_adj_2418_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n22_adj_762_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20694_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19729_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20676\ : std_logic;
signal \bfn_20_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n63\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n109\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18204\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n158\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18205\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n207\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18206\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n256\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18207\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n305\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18208\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n354\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18209\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n403\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18210\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18211\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n452\ : std_logic;
signal \bfn_20_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n501\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18212\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n550\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18213\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n599\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18214\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n648\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18215\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n697\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18216\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n750\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18217\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n751\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_CO\ : std_logic;
signal \bfn_20_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n66\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n112\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18219\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n161\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18220\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n210\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18221\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n259\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18222\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n308\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18223\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n357\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18224\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n406\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18225\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18226\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n455\ : std_logic;
signal \bfn_20_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n504\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18227\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n553\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18228\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n602\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18229\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n651\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18230\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n700\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18231\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n754\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18232\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n755\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_CO\ : std_logic;
signal \bfn_20_28_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n84\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18309\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n133\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18310\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n182\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18311\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n231\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18312\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n280\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18313\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n329\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18314\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n378\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18315\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18316\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n427\ : std_logic;
signal \bfn_20_29_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n476\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18317\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n525\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18318\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n574\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18319\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n623\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18320\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n672\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18321\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n721\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n778\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18322\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n779\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n66\ : std_logic;
signal \bfn_21_7_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n69_adj_489\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n115_adj_488\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17596\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n118_adj_487\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n164_adj_466\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17597\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n167_adj_486\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n213_adj_445\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17598\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n216_adj_485\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n262\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17599\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n265_adj_471\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n311\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17600\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n314\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n360_adj_484\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17601\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n363\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n409_adj_483\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17602\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17603\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n412_adj_482\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n458_adj_468\ : std_logic;
signal \bfn_21_8_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n461_adj_470\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n507_adj_447\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17604\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n510_adj_458\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n556\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17605\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n559\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n605\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17606\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n608\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n654\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17607\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n657\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n703\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17608\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n757\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n706\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n758_adj_403\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17609\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n759\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_CO\ : std_logic;
signal \bfn_21_9_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n63\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17566\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n112_adj_442\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17567\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n161_adj_395\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17568\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n210_adj_393\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17569\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n259_adj_391\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17570\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n308\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17571\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n357\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17572\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17573\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n406\ : std_logic;
signal \bfn_21_10_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n455\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17574\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n504_adj_467\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17575\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n553_adj_446\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17576\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n602_adj_355\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17577\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n651\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17578\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n749\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n700\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n750_adj_407\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17579\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_CO\ : std_logic;
signal \bfn_21_11_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n60_adj_495\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17551\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n109\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17552\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n158\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17553\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n207_adj_394\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17554\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n256_adj_392\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17555\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n305_adj_390\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17556\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n354\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17557\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17558\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n403\ : std_logic;
signal \bfn_21_12_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n452\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17559\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n501_adj_481\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17560\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n550_adj_441\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17561\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n599_adj_376\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17562\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n648\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17563\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n745\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n697_adj_444\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n746_adj_409\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17564\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_CO\ : std_logic;
signal \foc.dVoltage_2_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20548_cascade_\ : std_logic;
signal \foc.dVoltage_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20562_cascade_\ : std_logic;
signal \foc.dVoltage_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20574_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19727_cascade_\ : std_logic;
signal \foc.qVoltage_5_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20596_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20604\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20588\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19896\ : std_logic;
signal \foc.Out_31__N_333_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19920\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Voltage_1_31\ : std_logic;
signal \foc.Out_31__N_332_cascade_\ : std_logic;
signal \foc.qVoltage_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18\ : std_logic;
signal \foc.qVoltage_14_cascade_\ : std_logic;
signal \foc.preSatVoltage_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_24\ : std_logic;
signal \foc.qVoltage_15\ : std_logic;
signal \bfn_21_17_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n57\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17736\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n108\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n106\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17737\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n155_adj_369\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n111\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17738\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n204_adj_361\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n114\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17739\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n253\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n117\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17740\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n302_adj_364\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n120\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17741\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n351\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n123\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17742\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17743\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n400_adj_511\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n126\ : std_logic;
signal \bfn_21_18_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n449_adj_492\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n129\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17744\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n498_adj_469\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n132\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17745\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n547_adj_454\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n135\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17746\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n596_adj_434\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n138\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17747\ : std_logic;
signal n141 : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n645_adj_429\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n691\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17748\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n694_adj_427\ : std_logic;
signal n146 : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n742\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17749\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n743\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_CO\ : std_logic;
signal \Saturate_out1_31__N_266_adj_2417\ : std_logic;
signal \Saturate_out1_31__N_267_adj_2418\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20660_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20654_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20640_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19308\ : std_logic;
signal \bfn_21_21_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n57\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18174\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n106\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18175\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n155\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18176\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n204\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18177\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n253\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18178\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n302\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18179\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n351\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18180\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18181\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n400\ : std_logic;
signal \bfn_21_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n449\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18182\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n498\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18183\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n547\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18184\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n596\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18185\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n645\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n691\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18186\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n694\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n742\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18187\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n743\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_0\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_4\ : std_logic;
signal \bfn_21_23_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_1\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15913\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15914\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15915\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_4\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15916\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15917\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15918\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15919\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15920\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_12\ : std_logic;
signal \bfn_21_24_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15921\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_14\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15922\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15923\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15924\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15925\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15926\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15927\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15928\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_20\ : std_logic;
signal \bfn_21_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_21\ : std_logic;
signal \Add_add_temp_21_adj_2399\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15929\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_22\ : std_logic;
signal \Add_add_temp_22_adj_2398\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15930\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_23\ : std_logic;
signal \Add_add_temp_23_adj_2397\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15931\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_24\ : std_logic;
signal \Add_add_temp_24_adj_2396\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15932\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_25\ : std_logic;
signal \Add_add_temp_25_adj_2395\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15933\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_26\ : std_logic;
signal \Add_add_temp_26_adj_2394\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15934\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_27\ : std_logic;
signal \Add_add_temp_27_adj_2393\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15935\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15936\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_28\ : std_logic;
signal \Add_add_temp_28_adj_2392\ : std_logic;
signal \bfn_21_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_29\ : std_logic;
signal \Add_add_temp_29_adj_2391\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15937\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_30\ : std_logic;
signal \Add_add_temp_30_adj_2390\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15938\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_27\ : std_logic;
signal \Add_add_temp_31_adj_2389\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15939\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28\ : std_logic;
signal \Add_add_temp_32_adj_2388\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15940\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_29\ : std_logic;
signal \Add_add_temp_33_adj_2387\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15941\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30\ : std_logic;
signal \Add_add_temp_34_adj_2386\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15942\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_31\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15943\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31\ : std_logic;
signal \bfn_21_28_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n81\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18294\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n130\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18295\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n179\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18296\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n228\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18297\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n277\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18298\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n326_adj_588\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18299\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n375_adj_587\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18300\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18301\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n424_adj_586\ : std_logic;
signal \bfn_21_29_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n473_adj_585\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18302\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n522_adj_584\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18303\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n571\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18304\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n620\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18305\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n669\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18306\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n718\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n774_adj_589\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18307\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n105\ : std_logic;
signal \bfn_22_11_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n57_adj_491\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17536\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n106_adj_509\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17537\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n155\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17538\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n204\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17539\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n253_adj_464\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17540\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n302\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17541\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n351_adj_396\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17542\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17543\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n400\ : std_logic;
signal \bfn_22_12_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n449\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17544\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n498\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17545\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n547\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17546\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n596\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17547\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n645\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17548\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n694\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n741\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n742_adj_411\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17549\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20550_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20556\ : std_logic;
signal \foc.dVoltage_5_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20554\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15_cascade_\ : std_logic;
signal \foc.dVoltage_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20560\ : std_logic;
signal \foc.Out_31__N_332_adj_2312_cascade_\ : std_logic;
signal \foc.dVoltage_8\ : std_logic;
signal \foc.Out_31__N_333_adj_2310_cascade_\ : std_logic;
signal \foc.dVoltage_14\ : std_logic;
signal \foc.dVoltage_3_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20572\ : std_logic;
signal \foc.dVoltage_11_cascade_\ : std_logic;
signal \foc.dVoltage_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20566\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11\ : std_logic;
signal \foc.qVoltage_2_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20594\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20612\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20618\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15\ : std_logic;
signal \foc.qVoltage_6\ : std_logic;
signal \foc.Out_31__N_332\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21\ : std_logic;
signal \foc.Out_31__N_333\ : std_logic;
signal \foc.qVoltage_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15264_cascade_\ : std_logic;
signal \Saturate_out1_31__N_267_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19842_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20666_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20658_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20648_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20634\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_0\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_4\ : std_logic;
signal \bfn_22_19_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_1\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15973\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15974\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15975\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15976\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15977\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15978\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15979\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15980\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_12\ : std_logic;
signal \bfn_22_20_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15981\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_14\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15982\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15983\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15984\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15985\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15986\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15987\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15988\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_20\ : std_logic;
signal \bfn_22_21_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15989\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15990\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15991\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_24\ : std_logic;
signal \Add_add_temp_24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15992\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15993\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15994\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15995\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15996\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_28\ : std_logic;
signal \Add_add_temp_28\ : std_logic;
signal \bfn_22_22_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_29\ : std_logic;
signal \Add_add_temp_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15997\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15998\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15999\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n16000\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n16001\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n16002\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_31\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n16003\ : std_logic;
signal \Add_add_temp_14_adj_2406\ : std_logic;
signal \Add_add_temp_12_adj_2408\ : std_logic;
signal \Add_add_temp_13_adj_2407\ : std_logic;
signal \Add_add_temp_16_adj_2404\ : std_logic;
signal \Add_add_temp_17_adj_2403\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n15200_cascade_\ : std_logic;
signal \Add_add_temp_15_adj_2405\ : std_logic;
signal \Add_add_temp_20_adj_2400\ : std_logic;
signal \Add_add_temp_19_adj_2401\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20680_cascade_\ : std_logic;
signal \Add_add_temp_18_adj_2402\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19733\ : std_logic;
signal \Add_add_temp_5_adj_2415\ : std_logic;
signal \Add_add_temp_4_adj_2416\ : std_logic;
signal \Add_add_temp_8_adj_2412\ : std_logic;
signal \Add_add_temp_7_adj_2413\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20722_cascade_\ : std_logic;
signal \Add_add_temp_6_adj_2414\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19761_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20704\ : std_logic;
signal \bfn_22_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n69\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n115\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18234\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n164\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18235\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n213\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18236\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n262\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18237\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n311\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18238\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n360\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18239\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n409\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18240\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18241\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n458\ : std_logic;
signal \bfn_22_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n507\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18242\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n556\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18243\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n605\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18244\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n654\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18245\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n703\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18246\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n758\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18247\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n759\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_CO\ : std_logic;
signal \bfn_22_28_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n78\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18279\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n127\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18280\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n176\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18281\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n225\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18282\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n274\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18283\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n323\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18284\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n372_adj_596\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18285\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18286\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n421_adj_595\ : std_logic;
signal \bfn_22_29_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n470_adj_594\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18287\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n519_adj_593\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18288\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n568_adj_592\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18289\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n617_adj_591\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18290\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n666\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18291\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n715\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n770\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18292\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n771\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n102\ : std_logic;
signal \bfn_23_11_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n54\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17521\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n103\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17522\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n152\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17523\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n201\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17524\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n250\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17525\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n299\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17526\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n348\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17527\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17528\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n397\ : std_logic;
signal \bfn_23_12_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n446\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17529\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n495\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17530\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n544\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17531\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n593\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17532\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n642\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17533\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n737\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n691_adj_440\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n738\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n17534\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n739\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19932\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20546\ : std_logic;
signal \foc.dVoltage_13_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20568_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20576\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n14\ : std_logic;
signal \foc.dVoltage_6\ : std_logic;
signal \foc.Out_31__N_332_adj_2312\ : std_logic;
signal \foc.Out_31__N_333_adj_2310\ : std_logic;
signal \foc.dVoltage_7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19747\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19858\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19904\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n22_cascade_\ : std_logic;
signal \Add_add_temp_31\ : std_logic;
signal \Add_add_temp_32\ : std_logic;
signal \Add_add_temp_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20644\ : std_logic;
signal \Add_add_temp_34\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n58_cascade_\ : std_logic;
signal \Add_add_temp_33\ : std_logic;
signal \Saturate_out1_31__N_266_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_4\ : std_logic;
signal \Add_add_temp_26\ : std_logic;
signal \Add_add_temp_27\ : std_logic;
signal \Add_add_temp_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_5\ : std_logic;
signal \Saturate_out1_31__N_267\ : std_logic;
signal \Saturate_out1_31__N_266\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19723_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20708_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n22_adj_519_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20688\ : std_logic;
signal \Add_add_temp_17\ : std_logic;
signal \Add_add_temp_16\ : std_logic;
signal \Add_add_temp_15\ : std_logic;
signal \Add_add_temp_5\ : std_logic;
signal \Add_add_temp_4\ : std_logic;
signal \Add_add_temp_8\ : std_logic;
signal \Add_add_temp_7\ : std_logic;
signal \Add_add_temp_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20712\ : std_logic;
signal \Add_add_temp_9\ : std_logic;
signal \Add_add_temp_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19777_cascade_\ : std_logic;
signal \Add_add_temp_10\ : std_logic;
signal \Add_add_temp_14\ : std_logic;
signal \Add_add_temp_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20700_cascade_\ : std_logic;
signal \Add_add_temp_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15205\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20670\ : std_logic;
signal \Add_add_temp_20\ : std_logic;
signal \Add_add_temp_18\ : std_logic;
signal \Add_add_temp_19\ : std_logic;
signal \Add_add_temp_21\ : std_logic;
signal \Add_add_temp_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n19746_cascade_\ : std_logic;
signal \Add_add_temp_22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20656\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31\ : std_logic;
signal \pin3_clk_16mhz_N\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n19755\ : std_logic;
signal \Add_add_temp_11_adj_2409\ : std_logic;
signal \Add_add_temp_9_adj_2411\ : std_logic;
signal \Add_add_temp_10_adj_2410\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n20718\ : std_logic;
signal \bfn_23_25_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n72\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n118\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18249\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n167\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18250\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n216\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18251\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n265\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18252\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n314\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18253\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n363\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18254\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n412\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18255\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18256\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n461\ : std_logic;
signal \bfn_23_26_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n510\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18257\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n559\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18258\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n608\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18259\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n657\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18260\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n706\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18261\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n762\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18262\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n763\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n102\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0\ : std_logic;
signal \bfn_23_27_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n75\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n105\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n121\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18264\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n124\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n108\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n170\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18265\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n173\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n111\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n219\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18266\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n222\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n114\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n268\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18267\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n271\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n317\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18268\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n120\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n320\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n366\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18269\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n369\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n123\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n415\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18270\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18271\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n126\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n418\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n464\ : std_logic;
signal \bfn_23_28_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n467\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n129\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n513\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18272\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n516\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n132\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n562\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18273\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n565\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n135\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n611\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18274\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n614\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n138\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n660\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18275\ : std_logic;
signal n141_adj_2421 : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n663\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n709\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18276\ : std_logic;
signal n146_adj_2423 : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n712\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n766\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n18277\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n767\ : std_logic;
signal \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19926\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20112_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20098\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15171_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15188_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19688_cascade_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19424\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n14851\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19455\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19690\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0\ : std_logic;
signal \bfn_24_16_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20184\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_1\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15568\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20186\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_2\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15569\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20188\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_3\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15570\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20190\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_4\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15571\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20192\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_5\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15572\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15573\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_0_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_1_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20194\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_6\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14\ : std_logic;
signal \bfn_24_17_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20196\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_7\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n20198\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15574\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_8\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15575\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_9\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17\ : std_logic;
signal \foc.preSatVoltage_10_adj_2311\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15576\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_10\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15577\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_11\ : std_logic;
signal \foc.preSatVoltage_12_adj_2330\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15578\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_12\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15579\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15580\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15580_THRU_CRY_0_THRU_CO\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_13\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14\ : std_logic;
signal \bfn_24_18_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_14\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15581\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_15\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15582\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_16\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15583\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_17\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15584\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_18\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26\ : std_logic;
signal \foc.preSatVoltage_19_adj_2329\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15585\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_19\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15586\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_20\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15587\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15588\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_21\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_22\ : std_logic;
signal \bfn_24_19_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_22\ : std_logic;
signal \foc.preSatVoltage_23_adj_2328\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15589\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_23\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15590\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_24\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15591\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_25\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15592\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_26\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15593\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_27\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15594\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_28\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15595\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15596\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_29\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30\ : std_logic;
signal \bfn_24_20_0_\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_30\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.n15597\ : std_logic;
signal \foc.u_DQ_Current_Control.u_D_Current_Control.Voltage_1_31\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal pin10_wire : std_logic;
signal pin11_wire : std_logic;
signal pin12_wire : std_logic;
signal pin13_wire : std_logic;
signal pin14_sdo_wire : std_logic;
signal pin15_sdi_wire : std_logic;
signal pin16_sck_wire : std_logic;
signal pin17_ss_wire : std_logic;
signal pin18_wire : std_logic;
signal pin19_wire : std_logic;
signal pin1_usb_dp_wire : std_logic;
signal pin20_wire : std_logic;
signal pin21_wire : std_logic;
signal pin22_wire : std_logic;
signal pin23_wire : std_logic;
signal pin24_wire : std_logic;
signal pin2_usb_dn_wire : std_logic;
signal pin7_wire : std_logic;
signal pin8_wire : std_logic;
signal pin9_wire : std_logic;
signal pin3_clk_16mhz_wire : std_logic;

begin
    pin10 <= pin10_wire;
    pin11 <= pin11_wire;
    pin12 <= pin12_wire;
    pin13 <= pin13_wire;
    pin14_sdo <= pin14_sdo_wire;
    pin15_sdi <= pin15_sdi_wire;
    pin16_sck <= pin16_sck_wire;
    pin17_ss <= pin17_ss_wire;
    pin18 <= pin18_wire;
    pin19 <= pin19_wire;
    pin1_usb_dp <= pin1_usb_dp_wire;
    pin20 <= pin20_wire;
    pin21 <= pin21_wire;
    pin22 <= pin22_wire;
    pin23 <= pin23_wire;
    pin24 <= pin24_wire;
    pin2_usb_dn <= pin2_usb_dn_wire;
    pin7 <= pin7_wire;
    pin8 <= pin8_wire;
    pin9 <= pin9_wire;
    pin3_clk_16mhz_wire <= pin3_clk_16mhz;

    \pin10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69497\,
            DIN => \N__69496\,
            DOUT => \N__69495\,
            PACKAGEPIN => pin10_wire
        );

    \pin10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69497\,
            PADOUT => \N__69496\,
            PADIN => \N__69495\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69488\,
            DIN => \N__69487\,
            DOUT => \N__69486\,
            PACKAGEPIN => pin11_wire
        );

    \pin11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69488\,
            PADOUT => \N__69487\,
            PADIN => \N__69486\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69479\,
            DIN => \N__69478\,
            DOUT => \N__69477\,
            PACKAGEPIN => pin12_wire
        );

    \pin12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69479\,
            PADOUT => \N__69478\,
            PADIN => \N__69477\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69470\,
            DIN => \N__69469\,
            DOUT => \N__69468\,
            PACKAGEPIN => pin13_wire
        );

    \pin13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69470\,
            PADOUT => \N__69469\,
            PADIN => \N__69468\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin14_sdo_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69461\,
            DIN => \N__69460\,
            DOUT => \N__69459\,
            PACKAGEPIN => pin14_sdo_wire
        );

    \pin14_sdo_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69461\,
            PADOUT => \N__69460\,
            PADIN => \N__69459\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin15_sdi_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69452\,
            DIN => \N__69451\,
            DOUT => \N__69450\,
            PACKAGEPIN => pin15_sdi_wire
        );

    \pin15_sdi_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69452\,
            PADOUT => \N__69451\,
            PADIN => \N__69450\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin16_sck_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69443\,
            DIN => \N__69442\,
            DOUT => \N__69441\,
            PACKAGEPIN => pin16_sck_wire
        );

    \pin16_sck_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69443\,
            PADOUT => \N__69442\,
            PADIN => \N__69441\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin17_ss_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69434\,
            DIN => \N__69433\,
            DOUT => \N__69432\,
            PACKAGEPIN => pin17_ss_wire
        );

    \pin17_ss_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69434\,
            PADOUT => \N__69433\,
            PADIN => \N__69432\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69425\,
            DIN => \N__69424\,
            DOUT => \N__69423\,
            PACKAGEPIN => pin18_wire
        );

    \pin18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69425\,
            PADOUT => \N__69424\,
            PADIN => \N__69423\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69416\,
            DIN => \N__69415\,
            DOUT => \N__69414\,
            PACKAGEPIN => pin19_wire
        );

    \pin19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69416\,
            PADOUT => \N__69415\,
            PADIN => \N__69414\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin1_usb_dp_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69407\,
            DIN => \N__69406\,
            DOUT => \N__69405\,
            PACKAGEPIN => pin1_usb_dp_wire
        );

    \pin1_usb_dp_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69407\,
            PADOUT => \N__69406\,
            PADIN => \N__69405\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69398\,
            DIN => \N__69397\,
            DOUT => \N__69396\,
            PACKAGEPIN => pin20_wire
        );

    \pin20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69398\,
            PADOUT => \N__69397\,
            PADIN => \N__69396\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69389\,
            DIN => \N__69388\,
            DOUT => \N__69387\,
            PACKAGEPIN => pin21_wire
        );

    \pin21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69389\,
            PADOUT => \N__69388\,
            PADIN => \N__69387\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69380\,
            DIN => \N__69379\,
            DOUT => \N__69378\,
            PACKAGEPIN => pin22_wire
        );

    \pin22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69380\,
            PADOUT => \N__69379\,
            PADIN => \N__69378\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69371\,
            DIN => \N__69370\,
            DOUT => \N__69369\,
            PACKAGEPIN => pin23_wire
        );

    \pin23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69371\,
            PADOUT => \N__69370\,
            PADIN => \N__69369\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69362\,
            DIN => \N__69361\,
            DOUT => \N__69360\,
            PACKAGEPIN => pin24_wire
        );

    \pin24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69362\,
            PADOUT => \N__69361\,
            PADIN => \N__69360\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin2_usb_dn_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69353\,
            DIN => \N__69352\,
            DOUT => \N__69351\,
            PACKAGEPIN => pin2_usb_dn_wire
        );

    \pin2_usb_dn_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69353\,
            PADOUT => \N__69352\,
            PADIN => \N__69351\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69344\,
            DIN => \N__69343\,
            DOUT => \N__69342\,
            PACKAGEPIN => pin7_wire
        );

    \pin7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69344\,
            PADOUT => \N__69343\,
            PADIN => \N__69342\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69335\,
            DIN => \N__69334\,
            DOUT => \N__69333\,
            PACKAGEPIN => pin8_wire
        );

    \pin8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69335\,
            PADOUT => \N__69334\,
            PADIN => \N__69333\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69326\,
            DIN => \N__69325\,
            DOUT => \N__69324\,
            PACKAGEPIN => pin9_wire
        );

    \pin9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69326\,
            PADOUT => \N__69325\,
            PADIN => \N__69324\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin3_clk_16mhz_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69317\,
            DIN => \N__69316\,
            DOUT => \N__69315\,
            PACKAGEPIN => pin3_clk_16mhz_wire
        );

    \pin3_clk_16mhz_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69317\,
            PADOUT => \N__69316\,
            PADIN => \N__69315\,
            CLOCKENABLE => 'H',
            DIN0 => pin3_clk_16mhz_pad_gb_input,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__15992\ : CascadeMux
    port map (
            O => \N__69298\,
            I => \N__69295\
        );

    \I__15991\ : InMux
    port map (
            O => \N__69295\,
            I => \N__69288\
        );

    \I__15990\ : InMux
    port map (
            O => \N__69294\,
            I => \N__69288\
        );

    \I__15989\ : InMux
    port map (
            O => \N__69293\,
            I => \N__69285\
        );

    \I__15988\ : LocalMux
    port map (
            O => \N__69288\,
            I => \N__69282\
        );

    \I__15987\ : LocalMux
    port map (
            O => \N__69285\,
            I => \N__69279\
        );

    \I__15986\ : Sp12to4
    port map (
            O => \N__69282\,
            I => \N__69276\
        );

    \I__15985\ : Span4Mux_h
    port map (
            O => \N__69279\,
            I => \N__69273\
        );

    \I__15984\ : Odrv12
    port map (
            O => \N__69276\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26\
        );

    \I__15983\ : Odrv4
    port map (
            O => \N__69273\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26\
        );

    \I__15982\ : InMux
    port map (
            O => \N__69268\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15592\
        );

    \I__15981\ : InMux
    port map (
            O => \N__69265\,
            I => \N__69262\
        );

    \I__15980\ : LocalMux
    port map (
            O => \N__69262\,
            I => \N__69259\
        );

    \I__15979\ : Span12Mux_v
    port map (
            O => \N__69259\,
            I => \N__69256\
        );

    \I__15978\ : Odrv12
    port map (
            O => \N__69256\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_26\
        );

    \I__15977\ : InMux
    port map (
            O => \N__69253\,
            I => \N__69246\
        );

    \I__15976\ : InMux
    port map (
            O => \N__69252\,
            I => \N__69246\
        );

    \I__15975\ : InMux
    port map (
            O => \N__69251\,
            I => \N__69243\
        );

    \I__15974\ : LocalMux
    port map (
            O => \N__69246\,
            I => \N__69240\
        );

    \I__15973\ : LocalMux
    port map (
            O => \N__69243\,
            I => \N__69237\
        );

    \I__15972\ : Span12Mux_v
    port map (
            O => \N__69240\,
            I => \N__69234\
        );

    \I__15971\ : Span4Mux_h
    port map (
            O => \N__69237\,
            I => \N__69231\
        );

    \I__15970\ : Odrv12
    port map (
            O => \N__69234\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27\
        );

    \I__15969\ : Odrv4
    port map (
            O => \N__69231\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27\
        );

    \I__15968\ : InMux
    port map (
            O => \N__69226\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15593\
        );

    \I__15967\ : CascadeMux
    port map (
            O => \N__69223\,
            I => \N__69220\
        );

    \I__15966\ : InMux
    port map (
            O => \N__69220\,
            I => \N__69217\
        );

    \I__15965\ : LocalMux
    port map (
            O => \N__69217\,
            I => \N__69214\
        );

    \I__15964\ : Span4Mux_v
    port map (
            O => \N__69214\,
            I => \N__69211\
        );

    \I__15963\ : Odrv4
    port map (
            O => \N__69211\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_27\
        );

    \I__15962\ : InMux
    port map (
            O => \N__69208\,
            I => \N__69205\
        );

    \I__15961\ : LocalMux
    port map (
            O => \N__69205\,
            I => \N__69200\
        );

    \I__15960\ : InMux
    port map (
            O => \N__69204\,
            I => \N__69197\
        );

    \I__15959\ : InMux
    port map (
            O => \N__69203\,
            I => \N__69194\
        );

    \I__15958\ : Span4Mux_v
    port map (
            O => \N__69200\,
            I => \N__69191\
        );

    \I__15957\ : LocalMux
    port map (
            O => \N__69197\,
            I => \N__69186\
        );

    \I__15956\ : LocalMux
    port map (
            O => \N__69194\,
            I => \N__69186\
        );

    \I__15955\ : Span4Mux_h
    port map (
            O => \N__69191\,
            I => \N__69183\
        );

    \I__15954\ : Span4Mux_v
    port map (
            O => \N__69186\,
            I => \N__69180\
        );

    \I__15953\ : Odrv4
    port map (
            O => \N__69183\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28\
        );

    \I__15952\ : Odrv4
    port map (
            O => \N__69180\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28\
        );

    \I__15951\ : InMux
    port map (
            O => \N__69175\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15594\
        );

    \I__15950\ : InMux
    port map (
            O => \N__69172\,
            I => \N__69169\
        );

    \I__15949\ : LocalMux
    port map (
            O => \N__69169\,
            I => \N__69166\
        );

    \I__15948\ : Span4Mux_v
    port map (
            O => \N__69166\,
            I => \N__69163\
        );

    \I__15947\ : Span4Mux_h
    port map (
            O => \N__69163\,
            I => \N__69160\
        );

    \I__15946\ : Odrv4
    port map (
            O => \N__69160\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_28\
        );

    \I__15945\ : InMux
    port map (
            O => \N__69157\,
            I => \N__69150\
        );

    \I__15944\ : InMux
    port map (
            O => \N__69156\,
            I => \N__69150\
        );

    \I__15943\ : CascadeMux
    port map (
            O => \N__69155\,
            I => \N__69147\
        );

    \I__15942\ : LocalMux
    port map (
            O => \N__69150\,
            I => \N__69144\
        );

    \I__15941\ : InMux
    port map (
            O => \N__69147\,
            I => \N__69141\
        );

    \I__15940\ : Span4Mux_h
    port map (
            O => \N__69144\,
            I => \N__69136\
        );

    \I__15939\ : LocalMux
    port map (
            O => \N__69141\,
            I => \N__69136\
        );

    \I__15938\ : Sp12to4
    port map (
            O => \N__69136\,
            I => \N__69133\
        );

    \I__15937\ : Odrv12
    port map (
            O => \N__69133\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_29\
        );

    \I__15936\ : InMux
    port map (
            O => \N__69130\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15595\
        );

    \I__15935\ : CascadeMux
    port map (
            O => \N__69127\,
            I => \N__69124\
        );

    \I__15934\ : InMux
    port map (
            O => \N__69124\,
            I => \N__69121\
        );

    \I__15933\ : LocalMux
    port map (
            O => \N__69121\,
            I => \N__69118\
        );

    \I__15932\ : Span4Mux_h
    port map (
            O => \N__69118\,
            I => \N__69115\
        );

    \I__15931\ : Span4Mux_v
    port map (
            O => \N__69115\,
            I => \N__69112\
        );

    \I__15930\ : Odrv4
    port map (
            O => \N__69112\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_29\
        );

    \I__15929\ : InMux
    port map (
            O => \N__69109\,
            I => \N__69102\
        );

    \I__15928\ : InMux
    port map (
            O => \N__69108\,
            I => \N__69102\
        );

    \I__15927\ : InMux
    port map (
            O => \N__69107\,
            I => \N__69099\
        );

    \I__15926\ : LocalMux
    port map (
            O => \N__69102\,
            I => \N__69096\
        );

    \I__15925\ : LocalMux
    port map (
            O => \N__69099\,
            I => \N__69093\
        );

    \I__15924\ : Span4Mux_h
    port map (
            O => \N__69096\,
            I => \N__69090\
        );

    \I__15923\ : Span4Mux_h
    port map (
            O => \N__69093\,
            I => \N__69087\
        );

    \I__15922\ : Span4Mux_v
    port map (
            O => \N__69090\,
            I => \N__69084\
        );

    \I__15921\ : Span4Mux_v
    port map (
            O => \N__69087\,
            I => \N__69081\
        );

    \I__15920\ : Odrv4
    port map (
            O => \N__69084\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30\
        );

    \I__15919\ : Odrv4
    port map (
            O => \N__69081\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30\
        );

    \I__15918\ : InMux
    port map (
            O => \N__69076\,
            I => \bfn_24_20_0_\
        );

    \I__15917\ : CascadeMux
    port map (
            O => \N__69073\,
            I => \N__69068\
        );

    \I__15916\ : CascadeMux
    port map (
            O => \N__69072\,
            I => \N__69064\
        );

    \I__15915\ : CascadeMux
    port map (
            O => \N__69071\,
            I => \N__69060\
        );

    \I__15914\ : InMux
    port map (
            O => \N__69068\,
            I => \N__69046\
        );

    \I__15913\ : InMux
    port map (
            O => \N__69067\,
            I => \N__69046\
        );

    \I__15912\ : InMux
    port map (
            O => \N__69064\,
            I => \N__69046\
        );

    \I__15911\ : InMux
    port map (
            O => \N__69063\,
            I => \N__69046\
        );

    \I__15910\ : InMux
    port map (
            O => \N__69060\,
            I => \N__69046\
        );

    \I__15909\ : InMux
    port map (
            O => \N__69059\,
            I => \N__69046\
        );

    \I__15908\ : LocalMux
    port map (
            O => \N__69046\,
            I => \N__69040\
        );

    \I__15907\ : InMux
    port map (
            O => \N__69045\,
            I => \N__69037\
        );

    \I__15906\ : InMux
    port map (
            O => \N__69044\,
            I => \N__69032\
        );

    \I__15905\ : InMux
    port map (
            O => \N__69043\,
            I => \N__69032\
        );

    \I__15904\ : Odrv4
    port map (
            O => \N__69040\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31\
        );

    \I__15903\ : LocalMux
    port map (
            O => \N__69037\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31\
        );

    \I__15902\ : LocalMux
    port map (
            O => \N__69032\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31\
        );

    \I__15901\ : InMux
    port map (
            O => \N__69025\,
            I => \N__69022\
        );

    \I__15900\ : LocalMux
    port map (
            O => \N__69022\,
            I => \N__69019\
        );

    \I__15899\ : Span4Mux_v
    port map (
            O => \N__69019\,
            I => \N__69016\
        );

    \I__15898\ : Odrv4
    port map (
            O => \N__69016\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_30\
        );

    \I__15897\ : InMux
    port map (
            O => \N__69013\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15597\
        );

    \I__15896\ : CascadeMux
    port map (
            O => \N__69010\,
            I => \N__69007\
        );

    \I__15895\ : InMux
    port map (
            O => \N__69007\,
            I => \N__69003\
        );

    \I__15894\ : CascadeMux
    port map (
            O => \N__69006\,
            I => \N__69000\
        );

    \I__15893\ : LocalMux
    port map (
            O => \N__69003\,
            I => \N__68997\
        );

    \I__15892\ : InMux
    port map (
            O => \N__69000\,
            I => \N__68994\
        );

    \I__15891\ : Span4Mux_v
    port map (
            O => \N__68997\,
            I => \N__68991\
        );

    \I__15890\ : LocalMux
    port map (
            O => \N__68994\,
            I => \N__68988\
        );

    \I__15889\ : Span4Mux_h
    port map (
            O => \N__68991\,
            I => \N__68983\
        );

    \I__15888\ : Span4Mux_v
    port map (
            O => \N__68988\,
            I => \N__68983\
        );

    \I__15887\ : Span4Mux_v
    port map (
            O => \N__68983\,
            I => \N__68980\
        );

    \I__15886\ : Odrv4
    port map (
            O => \N__68980\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Voltage_1_31\
        );

    \I__15885\ : InMux
    port map (
            O => \N__68977\,
            I => \N__68974\
        );

    \I__15884\ : LocalMux
    port map (
            O => \N__68974\,
            I => \N__68971\
        );

    \I__15883\ : Span4Mux_v
    port map (
            O => \N__68971\,
            I => \N__68968\
        );

    \I__15882\ : Odrv4
    port map (
            O => \N__68968\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_18\
        );

    \I__15881\ : InMux
    port map (
            O => \N__68965\,
            I => \N__68962\
        );

    \I__15880\ : LocalMux
    port map (
            O => \N__68962\,
            I => \N__68958\
        );

    \I__15879\ : CascadeMux
    port map (
            O => \N__68961\,
            I => \N__68955\
        );

    \I__15878\ : Sp12to4
    port map (
            O => \N__68958\,
            I => \N__68952\
        );

    \I__15877\ : InMux
    port map (
            O => \N__68955\,
            I => \N__68949\
        );

    \I__15876\ : Odrv12
    port map (
            O => \N__68952\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26\
        );

    \I__15875\ : LocalMux
    port map (
            O => \N__68949\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26\
        );

    \I__15874\ : InMux
    port map (
            O => \N__68944\,
            I => \N__68937\
        );

    \I__15873\ : InMux
    port map (
            O => \N__68943\,
            I => \N__68937\
        );

    \I__15872\ : InMux
    port map (
            O => \N__68942\,
            I => \N__68933\
        );

    \I__15871\ : LocalMux
    port map (
            O => \N__68937\,
            I => \N__68930\
        );

    \I__15870\ : InMux
    port map (
            O => \N__68936\,
            I => \N__68927\
        );

    \I__15869\ : LocalMux
    port map (
            O => \N__68933\,
            I => \N__68924\
        );

    \I__15868\ : Span4Mux_h
    port map (
            O => \N__68930\,
            I => \N__68919\
        );

    \I__15867\ : LocalMux
    port map (
            O => \N__68927\,
            I => \N__68919\
        );

    \I__15866\ : Odrv12
    port map (
            O => \N__68924\,
            I => \foc.preSatVoltage_19_adj_2329\
        );

    \I__15865\ : Odrv4
    port map (
            O => \N__68919\,
            I => \foc.preSatVoltage_19_adj_2329\
        );

    \I__15864\ : InMux
    port map (
            O => \N__68914\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15585\
        );

    \I__15863\ : InMux
    port map (
            O => \N__68911\,
            I => \N__68907\
        );

    \I__15862\ : InMux
    port map (
            O => \N__68910\,
            I => \N__68904\
        );

    \I__15861\ : LocalMux
    port map (
            O => \N__68907\,
            I => \N__68901\
        );

    \I__15860\ : LocalMux
    port map (
            O => \N__68904\,
            I => \N__68898\
        );

    \I__15859\ : Span4Mux_v
    port map (
            O => \N__68901\,
            I => \N__68895\
        );

    \I__15858\ : Odrv12
    port map (
            O => \N__68898\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27\
        );

    \I__15857\ : Odrv4
    port map (
            O => \N__68895\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27\
        );

    \I__15856\ : CascadeMux
    port map (
            O => \N__68890\,
            I => \N__68887\
        );

    \I__15855\ : InMux
    port map (
            O => \N__68887\,
            I => \N__68884\
        );

    \I__15854\ : LocalMux
    port map (
            O => \N__68884\,
            I => \N__68881\
        );

    \I__15853\ : Span4Mux_v
    port map (
            O => \N__68881\,
            I => \N__68878\
        );

    \I__15852\ : Span4Mux_h
    port map (
            O => \N__68878\,
            I => \N__68875\
        );

    \I__15851\ : Odrv4
    port map (
            O => \N__68875\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_19\
        );

    \I__15850\ : InMux
    port map (
            O => \N__68872\,
            I => \N__68866\
        );

    \I__15849\ : InMux
    port map (
            O => \N__68871\,
            I => \N__68866\
        );

    \I__15848\ : LocalMux
    port map (
            O => \N__68866\,
            I => \N__68863\
        );

    \I__15847\ : Span4Mux_h
    port map (
            O => \N__68863\,
            I => \N__68858\
        );

    \I__15846\ : InMux
    port map (
            O => \N__68862\,
            I => \N__68855\
        );

    \I__15845\ : InMux
    port map (
            O => \N__68861\,
            I => \N__68852\
        );

    \I__15844\ : Sp12to4
    port map (
            O => \N__68858\,
            I => \N__68845\
        );

    \I__15843\ : LocalMux
    port map (
            O => \N__68855\,
            I => \N__68845\
        );

    \I__15842\ : LocalMux
    port map (
            O => \N__68852\,
            I => \N__68845\
        );

    \I__15841\ : Odrv12
    port map (
            O => \N__68845\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_20\
        );

    \I__15840\ : InMux
    port map (
            O => \N__68842\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15586\
        );

    \I__15839\ : CascadeMux
    port map (
            O => \N__68839\,
            I => \N__68836\
        );

    \I__15838\ : InMux
    port map (
            O => \N__68836\,
            I => \N__68833\
        );

    \I__15837\ : LocalMux
    port map (
            O => \N__68833\,
            I => \N__68830\
        );

    \I__15836\ : Span4Mux_v
    port map (
            O => \N__68830\,
            I => \N__68826\
        );

    \I__15835\ : InMux
    port map (
            O => \N__68829\,
            I => \N__68823\
        );

    \I__15834\ : Odrv4
    port map (
            O => \N__68826\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28\
        );

    \I__15833\ : LocalMux
    port map (
            O => \N__68823\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28\
        );

    \I__15832\ : CascadeMux
    port map (
            O => \N__68818\,
            I => \N__68815\
        );

    \I__15831\ : InMux
    port map (
            O => \N__68815\,
            I => \N__68812\
        );

    \I__15830\ : LocalMux
    port map (
            O => \N__68812\,
            I => \N__68809\
        );

    \I__15829\ : Span4Mux_h
    port map (
            O => \N__68809\,
            I => \N__68806\
        );

    \I__15828\ : Span4Mux_v
    port map (
            O => \N__68806\,
            I => \N__68803\
        );

    \I__15827\ : Odrv4
    port map (
            O => \N__68803\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_20\
        );

    \I__15826\ : InMux
    port map (
            O => \N__68800\,
            I => \N__68794\
        );

    \I__15825\ : InMux
    port map (
            O => \N__68799\,
            I => \N__68794\
        );

    \I__15824\ : LocalMux
    port map (
            O => \N__68794\,
            I => \N__68789\
        );

    \I__15823\ : InMux
    port map (
            O => \N__68793\,
            I => \N__68786\
        );

    \I__15822\ : InMux
    port map (
            O => \N__68792\,
            I => \N__68783\
        );

    \I__15821\ : Span12Mux_h
    port map (
            O => \N__68789\,
            I => \N__68776\
        );

    \I__15820\ : LocalMux
    port map (
            O => \N__68786\,
            I => \N__68776\
        );

    \I__15819\ : LocalMux
    port map (
            O => \N__68783\,
            I => \N__68776\
        );

    \I__15818\ : Odrv12
    port map (
            O => \N__68776\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_21\
        );

    \I__15817\ : InMux
    port map (
            O => \N__68773\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15587\
        );

    \I__15816\ : CascadeMux
    port map (
            O => \N__68770\,
            I => \N__68766\
        );

    \I__15815\ : InMux
    port map (
            O => \N__68769\,
            I => \N__68763\
        );

    \I__15814\ : InMux
    port map (
            O => \N__68766\,
            I => \N__68760\
        );

    \I__15813\ : LocalMux
    port map (
            O => \N__68763\,
            I => \N__68757\
        );

    \I__15812\ : LocalMux
    port map (
            O => \N__68760\,
            I => \N__68754\
        );

    \I__15811\ : Span4Mux_v
    port map (
            O => \N__68757\,
            I => \N__68751\
        );

    \I__15810\ : Odrv12
    port map (
            O => \N__68754\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29\
        );

    \I__15809\ : Odrv4
    port map (
            O => \N__68751\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29\
        );

    \I__15808\ : CascadeMux
    port map (
            O => \N__68746\,
            I => \N__68743\
        );

    \I__15807\ : InMux
    port map (
            O => \N__68743\,
            I => \N__68740\
        );

    \I__15806\ : LocalMux
    port map (
            O => \N__68740\,
            I => \N__68737\
        );

    \I__15805\ : Span4Mux_v
    port map (
            O => \N__68737\,
            I => \N__68734\
        );

    \I__15804\ : Span4Mux_h
    port map (
            O => \N__68734\,
            I => \N__68731\
        );

    \I__15803\ : Odrv4
    port map (
            O => \N__68731\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_21\
        );

    \I__15802\ : InMux
    port map (
            O => \N__68728\,
            I => \N__68722\
        );

    \I__15801\ : InMux
    port map (
            O => \N__68727\,
            I => \N__68722\
        );

    \I__15800\ : LocalMux
    port map (
            O => \N__68722\,
            I => \N__68717\
        );

    \I__15799\ : InMux
    port map (
            O => \N__68721\,
            I => \N__68714\
        );

    \I__15798\ : InMux
    port map (
            O => \N__68720\,
            I => \N__68711\
        );

    \I__15797\ : Sp12to4
    port map (
            O => \N__68717\,
            I => \N__68704\
        );

    \I__15796\ : LocalMux
    port map (
            O => \N__68714\,
            I => \N__68704\
        );

    \I__15795\ : LocalMux
    port map (
            O => \N__68711\,
            I => \N__68704\
        );

    \I__15794\ : Odrv12
    port map (
            O => \N__68704\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_22\
        );

    \I__15793\ : InMux
    port map (
            O => \N__68701\,
            I => \bfn_24_19_0_\
        );

    \I__15792\ : InMux
    port map (
            O => \N__68698\,
            I => \N__68694\
        );

    \I__15791\ : InMux
    port map (
            O => \N__68697\,
            I => \N__68691\
        );

    \I__15790\ : LocalMux
    port map (
            O => \N__68694\,
            I => \N__68688\
        );

    \I__15789\ : LocalMux
    port map (
            O => \N__68691\,
            I => \N__68685\
        );

    \I__15788\ : Span4Mux_v
    port map (
            O => \N__68688\,
            I => \N__68682\
        );

    \I__15787\ : Span4Mux_v
    port map (
            O => \N__68685\,
            I => \N__68679\
        );

    \I__15786\ : Odrv4
    port map (
            O => \N__68682\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30\
        );

    \I__15785\ : Odrv4
    port map (
            O => \N__68679\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30\
        );

    \I__15784\ : CascadeMux
    port map (
            O => \N__68674\,
            I => \N__68671\
        );

    \I__15783\ : InMux
    port map (
            O => \N__68671\,
            I => \N__68668\
        );

    \I__15782\ : LocalMux
    port map (
            O => \N__68668\,
            I => \N__68665\
        );

    \I__15781\ : Span4Mux_v
    port map (
            O => \N__68665\,
            I => \N__68662\
        );

    \I__15780\ : Odrv4
    port map (
            O => \N__68662\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_22\
        );

    \I__15779\ : InMux
    port map (
            O => \N__68659\,
            I => \N__68653\
        );

    \I__15778\ : InMux
    port map (
            O => \N__68658\,
            I => \N__68653\
        );

    \I__15777\ : LocalMux
    port map (
            O => \N__68653\,
            I => \N__68650\
        );

    \I__15776\ : Span4Mux_v
    port map (
            O => \N__68650\,
            I => \N__68645\
        );

    \I__15775\ : InMux
    port map (
            O => \N__68649\,
            I => \N__68642\
        );

    \I__15774\ : InMux
    port map (
            O => \N__68648\,
            I => \N__68639\
        );

    \I__15773\ : Span4Mux_v
    port map (
            O => \N__68645\,
            I => \N__68636\
        );

    \I__15772\ : LocalMux
    port map (
            O => \N__68642\,
            I => \N__68631\
        );

    \I__15771\ : LocalMux
    port map (
            O => \N__68639\,
            I => \N__68631\
        );

    \I__15770\ : Odrv4
    port map (
            O => \N__68636\,
            I => \foc.preSatVoltage_23_adj_2328\
        );

    \I__15769\ : Odrv12
    port map (
            O => \N__68631\,
            I => \foc.preSatVoltage_23_adj_2328\
        );

    \I__15768\ : InMux
    port map (
            O => \N__68626\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15589\
        );

    \I__15767\ : CascadeMux
    port map (
            O => \N__68623\,
            I => \N__68620\
        );

    \I__15766\ : InMux
    port map (
            O => \N__68620\,
            I => \N__68617\
        );

    \I__15765\ : LocalMux
    port map (
            O => \N__68617\,
            I => \N__68614\
        );

    \I__15764\ : Span4Mux_v
    port map (
            O => \N__68614\,
            I => \N__68611\
        );

    \I__15763\ : Odrv4
    port map (
            O => \N__68611\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_23\
        );

    \I__15762\ : InMux
    port map (
            O => \N__68608\,
            I => \N__68602\
        );

    \I__15761\ : InMux
    port map (
            O => \N__68607\,
            I => \N__68602\
        );

    \I__15760\ : LocalMux
    port map (
            O => \N__68602\,
            I => \N__68598\
        );

    \I__15759\ : InMux
    port map (
            O => \N__68601\,
            I => \N__68595\
        );

    \I__15758\ : Span4Mux_v
    port map (
            O => \N__68598\,
            I => \N__68591\
        );

    \I__15757\ : LocalMux
    port map (
            O => \N__68595\,
            I => \N__68588\
        );

    \I__15756\ : InMux
    port map (
            O => \N__68594\,
            I => \N__68585\
        );

    \I__15755\ : Span4Mux_h
    port map (
            O => \N__68591\,
            I => \N__68582\
        );

    \I__15754\ : Sp12to4
    port map (
            O => \N__68588\,
            I => \N__68577\
        );

    \I__15753\ : LocalMux
    port map (
            O => \N__68585\,
            I => \N__68577\
        );

    \I__15752\ : Odrv4
    port map (
            O => \N__68582\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24\
        );

    \I__15751\ : Odrv12
    port map (
            O => \N__68577\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24\
        );

    \I__15750\ : InMux
    port map (
            O => \N__68572\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15590\
        );

    \I__15749\ : InMux
    port map (
            O => \N__68569\,
            I => \N__68566\
        );

    \I__15748\ : LocalMux
    port map (
            O => \N__68566\,
            I => \N__68563\
        );

    \I__15747\ : Span4Mux_v
    port map (
            O => \N__68563\,
            I => \N__68560\
        );

    \I__15746\ : Odrv4
    port map (
            O => \N__68560\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_24\
        );

    \I__15745\ : CascadeMux
    port map (
            O => \N__68557\,
            I => \N__68554\
        );

    \I__15744\ : InMux
    port map (
            O => \N__68554\,
            I => \N__68551\
        );

    \I__15743\ : LocalMux
    port map (
            O => \N__68551\,
            I => \N__68546\
        );

    \I__15742\ : InMux
    port map (
            O => \N__68550\,
            I => \N__68543\
        );

    \I__15741\ : CascadeMux
    port map (
            O => \N__68549\,
            I => \N__68540\
        );

    \I__15740\ : Span4Mux_v
    port map (
            O => \N__68546\,
            I => \N__68537\
        );

    \I__15739\ : LocalMux
    port map (
            O => \N__68543\,
            I => \N__68534\
        );

    \I__15738\ : InMux
    port map (
            O => \N__68540\,
            I => \N__68531\
        );

    \I__15737\ : Span4Mux_h
    port map (
            O => \N__68537\,
            I => \N__68528\
        );

    \I__15736\ : Sp12to4
    port map (
            O => \N__68534\,
            I => \N__68523\
        );

    \I__15735\ : LocalMux
    port map (
            O => \N__68531\,
            I => \N__68523\
        );

    \I__15734\ : Odrv4
    port map (
            O => \N__68528\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25\
        );

    \I__15733\ : Odrv12
    port map (
            O => \N__68523\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25\
        );

    \I__15732\ : InMux
    port map (
            O => \N__68518\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15591\
        );

    \I__15731\ : CascadeMux
    port map (
            O => \N__68515\,
            I => \N__68512\
        );

    \I__15730\ : InMux
    port map (
            O => \N__68512\,
            I => \N__68509\
        );

    \I__15729\ : LocalMux
    port map (
            O => \N__68509\,
            I => \N__68506\
        );

    \I__15728\ : Span4Mux_v
    port map (
            O => \N__68506\,
            I => \N__68503\
        );

    \I__15727\ : Odrv4
    port map (
            O => \N__68503\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_25\
        );

    \I__15726\ : CascadeMux
    port map (
            O => \N__68500\,
            I => \N__68497\
        );

    \I__15725\ : InMux
    port map (
            O => \N__68497\,
            I => \N__68493\
        );

    \I__15724\ : InMux
    port map (
            O => \N__68496\,
            I => \N__68490\
        );

    \I__15723\ : LocalMux
    port map (
            O => \N__68493\,
            I => \N__68487\
        );

    \I__15722\ : LocalMux
    port map (
            O => \N__68490\,
            I => \N__68484\
        );

    \I__15721\ : Odrv12
    port map (
            O => \N__68487\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20\
        );

    \I__15720\ : Odrv12
    port map (
            O => \N__68484\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20\
        );

    \I__15719\ : CascadeMux
    port map (
            O => \N__68479\,
            I => \N__68476\
        );

    \I__15718\ : InMux
    port map (
            O => \N__68476\,
            I => \N__68473\
        );

    \I__15717\ : LocalMux
    port map (
            O => \N__68473\,
            I => \N__68470\
        );

    \I__15716\ : Span4Mux_v
    port map (
            O => \N__68470\,
            I => \N__68467\
        );

    \I__15715\ : Odrv4
    port map (
            O => \N__68467\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_12\
        );

    \I__15714\ : InMux
    port map (
            O => \N__68464\,
            I => \N__68461\
        );

    \I__15713\ : LocalMux
    port map (
            O => \N__68461\,
            I => \N__68456\
        );

    \I__15712\ : InMux
    port map (
            O => \N__68460\,
            I => \N__68453\
        );

    \I__15711\ : InMux
    port map (
            O => \N__68459\,
            I => \N__68450\
        );

    \I__15710\ : Span4Mux_h
    port map (
            O => \N__68456\,
            I => \N__68445\
        );

    \I__15709\ : LocalMux
    port map (
            O => \N__68453\,
            I => \N__68445\
        );

    \I__15708\ : LocalMux
    port map (
            O => \N__68450\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13\
        );

    \I__15707\ : Odrv4
    port map (
            O => \N__68445\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13\
        );

    \I__15706\ : InMux
    port map (
            O => \N__68440\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15579\
        );

    \I__15705\ : InMux
    port map (
            O => \N__68437\,
            I => \N__68429\
        );

    \I__15704\ : InMux
    port map (
            O => \N__68436\,
            I => \N__68429\
        );

    \I__15703\ : InMux
    port map (
            O => \N__68435\,
            I => \N__68423\
        );

    \I__15702\ : CascadeMux
    port map (
            O => \N__68434\,
            I => \N__68419\
        );

    \I__15701\ : LocalMux
    port map (
            O => \N__68429\,
            I => \N__68415\
        );

    \I__15700\ : InMux
    port map (
            O => \N__68428\,
            I => \N__68412\
        );

    \I__15699\ : CascadeMux
    port map (
            O => \N__68427\,
            I => \N__68408\
        );

    \I__15698\ : CascadeMux
    port map (
            O => \N__68426\,
            I => \N__68404\
        );

    \I__15697\ : LocalMux
    port map (
            O => \N__68423\,
            I => \N__68387\
        );

    \I__15696\ : InMux
    port map (
            O => \N__68422\,
            I => \N__68384\
        );

    \I__15695\ : InMux
    port map (
            O => \N__68419\,
            I => \N__68379\
        );

    \I__15694\ : InMux
    port map (
            O => \N__68418\,
            I => \N__68379\
        );

    \I__15693\ : Span4Mux_v
    port map (
            O => \N__68415\,
            I => \N__68374\
        );

    \I__15692\ : LocalMux
    port map (
            O => \N__68412\,
            I => \N__68374\
        );

    \I__15691\ : InMux
    port map (
            O => \N__68411\,
            I => \N__68365\
        );

    \I__15690\ : InMux
    port map (
            O => \N__68408\,
            I => \N__68365\
        );

    \I__15689\ : InMux
    port map (
            O => \N__68407\,
            I => \N__68365\
        );

    \I__15688\ : InMux
    port map (
            O => \N__68404\,
            I => \N__68365\
        );

    \I__15687\ : CascadeMux
    port map (
            O => \N__68403\,
            I => \N__68361\
        );

    \I__15686\ : CascadeMux
    port map (
            O => \N__68402\,
            I => \N__68357\
        );

    \I__15685\ : CascadeMux
    port map (
            O => \N__68401\,
            I => \N__68353\
        );

    \I__15684\ : CascadeMux
    port map (
            O => \N__68400\,
            I => \N__68349\
        );

    \I__15683\ : CascadeMux
    port map (
            O => \N__68399\,
            I => \N__68345\
        );

    \I__15682\ : CascadeMux
    port map (
            O => \N__68398\,
            I => \N__68341\
        );

    \I__15681\ : CascadeMux
    port map (
            O => \N__68397\,
            I => \N__68337\
        );

    \I__15680\ : CascadeMux
    port map (
            O => \N__68396\,
            I => \N__68333\
        );

    \I__15679\ : CascadeMux
    port map (
            O => \N__68395\,
            I => \N__68329\
        );

    \I__15678\ : CascadeMux
    port map (
            O => \N__68394\,
            I => \N__68326\
        );

    \I__15677\ : CascadeMux
    port map (
            O => \N__68393\,
            I => \N__68323\
        );

    \I__15676\ : CascadeMux
    port map (
            O => \N__68392\,
            I => \N__68320\
        );

    \I__15675\ : CascadeMux
    port map (
            O => \N__68391\,
            I => \N__68317\
        );

    \I__15674\ : CascadeMux
    port map (
            O => \N__68390\,
            I => \N__68314\
        );

    \I__15673\ : Span4Mux_v
    port map (
            O => \N__68387\,
            I => \N__68311\
        );

    \I__15672\ : LocalMux
    port map (
            O => \N__68384\,
            I => \N__68306\
        );

    \I__15671\ : LocalMux
    port map (
            O => \N__68379\,
            I => \N__68306\
        );

    \I__15670\ : Span4Mux_v
    port map (
            O => \N__68374\,
            I => \N__68303\
        );

    \I__15669\ : LocalMux
    port map (
            O => \N__68365\,
            I => \N__68300\
        );

    \I__15668\ : InMux
    port map (
            O => \N__68364\,
            I => \N__68283\
        );

    \I__15667\ : InMux
    port map (
            O => \N__68361\,
            I => \N__68283\
        );

    \I__15666\ : InMux
    port map (
            O => \N__68360\,
            I => \N__68283\
        );

    \I__15665\ : InMux
    port map (
            O => \N__68357\,
            I => \N__68283\
        );

    \I__15664\ : InMux
    port map (
            O => \N__68356\,
            I => \N__68283\
        );

    \I__15663\ : InMux
    port map (
            O => \N__68353\,
            I => \N__68283\
        );

    \I__15662\ : InMux
    port map (
            O => \N__68352\,
            I => \N__68283\
        );

    \I__15661\ : InMux
    port map (
            O => \N__68349\,
            I => \N__68283\
        );

    \I__15660\ : InMux
    port map (
            O => \N__68348\,
            I => \N__68266\
        );

    \I__15659\ : InMux
    port map (
            O => \N__68345\,
            I => \N__68266\
        );

    \I__15658\ : InMux
    port map (
            O => \N__68344\,
            I => \N__68266\
        );

    \I__15657\ : InMux
    port map (
            O => \N__68341\,
            I => \N__68266\
        );

    \I__15656\ : InMux
    port map (
            O => \N__68340\,
            I => \N__68266\
        );

    \I__15655\ : InMux
    port map (
            O => \N__68337\,
            I => \N__68266\
        );

    \I__15654\ : InMux
    port map (
            O => \N__68336\,
            I => \N__68266\
        );

    \I__15653\ : InMux
    port map (
            O => \N__68333\,
            I => \N__68266\
        );

    \I__15652\ : InMux
    port map (
            O => \N__68332\,
            I => \N__68257\
        );

    \I__15651\ : InMux
    port map (
            O => \N__68329\,
            I => \N__68257\
        );

    \I__15650\ : InMux
    port map (
            O => \N__68326\,
            I => \N__68257\
        );

    \I__15649\ : InMux
    port map (
            O => \N__68323\,
            I => \N__68257\
        );

    \I__15648\ : InMux
    port map (
            O => \N__68320\,
            I => \N__68250\
        );

    \I__15647\ : InMux
    port map (
            O => \N__68317\,
            I => \N__68250\
        );

    \I__15646\ : InMux
    port map (
            O => \N__68314\,
            I => \N__68250\
        );

    \I__15645\ : Span4Mux_v
    port map (
            O => \N__68311\,
            I => \N__68247\
        );

    \I__15644\ : Span4Mux_v
    port map (
            O => \N__68306\,
            I => \N__68244\
        );

    \I__15643\ : Span4Mux_h
    port map (
            O => \N__68303\,
            I => \N__68231\
        );

    \I__15642\ : Span4Mux_v
    port map (
            O => \N__68300\,
            I => \N__68231\
        );

    \I__15641\ : LocalMux
    port map (
            O => \N__68283\,
            I => \N__68231\
        );

    \I__15640\ : LocalMux
    port map (
            O => \N__68266\,
            I => \N__68231\
        );

    \I__15639\ : LocalMux
    port map (
            O => \N__68257\,
            I => \N__68231\
        );

    \I__15638\ : LocalMux
    port map (
            O => \N__68250\,
            I => \N__68231\
        );

    \I__15637\ : Span4Mux_v
    port map (
            O => \N__68247\,
            I => \N__68226\
        );

    \I__15636\ : Span4Mux_h
    port map (
            O => \N__68244\,
            I => \N__68226\
        );

    \I__15635\ : Span4Mux_v
    port map (
            O => \N__68231\,
            I => \N__68223\
        );

    \I__15634\ : Odrv4
    port map (
            O => \N__68226\,
            I => \CONSTANT_ONE_NET\
        );

    \I__15633\ : Odrv4
    port map (
            O => \N__68223\,
            I => \CONSTANT_ONE_NET\
        );

    \I__15632\ : InMux
    port map (
            O => \N__68218\,
            I => \N__68215\
        );

    \I__15631\ : LocalMux
    port map (
            O => \N__68215\,
            I => \N__68211\
        );

    \I__15630\ : InMux
    port map (
            O => \N__68214\,
            I => \N__68208\
        );

    \I__15629\ : Odrv4
    port map (
            O => \N__68211\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21\
        );

    \I__15628\ : LocalMux
    port map (
            O => \N__68208\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21\
        );

    \I__15627\ : CascadeMux
    port map (
            O => \N__68203\,
            I => \N__68200\
        );

    \I__15626\ : InMux
    port map (
            O => \N__68200\,
            I => \N__68197\
        );

    \I__15625\ : LocalMux
    port map (
            O => \N__68197\,
            I => \N__68194\
        );

    \I__15624\ : Span4Mux_v
    port map (
            O => \N__68194\,
            I => \N__68191\
        );

    \I__15623\ : Odrv4
    port map (
            O => \N__68191\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_13\
        );

    \I__15622\ : InMux
    port map (
            O => \N__68188\,
            I => \N__68184\
        );

    \I__15621\ : InMux
    port map (
            O => \N__68187\,
            I => \N__68181\
        );

    \I__15620\ : LocalMux
    port map (
            O => \N__68184\,
            I => \N__68174\
        );

    \I__15619\ : LocalMux
    port map (
            O => \N__68181\,
            I => \N__68174\
        );

    \I__15618\ : CascadeMux
    port map (
            O => \N__68180\,
            I => \N__68171\
        );

    \I__15617\ : CascadeMux
    port map (
            O => \N__68179\,
            I => \N__68168\
        );

    \I__15616\ : Span4Mux_v
    port map (
            O => \N__68174\,
            I => \N__68165\
        );

    \I__15615\ : InMux
    port map (
            O => \N__68171\,
            I => \N__68162\
        );

    \I__15614\ : InMux
    port map (
            O => \N__68168\,
            I => \N__68159\
        );

    \I__15613\ : Span4Mux_v
    port map (
            O => \N__68165\,
            I => \N__68156\
        );

    \I__15612\ : LocalMux
    port map (
            O => \N__68162\,
            I => \N__68151\
        );

    \I__15611\ : LocalMux
    port map (
            O => \N__68159\,
            I => \N__68151\
        );

    \I__15610\ : Odrv4
    port map (
            O => \N__68156\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14\
        );

    \I__15609\ : Odrv12
    port map (
            O => \N__68151\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14\
        );

    \I__15608\ : InMux
    port map (
            O => \N__68146\,
            I => \bfn_24_18_0_\
        );

    \I__15607\ : CascadeMux
    port map (
            O => \N__68143\,
            I => \N__68140\
        );

    \I__15606\ : InMux
    port map (
            O => \N__68140\,
            I => \N__68137\
        );

    \I__15605\ : LocalMux
    port map (
            O => \N__68137\,
            I => \N__68133\
        );

    \I__15604\ : InMux
    port map (
            O => \N__68136\,
            I => \N__68130\
        );

    \I__15603\ : Odrv4
    port map (
            O => \N__68133\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22\
        );

    \I__15602\ : LocalMux
    port map (
            O => \N__68130\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22\
        );

    \I__15601\ : CascadeMux
    port map (
            O => \N__68125\,
            I => \N__68122\
        );

    \I__15600\ : InMux
    port map (
            O => \N__68122\,
            I => \N__68119\
        );

    \I__15599\ : LocalMux
    port map (
            O => \N__68119\,
            I => \N__68116\
        );

    \I__15598\ : Span4Mux_h
    port map (
            O => \N__68116\,
            I => \N__68113\
        );

    \I__15597\ : Span4Mux_v
    port map (
            O => \N__68113\,
            I => \N__68110\
        );

    \I__15596\ : Odrv4
    port map (
            O => \N__68110\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_14\
        );

    \I__15595\ : InMux
    port map (
            O => \N__68107\,
            I => \N__68101\
        );

    \I__15594\ : InMux
    port map (
            O => \N__68106\,
            I => \N__68101\
        );

    \I__15593\ : LocalMux
    port map (
            O => \N__68101\,
            I => \N__68096\
        );

    \I__15592\ : InMux
    port map (
            O => \N__68100\,
            I => \N__68091\
        );

    \I__15591\ : InMux
    port map (
            O => \N__68099\,
            I => \N__68091\
        );

    \I__15590\ : Sp12to4
    port map (
            O => \N__68096\,
            I => \N__68086\
        );

    \I__15589\ : LocalMux
    port map (
            O => \N__68091\,
            I => \N__68086\
        );

    \I__15588\ : Odrv12
    port map (
            O => \N__68086\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_15\
        );

    \I__15587\ : InMux
    port map (
            O => \N__68083\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15581\
        );

    \I__15586\ : InMux
    port map (
            O => \N__68080\,
            I => \N__68077\
        );

    \I__15585\ : LocalMux
    port map (
            O => \N__68077\,
            I => \N__68073\
        );

    \I__15584\ : InMux
    port map (
            O => \N__68076\,
            I => \N__68070\
        );

    \I__15583\ : Odrv4
    port map (
            O => \N__68073\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23\
        );

    \I__15582\ : LocalMux
    port map (
            O => \N__68070\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23\
        );

    \I__15581\ : CascadeMux
    port map (
            O => \N__68065\,
            I => \N__68062\
        );

    \I__15580\ : InMux
    port map (
            O => \N__68062\,
            I => \N__68059\
        );

    \I__15579\ : LocalMux
    port map (
            O => \N__68059\,
            I => \N__68056\
        );

    \I__15578\ : Span4Mux_v
    port map (
            O => \N__68056\,
            I => \N__68053\
        );

    \I__15577\ : Odrv4
    port map (
            O => \N__68053\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_15\
        );

    \I__15576\ : InMux
    port map (
            O => \N__68050\,
            I => \N__68042\
        );

    \I__15575\ : InMux
    port map (
            O => \N__68049\,
            I => \N__68042\
        );

    \I__15574\ : InMux
    port map (
            O => \N__68048\,
            I => \N__68037\
        );

    \I__15573\ : InMux
    port map (
            O => \N__68047\,
            I => \N__68037\
        );

    \I__15572\ : LocalMux
    port map (
            O => \N__68042\,
            I => \N__68034\
        );

    \I__15571\ : LocalMux
    port map (
            O => \N__68037\,
            I => \N__68031\
        );

    \I__15570\ : Sp12to4
    port map (
            O => \N__68034\,
            I => \N__68028\
        );

    \I__15569\ : Span4Mux_v
    port map (
            O => \N__68031\,
            I => \N__68025\
        );

    \I__15568\ : Odrv12
    port map (
            O => \N__68028\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16\
        );

    \I__15567\ : Odrv4
    port map (
            O => \N__68025\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16\
        );

    \I__15566\ : InMux
    port map (
            O => \N__68020\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15582\
        );

    \I__15565\ : InMux
    port map (
            O => \N__68017\,
            I => \N__68014\
        );

    \I__15564\ : LocalMux
    port map (
            O => \N__68014\,
            I => \N__68010\
        );

    \I__15563\ : InMux
    port map (
            O => \N__68013\,
            I => \N__68007\
        );

    \I__15562\ : Span4Mux_v
    port map (
            O => \N__68010\,
            I => \N__68004\
        );

    \I__15561\ : LocalMux
    port map (
            O => \N__68007\,
            I => \N__68001\
        );

    \I__15560\ : Odrv4
    port map (
            O => \N__68004\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24\
        );

    \I__15559\ : Odrv4
    port map (
            O => \N__68001\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24\
        );

    \I__15558\ : CascadeMux
    port map (
            O => \N__67996\,
            I => \N__67993\
        );

    \I__15557\ : InMux
    port map (
            O => \N__67993\,
            I => \N__67990\
        );

    \I__15556\ : LocalMux
    port map (
            O => \N__67990\,
            I => \N__67987\
        );

    \I__15555\ : Span4Mux_v
    port map (
            O => \N__67987\,
            I => \N__67984\
        );

    \I__15554\ : Span4Mux_h
    port map (
            O => \N__67984\,
            I => \N__67981\
        );

    \I__15553\ : Odrv4
    port map (
            O => \N__67981\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_16\
        );

    \I__15552\ : InMux
    port map (
            O => \N__67978\,
            I => \N__67974\
        );

    \I__15551\ : InMux
    port map (
            O => \N__67977\,
            I => \N__67971\
        );

    \I__15550\ : LocalMux
    port map (
            O => \N__67974\,
            I => \N__67965\
        );

    \I__15549\ : LocalMux
    port map (
            O => \N__67971\,
            I => \N__67965\
        );

    \I__15548\ : InMux
    port map (
            O => \N__67970\,
            I => \N__67961\
        );

    \I__15547\ : Span4Mux_h
    port map (
            O => \N__67965\,
            I => \N__67958\
        );

    \I__15546\ : InMux
    port map (
            O => \N__67964\,
            I => \N__67955\
        );

    \I__15545\ : LocalMux
    port map (
            O => \N__67961\,
            I => \N__67952\
        );

    \I__15544\ : Span4Mux_v
    port map (
            O => \N__67958\,
            I => \N__67949\
        );

    \I__15543\ : LocalMux
    port map (
            O => \N__67955\,
            I => \N__67946\
        );

    \I__15542\ : Span4Mux_v
    port map (
            O => \N__67952\,
            I => \N__67943\
        );

    \I__15541\ : Odrv4
    port map (
            O => \N__67949\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17\
        );

    \I__15540\ : Odrv12
    port map (
            O => \N__67946\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17\
        );

    \I__15539\ : Odrv4
    port map (
            O => \N__67943\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17\
        );

    \I__15538\ : InMux
    port map (
            O => \N__67936\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15583\
        );

    \I__15537\ : InMux
    port map (
            O => \N__67933\,
            I => \N__67930\
        );

    \I__15536\ : LocalMux
    port map (
            O => \N__67930\,
            I => \N__67926\
        );

    \I__15535\ : InMux
    port map (
            O => \N__67929\,
            I => \N__67923\
        );

    \I__15534\ : Span4Mux_v
    port map (
            O => \N__67926\,
            I => \N__67918\
        );

    \I__15533\ : LocalMux
    port map (
            O => \N__67923\,
            I => \N__67918\
        );

    \I__15532\ : Odrv4
    port map (
            O => \N__67918\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_25\
        );

    \I__15531\ : CascadeMux
    port map (
            O => \N__67915\,
            I => \N__67912\
        );

    \I__15530\ : InMux
    port map (
            O => \N__67912\,
            I => \N__67909\
        );

    \I__15529\ : LocalMux
    port map (
            O => \N__67909\,
            I => \N__67906\
        );

    \I__15528\ : Span4Mux_v
    port map (
            O => \N__67906\,
            I => \N__67903\
        );

    \I__15527\ : Odrv4
    port map (
            O => \N__67903\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_17\
        );

    \I__15526\ : CascadeMux
    port map (
            O => \N__67900\,
            I => \N__67895\
        );

    \I__15525\ : InMux
    port map (
            O => \N__67899\,
            I => \N__67892\
        );

    \I__15524\ : InMux
    port map (
            O => \N__67898\,
            I => \N__67889\
        );

    \I__15523\ : InMux
    port map (
            O => \N__67895\,
            I => \N__67886\
        );

    \I__15522\ : LocalMux
    port map (
            O => \N__67892\,
            I => \N__67880\
        );

    \I__15521\ : LocalMux
    port map (
            O => \N__67889\,
            I => \N__67880\
        );

    \I__15520\ : LocalMux
    port map (
            O => \N__67886\,
            I => \N__67877\
        );

    \I__15519\ : InMux
    port map (
            O => \N__67885\,
            I => \N__67874\
        );

    \I__15518\ : Span4Mux_h
    port map (
            O => \N__67880\,
            I => \N__67867\
        );

    \I__15517\ : Span4Mux_v
    port map (
            O => \N__67877\,
            I => \N__67867\
        );

    \I__15516\ : LocalMux
    port map (
            O => \N__67874\,
            I => \N__67867\
        );

    \I__15515\ : Odrv4
    port map (
            O => \N__67867\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_18\
        );

    \I__15514\ : InMux
    port map (
            O => \N__67864\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15584\
        );

    \I__15513\ : InMux
    port map (
            O => \N__67861\,
            I => \N__67858\
        );

    \I__15512\ : LocalMux
    port map (
            O => \N__67858\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20194\
        );

    \I__15511\ : InMux
    port map (
            O => \N__67855\,
            I => \N__67852\
        );

    \I__15510\ : LocalMux
    port map (
            O => \N__67852\,
            I => \N__67849\
        );

    \I__15509\ : Span4Mux_v
    port map (
            O => \N__67849\,
            I => \N__67846\
        );

    \I__15508\ : Odrv4
    port map (
            O => \N__67846\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_6\
        );

    \I__15507\ : InMux
    port map (
            O => \N__67843\,
            I => \N__67839\
        );

    \I__15506\ : CascadeMux
    port map (
            O => \N__67842\,
            I => \N__67836\
        );

    \I__15505\ : LocalMux
    port map (
            O => \N__67839\,
            I => \N__67833\
        );

    \I__15504\ : InMux
    port map (
            O => \N__67836\,
            I => \N__67830\
        );

    \I__15503\ : Odrv4
    port map (
            O => \N__67833\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14\
        );

    \I__15502\ : LocalMux
    port map (
            O => \N__67830\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14\
        );

    \I__15501\ : InMux
    port map (
            O => \N__67825\,
            I => \bfn_24_17_0_\
        );

    \I__15500\ : InMux
    port map (
            O => \N__67822\,
            I => \N__67819\
        );

    \I__15499\ : LocalMux
    port map (
            O => \N__67819\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20196\
        );

    \I__15498\ : CascadeMux
    port map (
            O => \N__67816\,
            I => \N__67813\
        );

    \I__15497\ : InMux
    port map (
            O => \N__67813\,
            I => \N__67810\
        );

    \I__15496\ : LocalMux
    port map (
            O => \N__67810\,
            I => \N__67806\
        );

    \I__15495\ : InMux
    port map (
            O => \N__67809\,
            I => \N__67803\
        );

    \I__15494\ : Odrv4
    port map (
            O => \N__67806\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15\
        );

    \I__15493\ : LocalMux
    port map (
            O => \N__67803\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15\
        );

    \I__15492\ : CascadeMux
    port map (
            O => \N__67798\,
            I => \N__67795\
        );

    \I__15491\ : InMux
    port map (
            O => \N__67795\,
            I => \N__67792\
        );

    \I__15490\ : LocalMux
    port map (
            O => \N__67792\,
            I => \N__67789\
        );

    \I__15489\ : Span4Mux_v
    port map (
            O => \N__67789\,
            I => \N__67786\
        );

    \I__15488\ : Odrv4
    port map (
            O => \N__67786\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_7\
        );

    \I__15487\ : InMux
    port map (
            O => \N__67783\,
            I => \N__67780\
        );

    \I__15486\ : LocalMux
    port map (
            O => \N__67780\,
            I => \N__67776\
        );

    \I__15485\ : InMux
    port map (
            O => \N__67779\,
            I => \N__67773\
        );

    \I__15484\ : Odrv4
    port map (
            O => \N__67776\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20198\
        );

    \I__15483\ : LocalMux
    port map (
            O => \N__67773\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20198\
        );

    \I__15482\ : InMux
    port map (
            O => \N__67768\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15574\
        );

    \I__15481\ : InMux
    port map (
            O => \N__67765\,
            I => \N__67762\
        );

    \I__15480\ : LocalMux
    port map (
            O => \N__67762\,
            I => \N__67759\
        );

    \I__15479\ : Span4Mux_v
    port map (
            O => \N__67759\,
            I => \N__67755\
        );

    \I__15478\ : InMux
    port map (
            O => \N__67758\,
            I => \N__67752\
        );

    \I__15477\ : Odrv4
    port map (
            O => \N__67755\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16\
        );

    \I__15476\ : LocalMux
    port map (
            O => \N__67752\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16\
        );

    \I__15475\ : CascadeMux
    port map (
            O => \N__67747\,
            I => \N__67744\
        );

    \I__15474\ : InMux
    port map (
            O => \N__67744\,
            I => \N__67741\
        );

    \I__15473\ : LocalMux
    port map (
            O => \N__67741\,
            I => \N__67738\
        );

    \I__15472\ : Span4Mux_v
    port map (
            O => \N__67738\,
            I => \N__67735\
        );

    \I__15471\ : Odrv4
    port map (
            O => \N__67735\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_8\
        );

    \I__15470\ : InMux
    port map (
            O => \N__67732\,
            I => \N__67729\
        );

    \I__15469\ : LocalMux
    port map (
            O => \N__67729\,
            I => \N__67725\
        );

    \I__15468\ : InMux
    port map (
            O => \N__67728\,
            I => \N__67722\
        );

    \I__15467\ : Odrv4
    port map (
            O => \N__67725\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9\
        );

    \I__15466\ : LocalMux
    port map (
            O => \N__67722\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9\
        );

    \I__15465\ : InMux
    port map (
            O => \N__67717\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15575\
        );

    \I__15464\ : InMux
    port map (
            O => \N__67714\,
            I => \N__67711\
        );

    \I__15463\ : LocalMux
    port map (
            O => \N__67711\,
            I => \N__67708\
        );

    \I__15462\ : Span4Mux_v
    port map (
            O => \N__67708\,
            I => \N__67705\
        );

    \I__15461\ : Odrv4
    port map (
            O => \N__67705\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_9\
        );

    \I__15460\ : InMux
    port map (
            O => \N__67702\,
            I => \N__67699\
        );

    \I__15459\ : LocalMux
    port map (
            O => \N__67699\,
            I => \N__67696\
        );

    \I__15458\ : Span4Mux_v
    port map (
            O => \N__67696\,
            I => \N__67692\
        );

    \I__15457\ : CascadeMux
    port map (
            O => \N__67695\,
            I => \N__67689\
        );

    \I__15456\ : Sp12to4
    port map (
            O => \N__67692\,
            I => \N__67686\
        );

    \I__15455\ : InMux
    port map (
            O => \N__67689\,
            I => \N__67683\
        );

    \I__15454\ : Odrv12
    port map (
            O => \N__67686\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17\
        );

    \I__15453\ : LocalMux
    port map (
            O => \N__67683\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17\
        );

    \I__15452\ : InMux
    port map (
            O => \N__67678\,
            I => \N__67674\
        );

    \I__15451\ : InMux
    port map (
            O => \N__67677\,
            I => \N__67670\
        );

    \I__15450\ : LocalMux
    port map (
            O => \N__67674\,
            I => \N__67667\
        );

    \I__15449\ : InMux
    port map (
            O => \N__67673\,
            I => \N__67664\
        );

    \I__15448\ : LocalMux
    port map (
            O => \N__67670\,
            I => \N__67661\
        );

    \I__15447\ : Odrv4
    port map (
            O => \N__67667\,
            I => \foc.preSatVoltage_10_adj_2311\
        );

    \I__15446\ : LocalMux
    port map (
            O => \N__67664\,
            I => \foc.preSatVoltage_10_adj_2311\
        );

    \I__15445\ : Odrv4
    port map (
            O => \N__67661\,
            I => \foc.preSatVoltage_10_adj_2311\
        );

    \I__15444\ : InMux
    port map (
            O => \N__67654\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15576\
        );

    \I__15443\ : InMux
    port map (
            O => \N__67651\,
            I => \N__67647\
        );

    \I__15442\ : InMux
    port map (
            O => \N__67650\,
            I => \N__67644\
        );

    \I__15441\ : LocalMux
    port map (
            O => \N__67647\,
            I => \N__67641\
        );

    \I__15440\ : LocalMux
    port map (
            O => \N__67644\,
            I => \N__67638\
        );

    \I__15439\ : Odrv12
    port map (
            O => \N__67641\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18\
        );

    \I__15438\ : Odrv4
    port map (
            O => \N__67638\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18\
        );

    \I__15437\ : CascadeMux
    port map (
            O => \N__67633\,
            I => \N__67630\
        );

    \I__15436\ : InMux
    port map (
            O => \N__67630\,
            I => \N__67627\
        );

    \I__15435\ : LocalMux
    port map (
            O => \N__67627\,
            I => \N__67624\
        );

    \I__15434\ : Span4Mux_v
    port map (
            O => \N__67624\,
            I => \N__67621\
        );

    \I__15433\ : Odrv4
    port map (
            O => \N__67621\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_10\
        );

    \I__15432\ : InMux
    port map (
            O => \N__67618\,
            I => \N__67612\
        );

    \I__15431\ : InMux
    port map (
            O => \N__67617\,
            I => \N__67612\
        );

    \I__15430\ : LocalMux
    port map (
            O => \N__67612\,
            I => \N__67607\
        );

    \I__15429\ : InMux
    port map (
            O => \N__67611\,
            I => \N__67604\
        );

    \I__15428\ : InMux
    port map (
            O => \N__67610\,
            I => \N__67601\
        );

    \I__15427\ : Span4Mux_h
    port map (
            O => \N__67607\,
            I => \N__67596\
        );

    \I__15426\ : LocalMux
    port map (
            O => \N__67604\,
            I => \N__67596\
        );

    \I__15425\ : LocalMux
    port map (
            O => \N__67601\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11\
        );

    \I__15424\ : Odrv4
    port map (
            O => \N__67596\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11\
        );

    \I__15423\ : InMux
    port map (
            O => \N__67591\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15577\
        );

    \I__15422\ : CascadeMux
    port map (
            O => \N__67588\,
            I => \N__67585\
        );

    \I__15421\ : InMux
    port map (
            O => \N__67585\,
            I => \N__67582\
        );

    \I__15420\ : LocalMux
    port map (
            O => \N__67582\,
            I => \N__67578\
        );

    \I__15419\ : InMux
    port map (
            O => \N__67581\,
            I => \N__67575\
        );

    \I__15418\ : Odrv4
    port map (
            O => \N__67578\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19\
        );

    \I__15417\ : LocalMux
    port map (
            O => \N__67575\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19\
        );

    \I__15416\ : CascadeMux
    port map (
            O => \N__67570\,
            I => \N__67567\
        );

    \I__15415\ : InMux
    port map (
            O => \N__67567\,
            I => \N__67564\
        );

    \I__15414\ : LocalMux
    port map (
            O => \N__67564\,
            I => \N__67561\
        );

    \I__15413\ : Span4Mux_v
    port map (
            O => \N__67561\,
            I => \N__67558\
        );

    \I__15412\ : Odrv4
    port map (
            O => \N__67558\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_11\
        );

    \I__15411\ : InMux
    port map (
            O => \N__67555\,
            I => \N__67549\
        );

    \I__15410\ : InMux
    port map (
            O => \N__67554\,
            I => \N__67549\
        );

    \I__15409\ : LocalMux
    port map (
            O => \N__67549\,
            I => \N__67544\
        );

    \I__15408\ : InMux
    port map (
            O => \N__67548\,
            I => \N__67541\
        );

    \I__15407\ : InMux
    port map (
            O => \N__67547\,
            I => \N__67538\
        );

    \I__15406\ : Span4Mux_v
    port map (
            O => \N__67544\,
            I => \N__67535\
        );

    \I__15405\ : LocalMux
    port map (
            O => \N__67541\,
            I => \N__67530\
        );

    \I__15404\ : LocalMux
    port map (
            O => \N__67538\,
            I => \N__67530\
        );

    \I__15403\ : Odrv4
    port map (
            O => \N__67535\,
            I => \foc.preSatVoltage_12_adj_2330\
        );

    \I__15402\ : Odrv4
    port map (
            O => \N__67530\,
            I => \foc.preSatVoltage_12_adj_2330\
        );

    \I__15401\ : InMux
    port map (
            O => \N__67525\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15578\
        );

    \I__15400\ : InMux
    port map (
            O => \N__67522\,
            I => \N__67519\
        );

    \I__15399\ : LocalMux
    port map (
            O => \N__67519\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19455\
        );

    \I__15398\ : InMux
    port map (
            O => \N__67516\,
            I => \N__67513\
        );

    \I__15397\ : LocalMux
    port map (
            O => \N__67513\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19690\
        );

    \I__15396\ : CascadeMux
    port map (
            O => \N__67510\,
            I => \N__67507\
        );

    \I__15395\ : InMux
    port map (
            O => \N__67507\,
            I => \N__67504\
        );

    \I__15394\ : LocalMux
    port map (
            O => \N__67504\,
            I => \N__67500\
        );

    \I__15393\ : InMux
    port map (
            O => \N__67503\,
            I => \N__67497\
        );

    \I__15392\ : Odrv4
    port map (
            O => \N__67500\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0\
        );

    \I__15391\ : LocalMux
    port map (
            O => \N__67497\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0\
        );

    \I__15390\ : InMux
    port map (
            O => \N__67492\,
            I => \N__67489\
        );

    \I__15389\ : LocalMux
    port map (
            O => \N__67489\,
            I => \N__67486\
        );

    \I__15388\ : Span12Mux_h
    port map (
            O => \N__67486\,
            I => \N__67482\
        );

    \I__15387\ : InMux
    port map (
            O => \N__67485\,
            I => \N__67479\
        );

    \I__15386\ : Odrv12
    port map (
            O => \N__67482\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8\
        );

    \I__15385\ : LocalMux
    port map (
            O => \N__67479\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8\
        );

    \I__15384\ : CascadeMux
    port map (
            O => \N__67474\,
            I => \N__67471\
        );

    \I__15383\ : InMux
    port map (
            O => \N__67471\,
            I => \N__67468\
        );

    \I__15382\ : LocalMux
    port map (
            O => \N__67468\,
            I => \N__67452\
        );

    \I__15381\ : CascadeMux
    port map (
            O => \N__67467\,
            I => \N__67449\
        );

    \I__15380\ : CascadeMux
    port map (
            O => \N__67466\,
            I => \N__67446\
        );

    \I__15379\ : CascadeMux
    port map (
            O => \N__67465\,
            I => \N__67443\
        );

    \I__15378\ : CascadeMux
    port map (
            O => \N__67464\,
            I => \N__67439\
        );

    \I__15377\ : CascadeMux
    port map (
            O => \N__67463\,
            I => \N__67436\
        );

    \I__15376\ : CascadeMux
    port map (
            O => \N__67462\,
            I => \N__67433\
        );

    \I__15375\ : CascadeMux
    port map (
            O => \N__67461\,
            I => \N__67430\
        );

    \I__15374\ : CascadeMux
    port map (
            O => \N__67460\,
            I => \N__67427\
        );

    \I__15373\ : CascadeMux
    port map (
            O => \N__67459\,
            I => \N__67422\
        );

    \I__15372\ : CascadeMux
    port map (
            O => \N__67458\,
            I => \N__67418\
        );

    \I__15371\ : CascadeMux
    port map (
            O => \N__67457\,
            I => \N__67414\
        );

    \I__15370\ : CascadeMux
    port map (
            O => \N__67456\,
            I => \N__67410\
        );

    \I__15369\ : CascadeMux
    port map (
            O => \N__67455\,
            I => \N__67406\
        );

    \I__15368\ : Span4Mux_v
    port map (
            O => \N__67452\,
            I => \N__67401\
        );

    \I__15367\ : InMux
    port map (
            O => \N__67449\,
            I => \N__67398\
        );

    \I__15366\ : InMux
    port map (
            O => \N__67446\,
            I => \N__67392\
        );

    \I__15365\ : InMux
    port map (
            O => \N__67443\,
            I => \N__67389\
        );

    \I__15364\ : CascadeMux
    port map (
            O => \N__67442\,
            I => \N__67386\
        );

    \I__15363\ : InMux
    port map (
            O => \N__67439\,
            I => \N__67381\
        );

    \I__15362\ : InMux
    port map (
            O => \N__67436\,
            I => \N__67381\
        );

    \I__15361\ : InMux
    port map (
            O => \N__67433\,
            I => \N__67372\
        );

    \I__15360\ : InMux
    port map (
            O => \N__67430\,
            I => \N__67372\
        );

    \I__15359\ : InMux
    port map (
            O => \N__67427\,
            I => \N__67372\
        );

    \I__15358\ : InMux
    port map (
            O => \N__67426\,
            I => \N__67372\
        );

    \I__15357\ : InMux
    port map (
            O => \N__67425\,
            I => \N__67355\
        );

    \I__15356\ : InMux
    port map (
            O => \N__67422\,
            I => \N__67355\
        );

    \I__15355\ : InMux
    port map (
            O => \N__67421\,
            I => \N__67355\
        );

    \I__15354\ : InMux
    port map (
            O => \N__67418\,
            I => \N__67355\
        );

    \I__15353\ : InMux
    port map (
            O => \N__67417\,
            I => \N__67355\
        );

    \I__15352\ : InMux
    port map (
            O => \N__67414\,
            I => \N__67355\
        );

    \I__15351\ : InMux
    port map (
            O => \N__67413\,
            I => \N__67355\
        );

    \I__15350\ : InMux
    port map (
            O => \N__67410\,
            I => \N__67355\
        );

    \I__15349\ : CascadeMux
    port map (
            O => \N__67409\,
            I => \N__67352\
        );

    \I__15348\ : InMux
    port map (
            O => \N__67406\,
            I => \N__67348\
        );

    \I__15347\ : CascadeMux
    port map (
            O => \N__67405\,
            I => \N__67345\
        );

    \I__15346\ : CascadeMux
    port map (
            O => \N__67404\,
            I => \N__67342\
        );

    \I__15345\ : Span4Mux_h
    port map (
            O => \N__67401\,
            I => \N__67337\
        );

    \I__15344\ : LocalMux
    port map (
            O => \N__67398\,
            I => \N__67337\
        );

    \I__15343\ : CascadeMux
    port map (
            O => \N__67397\,
            I => \N__67334\
        );

    \I__15342\ : CascadeMux
    port map (
            O => \N__67396\,
            I => \N__67331\
        );

    \I__15341\ : CascadeMux
    port map (
            O => \N__67395\,
            I => \N__67328\
        );

    \I__15340\ : LocalMux
    port map (
            O => \N__67392\,
            I => \N__67323\
        );

    \I__15339\ : LocalMux
    port map (
            O => \N__67389\,
            I => \N__67323\
        );

    \I__15338\ : InMux
    port map (
            O => \N__67386\,
            I => \N__67320\
        );

    \I__15337\ : LocalMux
    port map (
            O => \N__67381\,
            I => \N__67315\
        );

    \I__15336\ : LocalMux
    port map (
            O => \N__67372\,
            I => \N__67315\
        );

    \I__15335\ : LocalMux
    port map (
            O => \N__67355\,
            I => \N__67312\
        );

    \I__15334\ : InMux
    port map (
            O => \N__67352\,
            I => \N__67309\
        );

    \I__15333\ : CascadeMux
    port map (
            O => \N__67351\,
            I => \N__67306\
        );

    \I__15332\ : LocalMux
    port map (
            O => \N__67348\,
            I => \N__67303\
        );

    \I__15331\ : InMux
    port map (
            O => \N__67345\,
            I => \N__67300\
        );

    \I__15330\ : InMux
    port map (
            O => \N__67342\,
            I => \N__67297\
        );

    \I__15329\ : Span4Mux_v
    port map (
            O => \N__67337\,
            I => \N__67293\
        );

    \I__15328\ : InMux
    port map (
            O => \N__67334\,
            I => \N__67290\
        );

    \I__15327\ : InMux
    port map (
            O => \N__67331\,
            I => \N__67287\
        );

    \I__15326\ : InMux
    port map (
            O => \N__67328\,
            I => \N__67284\
        );

    \I__15325\ : Span4Mux_v
    port map (
            O => \N__67323\,
            I => \N__67279\
        );

    \I__15324\ : LocalMux
    port map (
            O => \N__67320\,
            I => \N__67279\
        );

    \I__15323\ : Span4Mux_v
    port map (
            O => \N__67315\,
            I => \N__67272\
        );

    \I__15322\ : Span4Mux_v
    port map (
            O => \N__67312\,
            I => \N__67272\
        );

    \I__15321\ : LocalMux
    port map (
            O => \N__67309\,
            I => \N__67272\
        );

    \I__15320\ : InMux
    port map (
            O => \N__67306\,
            I => \N__67269\
        );

    \I__15319\ : Span4Mux_v
    port map (
            O => \N__67303\,
            I => \N__67262\
        );

    \I__15318\ : LocalMux
    port map (
            O => \N__67300\,
            I => \N__67262\
        );

    \I__15317\ : LocalMux
    port map (
            O => \N__67297\,
            I => \N__67262\
        );

    \I__15316\ : CascadeMux
    port map (
            O => \N__67296\,
            I => \N__67259\
        );

    \I__15315\ : Span4Mux_h
    port map (
            O => \N__67293\,
            I => \N__67254\
        );

    \I__15314\ : LocalMux
    port map (
            O => \N__67290\,
            I => \N__67254\
        );

    \I__15313\ : LocalMux
    port map (
            O => \N__67287\,
            I => \N__67243\
        );

    \I__15312\ : LocalMux
    port map (
            O => \N__67284\,
            I => \N__67243\
        );

    \I__15311\ : Span4Mux_h
    port map (
            O => \N__67279\,
            I => \N__67243\
        );

    \I__15310\ : Span4Mux_h
    port map (
            O => \N__67272\,
            I => \N__67243\
        );

    \I__15309\ : LocalMux
    port map (
            O => \N__67269\,
            I => \N__67243\
        );

    \I__15308\ : Span4Mux_v
    port map (
            O => \N__67262\,
            I => \N__67240\
        );

    \I__15307\ : InMux
    port map (
            O => \N__67259\,
            I => \N__67237\
        );

    \I__15306\ : Span4Mux_v
    port map (
            O => \N__67254\,
            I => \N__67234\
        );

    \I__15305\ : Span4Mux_v
    port map (
            O => \N__67243\,
            I => \N__67227\
        );

    \I__15304\ : Span4Mux_v
    port map (
            O => \N__67240\,
            I => \N__67227\
        );

    \I__15303\ : LocalMux
    port map (
            O => \N__67237\,
            I => \N__67227\
        );

    \I__15302\ : Span4Mux_v
    port map (
            O => \N__67234\,
            I => \N__67224\
        );

    \I__15301\ : Span4Mux_v
    port map (
            O => \N__67227\,
            I => \N__67221\
        );

    \I__15300\ : Odrv4
    port map (
            O => \N__67224\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0\
        );

    \I__15299\ : Odrv4
    port map (
            O => \N__67221\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0\
        );

    \I__15298\ : InMux
    port map (
            O => \N__67216\,
            I => \N__67213\
        );

    \I__15297\ : LocalMux
    port map (
            O => \N__67213\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20184\
        );

    \I__15296\ : InMux
    port map (
            O => \N__67210\,
            I => \N__67207\
        );

    \I__15295\ : LocalMux
    port map (
            O => \N__67207\,
            I => \N__67204\
        );

    \I__15294\ : Span4Mux_v
    port map (
            O => \N__67204\,
            I => \N__67200\
        );

    \I__15293\ : InMux
    port map (
            O => \N__67203\,
            I => \N__67197\
        );

    \I__15292\ : Odrv4
    port map (
            O => \N__67200\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9\
        );

    \I__15291\ : LocalMux
    port map (
            O => \N__67197\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9\
        );

    \I__15290\ : CascadeMux
    port map (
            O => \N__67192\,
            I => \N__67189\
        );

    \I__15289\ : InMux
    port map (
            O => \N__67189\,
            I => \N__67186\
        );

    \I__15288\ : LocalMux
    port map (
            O => \N__67186\,
            I => \N__67183\
        );

    \I__15287\ : Span4Mux_v
    port map (
            O => \N__67183\,
            I => \N__67180\
        );

    \I__15286\ : Odrv4
    port map (
            O => \N__67180\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_1\
        );

    \I__15285\ : InMux
    port map (
            O => \N__67177\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15568\
        );

    \I__15284\ : InMux
    port map (
            O => \N__67174\,
            I => \N__67171\
        );

    \I__15283\ : LocalMux
    port map (
            O => \N__67171\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20186\
        );

    \I__15282\ : InMux
    port map (
            O => \N__67168\,
            I => \N__67165\
        );

    \I__15281\ : LocalMux
    port map (
            O => \N__67165\,
            I => \N__67162\
        );

    \I__15280\ : Span4Mux_v
    port map (
            O => \N__67162\,
            I => \N__67158\
        );

    \I__15279\ : InMux
    port map (
            O => \N__67161\,
            I => \N__67155\
        );

    \I__15278\ : Odrv4
    port map (
            O => \N__67158\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10\
        );

    \I__15277\ : LocalMux
    port map (
            O => \N__67155\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10\
        );

    \I__15276\ : CascadeMux
    port map (
            O => \N__67150\,
            I => \N__67147\
        );

    \I__15275\ : InMux
    port map (
            O => \N__67147\,
            I => \N__67144\
        );

    \I__15274\ : LocalMux
    port map (
            O => \N__67144\,
            I => \N__67141\
        );

    \I__15273\ : Span4Mux_v
    port map (
            O => \N__67141\,
            I => \N__67138\
        );

    \I__15272\ : Odrv4
    port map (
            O => \N__67138\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_2\
        );

    \I__15271\ : InMux
    port map (
            O => \N__67135\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15569\
        );

    \I__15270\ : InMux
    port map (
            O => \N__67132\,
            I => \N__67129\
        );

    \I__15269\ : LocalMux
    port map (
            O => \N__67129\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20188\
        );

    \I__15268\ : CascadeMux
    port map (
            O => \N__67126\,
            I => \N__67123\
        );

    \I__15267\ : InMux
    port map (
            O => \N__67123\,
            I => \N__67120\
        );

    \I__15266\ : LocalMux
    port map (
            O => \N__67120\,
            I => \N__67117\
        );

    \I__15265\ : Span4Mux_v
    port map (
            O => \N__67117\,
            I => \N__67113\
        );

    \I__15264\ : InMux
    port map (
            O => \N__67116\,
            I => \N__67110\
        );

    \I__15263\ : Odrv4
    port map (
            O => \N__67113\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11\
        );

    \I__15262\ : LocalMux
    port map (
            O => \N__67110\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11\
        );

    \I__15261\ : CascadeMux
    port map (
            O => \N__67105\,
            I => \N__67102\
        );

    \I__15260\ : InMux
    port map (
            O => \N__67102\,
            I => \N__67099\
        );

    \I__15259\ : LocalMux
    port map (
            O => \N__67099\,
            I => \N__67096\
        );

    \I__15258\ : Span4Mux_v
    port map (
            O => \N__67096\,
            I => \N__67093\
        );

    \I__15257\ : Odrv4
    port map (
            O => \N__67093\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_3\
        );

    \I__15256\ : InMux
    port map (
            O => \N__67090\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15570\
        );

    \I__15255\ : InMux
    port map (
            O => \N__67087\,
            I => \N__67084\
        );

    \I__15254\ : LocalMux
    port map (
            O => \N__67084\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20190\
        );

    \I__15253\ : InMux
    port map (
            O => \N__67081\,
            I => \N__67078\
        );

    \I__15252\ : LocalMux
    port map (
            O => \N__67078\,
            I => \N__67074\
        );

    \I__15251\ : InMux
    port map (
            O => \N__67077\,
            I => \N__67071\
        );

    \I__15250\ : Odrv4
    port map (
            O => \N__67074\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12\
        );

    \I__15249\ : LocalMux
    port map (
            O => \N__67071\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12\
        );

    \I__15248\ : CascadeMux
    port map (
            O => \N__67066\,
            I => \N__67063\
        );

    \I__15247\ : InMux
    port map (
            O => \N__67063\,
            I => \N__67060\
        );

    \I__15246\ : LocalMux
    port map (
            O => \N__67060\,
            I => \N__67057\
        );

    \I__15245\ : Span4Mux_v
    port map (
            O => \N__67057\,
            I => \N__67054\
        );

    \I__15244\ : Odrv4
    port map (
            O => \N__67054\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_4\
        );

    \I__15243\ : InMux
    port map (
            O => \N__67051\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15571\
        );

    \I__15242\ : InMux
    port map (
            O => \N__67048\,
            I => \N__67045\
        );

    \I__15241\ : LocalMux
    port map (
            O => \N__67045\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20192\
        );

    \I__15240\ : InMux
    port map (
            O => \N__67042\,
            I => \N__67039\
        );

    \I__15239\ : LocalMux
    port map (
            O => \N__67039\,
            I => \N__67036\
        );

    \I__15238\ : Span4Mux_h
    port map (
            O => \N__67036\,
            I => \N__67033\
        );

    \I__15237\ : Span4Mux_v
    port map (
            O => \N__67033\,
            I => \N__67029\
        );

    \I__15236\ : InMux
    port map (
            O => \N__67032\,
            I => \N__67026\
        );

    \I__15235\ : Odrv4
    port map (
            O => \N__67029\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13\
        );

    \I__15234\ : LocalMux
    port map (
            O => \N__67026\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13\
        );

    \I__15233\ : CascadeMux
    port map (
            O => \N__67021\,
            I => \N__67018\
        );

    \I__15232\ : InMux
    port map (
            O => \N__67018\,
            I => \N__67015\
        );

    \I__15231\ : LocalMux
    port map (
            O => \N__67015\,
            I => \N__67012\
        );

    \I__15230\ : Span4Mux_v
    port map (
            O => \N__67012\,
            I => \N__67009\
        );

    \I__15229\ : Span4Mux_h
    port map (
            O => \N__67009\,
            I => \N__67006\
        );

    \I__15228\ : Odrv4
    port map (
            O => \N__67006\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_5\
        );

    \I__15227\ : InMux
    port map (
            O => \N__67003\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15572\
        );

    \I__15226\ : InMux
    port map (
            O => \N__67000\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18277\
        );

    \I__15225\ : InMux
    port map (
            O => \N__66997\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767\
        );

    \I__15224\ : CascadeMux
    port map (
            O => \N__66994\,
            I => \N__66991\
        );

    \I__15223\ : InMux
    port map (
            O => \N__66991\,
            I => \N__66988\
        );

    \I__15222\ : LocalMux
    port map (
            O => \N__66988\,
            I => \N__66985\
        );

    \I__15221\ : Span4Mux_h
    port map (
            O => \N__66985\,
            I => \N__66982\
        );

    \I__15220\ : Span4Mux_v
    port map (
            O => \N__66982\,
            I => \N__66979\
        );

    \I__15219\ : Odrv4
    port map (
            O => \N__66979\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_CO\
        );

    \I__15218\ : InMux
    port map (
            O => \N__66976\,
            I => \N__66973\
        );

    \I__15217\ : LocalMux
    port map (
            O => \N__66973\,
            I => \N__66970\
        );

    \I__15216\ : Odrv4
    port map (
            O => \N__66970\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19926\
        );

    \I__15215\ : CascadeMux
    port map (
            O => \N__66967\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20112_cascade_\
        );

    \I__15214\ : InMux
    port map (
            O => \N__66964\,
            I => \N__66961\
        );

    \I__15213\ : LocalMux
    port map (
            O => \N__66961\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20098\
        );

    \I__15212\ : CascadeMux
    port map (
            O => \N__66958\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15171_cascade_\
        );

    \I__15211\ : CascadeMux
    port map (
            O => \N__66955\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15188_cascade_\
        );

    \I__15210\ : CascadeMux
    port map (
            O => \N__66952\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19688_cascade_\
        );

    \I__15209\ : InMux
    port map (
            O => \N__66949\,
            I => \N__66946\
        );

    \I__15208\ : LocalMux
    port map (
            O => \N__66946\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19424\
        );

    \I__15207\ : InMux
    port map (
            O => \N__66943\,
            I => \N__66940\
        );

    \I__15206\ : LocalMux
    port map (
            O => \N__66940\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n14851\
        );

    \I__15205\ : InMux
    port map (
            O => \N__66937\,
            I => \N__66934\
        );

    \I__15204\ : LocalMux
    port map (
            O => \N__66934\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n369\
        );

    \I__15203\ : CascadeMux
    port map (
            O => \N__66931\,
            I => \N__66917\
        );

    \I__15202\ : CascadeMux
    port map (
            O => \N__66930\,
            I => \N__66914\
        );

    \I__15201\ : CascadeMux
    port map (
            O => \N__66929\,
            I => \N__66910\
        );

    \I__15200\ : CascadeMux
    port map (
            O => \N__66928\,
            I => \N__66907\
        );

    \I__15199\ : CascadeMux
    port map (
            O => \N__66927\,
            I => \N__66904\
        );

    \I__15198\ : CascadeMux
    port map (
            O => \N__66926\,
            I => \N__66901\
        );

    \I__15197\ : CascadeMux
    port map (
            O => \N__66925\,
            I => \N__66898\
        );

    \I__15196\ : CascadeMux
    port map (
            O => \N__66924\,
            I => \N__66895\
        );

    \I__15195\ : CascadeMux
    port map (
            O => \N__66923\,
            I => \N__66892\
        );

    \I__15194\ : InMux
    port map (
            O => \N__66922\,
            I => \N__66885\
        );

    \I__15193\ : CascadeMux
    port map (
            O => \N__66921\,
            I => \N__66881\
        );

    \I__15192\ : CascadeMux
    port map (
            O => \N__66920\,
            I => \N__66877\
        );

    \I__15191\ : InMux
    port map (
            O => \N__66917\,
            I => \N__66870\
        );

    \I__15190\ : InMux
    port map (
            O => \N__66914\,
            I => \N__66870\
        );

    \I__15189\ : InMux
    port map (
            O => \N__66913\,
            I => \N__66861\
        );

    \I__15188\ : InMux
    port map (
            O => \N__66910\,
            I => \N__66861\
        );

    \I__15187\ : InMux
    port map (
            O => \N__66907\,
            I => \N__66861\
        );

    \I__15186\ : InMux
    port map (
            O => \N__66904\,
            I => \N__66861\
        );

    \I__15185\ : InMux
    port map (
            O => \N__66901\,
            I => \N__66852\
        );

    \I__15184\ : InMux
    port map (
            O => \N__66898\,
            I => \N__66852\
        );

    \I__15183\ : InMux
    port map (
            O => \N__66895\,
            I => \N__66852\
        );

    \I__15182\ : InMux
    port map (
            O => \N__66892\,
            I => \N__66852\
        );

    \I__15181\ : CascadeMux
    port map (
            O => \N__66891\,
            I => \N__66849\
        );

    \I__15180\ : CascadeMux
    port map (
            O => \N__66890\,
            I => \N__66846\
        );

    \I__15179\ : CascadeMux
    port map (
            O => \N__66889\,
            I => \N__66843\
        );

    \I__15178\ : CascadeMux
    port map (
            O => \N__66888\,
            I => \N__66840\
        );

    \I__15177\ : LocalMux
    port map (
            O => \N__66885\,
            I => \N__66837\
        );

    \I__15176\ : InMux
    port map (
            O => \N__66884\,
            I => \N__66834\
        );

    \I__15175\ : InMux
    port map (
            O => \N__66881\,
            I => \N__66831\
        );

    \I__15174\ : CascadeMux
    port map (
            O => \N__66880\,
            I => \N__66825\
        );

    \I__15173\ : InMux
    port map (
            O => \N__66877\,
            I => \N__66819\
        );

    \I__15172\ : CascadeMux
    port map (
            O => \N__66876\,
            I => \N__66816\
        );

    \I__15171\ : CascadeMux
    port map (
            O => \N__66875\,
            I => \N__66813\
        );

    \I__15170\ : LocalMux
    port map (
            O => \N__66870\,
            I => \N__66808\
        );

    \I__15169\ : LocalMux
    port map (
            O => \N__66861\,
            I => \N__66808\
        );

    \I__15168\ : LocalMux
    port map (
            O => \N__66852\,
            I => \N__66805\
        );

    \I__15167\ : InMux
    port map (
            O => \N__66849\,
            I => \N__66796\
        );

    \I__15166\ : InMux
    port map (
            O => \N__66846\,
            I => \N__66796\
        );

    \I__15165\ : InMux
    port map (
            O => \N__66843\,
            I => \N__66796\
        );

    \I__15164\ : InMux
    port map (
            O => \N__66840\,
            I => \N__66796\
        );

    \I__15163\ : Span4Mux_h
    port map (
            O => \N__66837\,
            I => \N__66789\
        );

    \I__15162\ : LocalMux
    port map (
            O => \N__66834\,
            I => \N__66789\
        );

    \I__15161\ : LocalMux
    port map (
            O => \N__66831\,
            I => \N__66789\
        );

    \I__15160\ : CascadeMux
    port map (
            O => \N__66830\,
            I => \N__66786\
        );

    \I__15159\ : CascadeMux
    port map (
            O => \N__66829\,
            I => \N__66783\
        );

    \I__15158\ : CascadeMux
    port map (
            O => \N__66828\,
            I => \N__66779\
        );

    \I__15157\ : InMux
    port map (
            O => \N__66825\,
            I => \N__66776\
        );

    \I__15156\ : CascadeMux
    port map (
            O => \N__66824\,
            I => \N__66773\
        );

    \I__15155\ : CascadeMux
    port map (
            O => \N__66823\,
            I => \N__66770\
        );

    \I__15154\ : InMux
    port map (
            O => \N__66822\,
            I => \N__66767\
        );

    \I__15153\ : LocalMux
    port map (
            O => \N__66819\,
            I => \N__66764\
        );

    \I__15152\ : InMux
    port map (
            O => \N__66816\,
            I => \N__66761\
        );

    \I__15151\ : InMux
    port map (
            O => \N__66813\,
            I => \N__66757\
        );

    \I__15150\ : Span4Mux_v
    port map (
            O => \N__66808\,
            I => \N__66750\
        );

    \I__15149\ : Span4Mux_h
    port map (
            O => \N__66805\,
            I => \N__66750\
        );

    \I__15148\ : LocalMux
    port map (
            O => \N__66796\,
            I => \N__66750\
        );

    \I__15147\ : Span4Mux_h
    port map (
            O => \N__66789\,
            I => \N__66747\
        );

    \I__15146\ : InMux
    port map (
            O => \N__66786\,
            I => \N__66744\
        );

    \I__15145\ : InMux
    port map (
            O => \N__66783\,
            I => \N__66741\
        );

    \I__15144\ : InMux
    port map (
            O => \N__66782\,
            I => \N__66738\
        );

    \I__15143\ : InMux
    port map (
            O => \N__66779\,
            I => \N__66735\
        );

    \I__15142\ : LocalMux
    port map (
            O => \N__66776\,
            I => \N__66732\
        );

    \I__15141\ : InMux
    port map (
            O => \N__66773\,
            I => \N__66729\
        );

    \I__15140\ : InMux
    port map (
            O => \N__66770\,
            I => \N__66726\
        );

    \I__15139\ : LocalMux
    port map (
            O => \N__66767\,
            I => \N__66723\
        );

    \I__15138\ : Span4Mux_h
    port map (
            O => \N__66764\,
            I => \N__66720\
        );

    \I__15137\ : LocalMux
    port map (
            O => \N__66761\,
            I => \N__66717\
        );

    \I__15136\ : InMux
    port map (
            O => \N__66760\,
            I => \N__66714\
        );

    \I__15135\ : LocalMux
    port map (
            O => \N__66757\,
            I => \N__66711\
        );

    \I__15134\ : Span4Mux_v
    port map (
            O => \N__66750\,
            I => \N__66708\
        );

    \I__15133\ : Sp12to4
    port map (
            O => \N__66747\,
            I => \N__66705\
        );

    \I__15132\ : LocalMux
    port map (
            O => \N__66744\,
            I => \N__66698\
        );

    \I__15131\ : LocalMux
    port map (
            O => \N__66741\,
            I => \N__66698\
        );

    \I__15130\ : LocalMux
    port map (
            O => \N__66738\,
            I => \N__66698\
        );

    \I__15129\ : LocalMux
    port map (
            O => \N__66735\,
            I => \N__66695\
        );

    \I__15128\ : Span4Mux_v
    port map (
            O => \N__66732\,
            I => \N__66688\
        );

    \I__15127\ : LocalMux
    port map (
            O => \N__66729\,
            I => \N__66688\
        );

    \I__15126\ : LocalMux
    port map (
            O => \N__66726\,
            I => \N__66688\
        );

    \I__15125\ : Span4Mux_v
    port map (
            O => \N__66723\,
            I => \N__66685\
        );

    \I__15124\ : Span4Mux_v
    port map (
            O => \N__66720\,
            I => \N__66676\
        );

    \I__15123\ : Span4Mux_v
    port map (
            O => \N__66717\,
            I => \N__66676\
        );

    \I__15122\ : LocalMux
    port map (
            O => \N__66714\,
            I => \N__66676\
        );

    \I__15121\ : Span4Mux_v
    port map (
            O => \N__66711\,
            I => \N__66676\
        );

    \I__15120\ : Span4Mux_h
    port map (
            O => \N__66708\,
            I => \N__66673\
        );

    \I__15119\ : Span12Mux_s7_v
    port map (
            O => \N__66705\,
            I => \N__66668\
        );

    \I__15118\ : Span12Mux_h
    port map (
            O => \N__66698\,
            I => \N__66668\
        );

    \I__15117\ : Span4Mux_v
    port map (
            O => \N__66695\,
            I => \N__66663\
        );

    \I__15116\ : Span4Mux_v
    port map (
            O => \N__66688\,
            I => \N__66663\
        );

    \I__15115\ : Span4Mux_h
    port map (
            O => \N__66685\,
            I => \N__66658\
        );

    \I__15114\ : Span4Mux_h
    port map (
            O => \N__66676\,
            I => \N__66658\
        );

    \I__15113\ : Odrv4
    port map (
            O => \N__66673\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n123\
        );

    \I__15112\ : Odrv12
    port map (
            O => \N__66668\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n123\
        );

    \I__15111\ : Odrv4
    port map (
            O => \N__66663\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n123\
        );

    \I__15110\ : Odrv4
    port map (
            O => \N__66658\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n123\
        );

    \I__15109\ : InMux
    port map (
            O => \N__66649\,
            I => \N__66646\
        );

    \I__15108\ : LocalMux
    port map (
            O => \N__66646\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n415\
        );

    \I__15107\ : InMux
    port map (
            O => \N__66643\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18270\
        );

    \I__15106\ : CascadeMux
    port map (
            O => \N__66640\,
            I => \N__66635\
        );

    \I__15105\ : CascadeMux
    port map (
            O => \N__66639\,
            I => \N__66632\
        );

    \I__15104\ : InMux
    port map (
            O => \N__66638\,
            I => \N__66626\
        );

    \I__15103\ : InMux
    port map (
            O => \N__66635\,
            I => \N__66622\
        );

    \I__15102\ : InMux
    port map (
            O => \N__66632\,
            I => \N__66619\
        );

    \I__15101\ : CascadeMux
    port map (
            O => \N__66631\,
            I => \N__66616\
        );

    \I__15100\ : CascadeMux
    port map (
            O => \N__66630\,
            I => \N__66613\
        );

    \I__15099\ : CascadeMux
    port map (
            O => \N__66629\,
            I => \N__66609\
        );

    \I__15098\ : LocalMux
    port map (
            O => \N__66626\,
            I => \N__66605\
        );

    \I__15097\ : CascadeMux
    port map (
            O => \N__66625\,
            I => \N__66601\
        );

    \I__15096\ : LocalMux
    port map (
            O => \N__66622\,
            I => \N__66595\
        );

    \I__15095\ : LocalMux
    port map (
            O => \N__66619\,
            I => \N__66592\
        );

    \I__15094\ : InMux
    port map (
            O => \N__66616\,
            I => \N__66589\
        );

    \I__15093\ : InMux
    port map (
            O => \N__66613\,
            I => \N__66586\
        );

    \I__15092\ : InMux
    port map (
            O => \N__66612\,
            I => \N__66583\
        );

    \I__15091\ : InMux
    port map (
            O => \N__66609\,
            I => \N__66580\
        );

    \I__15090\ : CascadeMux
    port map (
            O => \N__66608\,
            I => \N__66577\
        );

    \I__15089\ : Span4Mux_v
    port map (
            O => \N__66605\,
            I => \N__66571\
        );

    \I__15088\ : CascadeMux
    port map (
            O => \N__66604\,
            I => \N__66568\
        );

    \I__15087\ : InMux
    port map (
            O => \N__66601\,
            I => \N__66565\
        );

    \I__15086\ : CascadeMux
    port map (
            O => \N__66600\,
            I => \N__66562\
        );

    \I__15085\ : CascadeMux
    port map (
            O => \N__66599\,
            I => \N__66559\
        );

    \I__15084\ : InMux
    port map (
            O => \N__66598\,
            I => \N__66556\
        );

    \I__15083\ : Span4Mux_v
    port map (
            O => \N__66595\,
            I => \N__66549\
        );

    \I__15082\ : Span4Mux_v
    port map (
            O => \N__66592\,
            I => \N__66549\
        );

    \I__15081\ : LocalMux
    port map (
            O => \N__66589\,
            I => \N__66549\
        );

    \I__15080\ : LocalMux
    port map (
            O => \N__66586\,
            I => \N__66542\
        );

    \I__15079\ : LocalMux
    port map (
            O => \N__66583\,
            I => \N__66542\
        );

    \I__15078\ : LocalMux
    port map (
            O => \N__66580\,
            I => \N__66542\
        );

    \I__15077\ : InMux
    port map (
            O => \N__66577\,
            I => \N__66539\
        );

    \I__15076\ : CascadeMux
    port map (
            O => \N__66576\,
            I => \N__66535\
        );

    \I__15075\ : CascadeMux
    port map (
            O => \N__66575\,
            I => \N__66531\
        );

    \I__15074\ : CascadeMux
    port map (
            O => \N__66574\,
            I => \N__66528\
        );

    \I__15073\ : Span4Mux_h
    port map (
            O => \N__66571\,
            I => \N__66525\
        );

    \I__15072\ : InMux
    port map (
            O => \N__66568\,
            I => \N__66522\
        );

    \I__15071\ : LocalMux
    port map (
            O => \N__66565\,
            I => \N__66512\
        );

    \I__15070\ : InMux
    port map (
            O => \N__66562\,
            I => \N__66509\
        );

    \I__15069\ : InMux
    port map (
            O => \N__66559\,
            I => \N__66506\
        );

    \I__15068\ : LocalMux
    port map (
            O => \N__66556\,
            I => \N__66503\
        );

    \I__15067\ : Span4Mux_h
    port map (
            O => \N__66549\,
            I => \N__66496\
        );

    \I__15066\ : Span4Mux_v
    port map (
            O => \N__66542\,
            I => \N__66496\
        );

    \I__15065\ : LocalMux
    port map (
            O => \N__66539\,
            I => \N__66496\
        );

    \I__15064\ : InMux
    port map (
            O => \N__66538\,
            I => \N__66493\
        );

    \I__15063\ : InMux
    port map (
            O => \N__66535\,
            I => \N__66486\
        );

    \I__15062\ : InMux
    port map (
            O => \N__66534\,
            I => \N__66486\
        );

    \I__15061\ : InMux
    port map (
            O => \N__66531\,
            I => \N__66486\
        );

    \I__15060\ : InMux
    port map (
            O => \N__66528\,
            I => \N__66483\
        );

    \I__15059\ : Span4Mux_v
    port map (
            O => \N__66525\,
            I => \N__66478\
        );

    \I__15058\ : LocalMux
    port map (
            O => \N__66522\,
            I => \N__66478\
        );

    \I__15057\ : CascadeMux
    port map (
            O => \N__66521\,
            I => \N__66475\
        );

    \I__15056\ : CascadeMux
    port map (
            O => \N__66520\,
            I => \N__66472\
        );

    \I__15055\ : CascadeMux
    port map (
            O => \N__66519\,
            I => \N__66469\
        );

    \I__15054\ : CascadeMux
    port map (
            O => \N__66518\,
            I => \N__66465\
        );

    \I__15053\ : CascadeMux
    port map (
            O => \N__66517\,
            I => \N__66461\
        );

    \I__15052\ : CascadeMux
    port map (
            O => \N__66516\,
            I => \N__66458\
        );

    \I__15051\ : CascadeMux
    port map (
            O => \N__66515\,
            I => \N__66455\
        );

    \I__15050\ : Span4Mux_v
    port map (
            O => \N__66512\,
            I => \N__66448\
        );

    \I__15049\ : LocalMux
    port map (
            O => \N__66509\,
            I => \N__66448\
        );

    \I__15048\ : LocalMux
    port map (
            O => \N__66506\,
            I => \N__66448\
        );

    \I__15047\ : Sp12to4
    port map (
            O => \N__66503\,
            I => \N__66445\
        );

    \I__15046\ : Span4Mux_v
    port map (
            O => \N__66496\,
            I => \N__66442\
        );

    \I__15045\ : LocalMux
    port map (
            O => \N__66493\,
            I => \N__66435\
        );

    \I__15044\ : LocalMux
    port map (
            O => \N__66486\,
            I => \N__66435\
        );

    \I__15043\ : LocalMux
    port map (
            O => \N__66483\,
            I => \N__66435\
        );

    \I__15042\ : Span4Mux_v
    port map (
            O => \N__66478\,
            I => \N__66432\
        );

    \I__15041\ : InMux
    port map (
            O => \N__66475\,
            I => \N__66429\
        );

    \I__15040\ : InMux
    port map (
            O => \N__66472\,
            I => \N__66416\
        );

    \I__15039\ : InMux
    port map (
            O => \N__66469\,
            I => \N__66416\
        );

    \I__15038\ : InMux
    port map (
            O => \N__66468\,
            I => \N__66416\
        );

    \I__15037\ : InMux
    port map (
            O => \N__66465\,
            I => \N__66416\
        );

    \I__15036\ : InMux
    port map (
            O => \N__66464\,
            I => \N__66416\
        );

    \I__15035\ : InMux
    port map (
            O => \N__66461\,
            I => \N__66416\
        );

    \I__15034\ : InMux
    port map (
            O => \N__66458\,
            I => \N__66411\
        );

    \I__15033\ : InMux
    port map (
            O => \N__66455\,
            I => \N__66411\
        );

    \I__15032\ : Span4Mux_v
    port map (
            O => \N__66448\,
            I => \N__66408\
        );

    \I__15031\ : Span12Mux_s10_v
    port map (
            O => \N__66445\,
            I => \N__66393\
        );

    \I__15030\ : Sp12to4
    port map (
            O => \N__66442\,
            I => \N__66393\
        );

    \I__15029\ : Span12Mux_s10_v
    port map (
            O => \N__66435\,
            I => \N__66393\
        );

    \I__15028\ : Sp12to4
    port map (
            O => \N__66432\,
            I => \N__66393\
        );

    \I__15027\ : LocalMux
    port map (
            O => \N__66429\,
            I => \N__66393\
        );

    \I__15026\ : LocalMux
    port map (
            O => \N__66416\,
            I => \N__66393\
        );

    \I__15025\ : LocalMux
    port map (
            O => \N__66411\,
            I => \N__66393\
        );

    \I__15024\ : Odrv4
    port map (
            O => \N__66408\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n126\
        );

    \I__15023\ : Odrv12
    port map (
            O => \N__66393\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n126\
        );

    \I__15022\ : CascadeMux
    port map (
            O => \N__66388\,
            I => \N__66385\
        );

    \I__15021\ : InMux
    port map (
            O => \N__66385\,
            I => \N__66382\
        );

    \I__15020\ : LocalMux
    port map (
            O => \N__66382\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n418\
        );

    \I__15019\ : InMux
    port map (
            O => \N__66379\,
            I => \N__66376\
        );

    \I__15018\ : LocalMux
    port map (
            O => \N__66376\,
            I => \N__66373\
        );

    \I__15017\ : Odrv4
    port map (
            O => \N__66373\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n464\
        );

    \I__15016\ : InMux
    port map (
            O => \N__66370\,
            I => \bfn_23_28_0_\
        );

    \I__15015\ : InMux
    port map (
            O => \N__66367\,
            I => \N__66364\
        );

    \I__15014\ : LocalMux
    port map (
            O => \N__66364\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n467\
        );

    \I__15013\ : CascadeMux
    port map (
            O => \N__66361\,
            I => \N__66356\
        );

    \I__15012\ : CascadeMux
    port map (
            O => \N__66360\,
            I => \N__66353\
        );

    \I__15011\ : CascadeMux
    port map (
            O => \N__66359\,
            I => \N__66350\
        );

    \I__15010\ : InMux
    port map (
            O => \N__66356\,
            I => \N__66340\
        );

    \I__15009\ : InMux
    port map (
            O => \N__66353\,
            I => \N__66337\
        );

    \I__15008\ : InMux
    port map (
            O => \N__66350\,
            I => \N__66334\
        );

    \I__15007\ : CascadeMux
    port map (
            O => \N__66349\,
            I => \N__66331\
        );

    \I__15006\ : CascadeMux
    port map (
            O => \N__66348\,
            I => \N__66328\
        );

    \I__15005\ : CascadeMux
    port map (
            O => \N__66347\,
            I => \N__66324\
        );

    \I__15004\ : CascadeMux
    port map (
            O => \N__66346\,
            I => \N__66321\
        );

    \I__15003\ : CascadeMux
    port map (
            O => \N__66345\,
            I => \N__66318\
        );

    \I__15002\ : CascadeMux
    port map (
            O => \N__66344\,
            I => \N__66315\
        );

    \I__15001\ : CascadeMux
    port map (
            O => \N__66343\,
            I => \N__66312\
        );

    \I__15000\ : LocalMux
    port map (
            O => \N__66340\,
            I => \N__66307\
        );

    \I__14999\ : LocalMux
    port map (
            O => \N__66337\,
            I => \N__66307\
        );

    \I__14998\ : LocalMux
    port map (
            O => \N__66334\,
            I => \N__66304\
        );

    \I__14997\ : InMux
    port map (
            O => \N__66331\,
            I => \N__66301\
        );

    \I__14996\ : InMux
    port map (
            O => \N__66328\,
            I => \N__66298\
        );

    \I__14995\ : CascadeMux
    port map (
            O => \N__66327\,
            I => \N__66295\
        );

    \I__14994\ : InMux
    port map (
            O => \N__66324\,
            I => \N__66290\
        );

    \I__14993\ : InMux
    port map (
            O => \N__66321\,
            I => \N__66287\
        );

    \I__14992\ : InMux
    port map (
            O => \N__66318\,
            I => \N__66283\
        );

    \I__14991\ : InMux
    port map (
            O => \N__66315\,
            I => \N__66280\
        );

    \I__14990\ : InMux
    port map (
            O => \N__66312\,
            I => \N__66277\
        );

    \I__14989\ : Span4Mux_v
    port map (
            O => \N__66307\,
            I => \N__66268\
        );

    \I__14988\ : Span4Mux_v
    port map (
            O => \N__66304\,
            I => \N__66268\
        );

    \I__14987\ : LocalMux
    port map (
            O => \N__66301\,
            I => \N__66268\
        );

    \I__14986\ : LocalMux
    port map (
            O => \N__66298\,
            I => \N__66268\
        );

    \I__14985\ : InMux
    port map (
            O => \N__66295\,
            I => \N__66265\
        );

    \I__14984\ : CascadeMux
    port map (
            O => \N__66294\,
            I => \N__66262\
        );

    \I__14983\ : CascadeMux
    port map (
            O => \N__66293\,
            I => \N__66256\
        );

    \I__14982\ : LocalMux
    port map (
            O => \N__66290\,
            I => \N__66253\
        );

    \I__14981\ : LocalMux
    port map (
            O => \N__66287\,
            I => \N__66250\
        );

    \I__14980\ : CascadeMux
    port map (
            O => \N__66286\,
            I => \N__66247\
        );

    \I__14979\ : LocalMux
    port map (
            O => \N__66283\,
            I => \N__66244\
        );

    \I__14978\ : LocalMux
    port map (
            O => \N__66280\,
            I => \N__66235\
        );

    \I__14977\ : LocalMux
    port map (
            O => \N__66277\,
            I => \N__66235\
        );

    \I__14976\ : Span4Mux_h
    port map (
            O => \N__66268\,
            I => \N__66235\
        );

    \I__14975\ : LocalMux
    port map (
            O => \N__66265\,
            I => \N__66235\
        );

    \I__14974\ : InMux
    port map (
            O => \N__66262\,
            I => \N__66232\
        );

    \I__14973\ : CascadeMux
    port map (
            O => \N__66261\,
            I => \N__66229\
        );

    \I__14972\ : InMux
    port map (
            O => \N__66260\,
            I => \N__66226\
        );

    \I__14971\ : InMux
    port map (
            O => \N__66259\,
            I => \N__66221\
        );

    \I__14970\ : InMux
    port map (
            O => \N__66256\,
            I => \N__66221\
        );

    \I__14969\ : Span4Mux_v
    port map (
            O => \N__66253\,
            I => \N__66214\
        );

    \I__14968\ : Span4Mux_v
    port map (
            O => \N__66250\,
            I => \N__66211\
        );

    \I__14967\ : InMux
    port map (
            O => \N__66247\,
            I => \N__66208\
        );

    \I__14966\ : Span4Mux_h
    port map (
            O => \N__66244\,
            I => \N__66201\
        );

    \I__14965\ : Span4Mux_v
    port map (
            O => \N__66235\,
            I => \N__66201\
        );

    \I__14964\ : LocalMux
    port map (
            O => \N__66232\,
            I => \N__66201\
        );

    \I__14963\ : InMux
    port map (
            O => \N__66229\,
            I => \N__66198\
        );

    \I__14962\ : LocalMux
    port map (
            O => \N__66226\,
            I => \N__66193\
        );

    \I__14961\ : LocalMux
    port map (
            O => \N__66221\,
            I => \N__66193\
        );

    \I__14960\ : CascadeMux
    port map (
            O => \N__66220\,
            I => \N__66189\
        );

    \I__14959\ : CascadeMux
    port map (
            O => \N__66219\,
            I => \N__66185\
        );

    \I__14958\ : CascadeMux
    port map (
            O => \N__66218\,
            I => \N__66181\
        );

    \I__14957\ : CascadeMux
    port map (
            O => \N__66217\,
            I => \N__66177\
        );

    \I__14956\ : Span4Mux_h
    port map (
            O => \N__66214\,
            I => \N__66174\
        );

    \I__14955\ : Span4Mux_v
    port map (
            O => \N__66211\,
            I => \N__66169\
        );

    \I__14954\ : LocalMux
    port map (
            O => \N__66208\,
            I => \N__66169\
        );

    \I__14953\ : Span4Mux_v
    port map (
            O => \N__66201\,
            I => \N__66166\
        );

    \I__14952\ : LocalMux
    port map (
            O => \N__66198\,
            I => \N__66163\
        );

    \I__14951\ : Span4Mux_v
    port map (
            O => \N__66193\,
            I => \N__66160\
        );

    \I__14950\ : InMux
    port map (
            O => \N__66192\,
            I => \N__66143\
        );

    \I__14949\ : InMux
    port map (
            O => \N__66189\,
            I => \N__66143\
        );

    \I__14948\ : InMux
    port map (
            O => \N__66188\,
            I => \N__66143\
        );

    \I__14947\ : InMux
    port map (
            O => \N__66185\,
            I => \N__66143\
        );

    \I__14946\ : InMux
    port map (
            O => \N__66184\,
            I => \N__66143\
        );

    \I__14945\ : InMux
    port map (
            O => \N__66181\,
            I => \N__66143\
        );

    \I__14944\ : InMux
    port map (
            O => \N__66180\,
            I => \N__66143\
        );

    \I__14943\ : InMux
    port map (
            O => \N__66177\,
            I => \N__66143\
        );

    \I__14942\ : Span4Mux_v
    port map (
            O => \N__66174\,
            I => \N__66140\
        );

    \I__14941\ : Span4Mux_v
    port map (
            O => \N__66169\,
            I => \N__66137\
        );

    \I__14940\ : Span4Mux_h
    port map (
            O => \N__66166\,
            I => \N__66132\
        );

    \I__14939\ : Span4Mux_h
    port map (
            O => \N__66163\,
            I => \N__66132\
        );

    \I__14938\ : Sp12to4
    port map (
            O => \N__66160\,
            I => \N__66127\
        );

    \I__14937\ : LocalMux
    port map (
            O => \N__66143\,
            I => \N__66127\
        );

    \I__14936\ : Odrv4
    port map (
            O => \N__66140\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n129\
        );

    \I__14935\ : Odrv4
    port map (
            O => \N__66137\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n129\
        );

    \I__14934\ : Odrv4
    port map (
            O => \N__66132\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n129\
        );

    \I__14933\ : Odrv12
    port map (
            O => \N__66127\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n129\
        );

    \I__14932\ : InMux
    port map (
            O => \N__66118\,
            I => \N__66115\
        );

    \I__14931\ : LocalMux
    port map (
            O => \N__66115\,
            I => \N__66112\
        );

    \I__14930\ : Odrv4
    port map (
            O => \N__66112\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n513\
        );

    \I__14929\ : InMux
    port map (
            O => \N__66109\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18272\
        );

    \I__14928\ : InMux
    port map (
            O => \N__66106\,
            I => \N__66103\
        );

    \I__14927\ : LocalMux
    port map (
            O => \N__66103\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n516\
        );

    \I__14926\ : CascadeMux
    port map (
            O => \N__66100\,
            I => \N__66095\
        );

    \I__14925\ : CascadeMux
    port map (
            O => \N__66099\,
            I => \N__66087\
        );

    \I__14924\ : CascadeMux
    port map (
            O => \N__66098\,
            I => \N__66083\
        );

    \I__14923\ : InMux
    port map (
            O => \N__66095\,
            I => \N__66080\
        );

    \I__14922\ : CascadeMux
    port map (
            O => \N__66094\,
            I => \N__66077\
        );

    \I__14921\ : CascadeMux
    port map (
            O => \N__66093\,
            I => \N__66074\
        );

    \I__14920\ : CascadeMux
    port map (
            O => \N__66092\,
            I => \N__66071\
        );

    \I__14919\ : CascadeMux
    port map (
            O => \N__66091\,
            I => \N__66067\
        );

    \I__14918\ : CascadeMux
    port map (
            O => \N__66090\,
            I => \N__66064\
        );

    \I__14917\ : InMux
    port map (
            O => \N__66087\,
            I => \N__66060\
        );

    \I__14916\ : CascadeMux
    port map (
            O => \N__66086\,
            I => \N__66057\
        );

    \I__14915\ : InMux
    port map (
            O => \N__66083\,
            I => \N__66053\
        );

    \I__14914\ : LocalMux
    port map (
            O => \N__66080\,
            I => \N__66050\
        );

    \I__14913\ : InMux
    port map (
            O => \N__66077\,
            I => \N__66047\
        );

    \I__14912\ : InMux
    port map (
            O => \N__66074\,
            I => \N__66044\
        );

    \I__14911\ : InMux
    port map (
            O => \N__66071\,
            I => \N__66041\
        );

    \I__14910\ : CascadeMux
    port map (
            O => \N__66070\,
            I => \N__66037\
        );

    \I__14909\ : InMux
    port map (
            O => \N__66067\,
            I => \N__66033\
        );

    \I__14908\ : InMux
    port map (
            O => \N__66064\,
            I => \N__66025\
        );

    \I__14907\ : CascadeMux
    port map (
            O => \N__66063\,
            I => \N__66022\
        );

    \I__14906\ : LocalMux
    port map (
            O => \N__66060\,
            I => \N__66019\
        );

    \I__14905\ : InMux
    port map (
            O => \N__66057\,
            I => \N__66016\
        );

    \I__14904\ : InMux
    port map (
            O => \N__66056\,
            I => \N__66013\
        );

    \I__14903\ : LocalMux
    port map (
            O => \N__66053\,
            I => \N__66005\
        );

    \I__14902\ : Span4Mux_v
    port map (
            O => \N__66050\,
            I => \N__66005\
        );

    \I__14901\ : LocalMux
    port map (
            O => \N__66047\,
            I => \N__66005\
        );

    \I__14900\ : LocalMux
    port map (
            O => \N__66044\,
            I => \N__66002\
        );

    \I__14899\ : LocalMux
    port map (
            O => \N__66041\,
            I => \N__65999\
        );

    \I__14898\ : InMux
    port map (
            O => \N__66040\,
            I => \N__65996\
        );

    \I__14897\ : InMux
    port map (
            O => \N__66037\,
            I => \N__65993\
        );

    \I__14896\ : CascadeMux
    port map (
            O => \N__66036\,
            I => \N__65990\
        );

    \I__14895\ : LocalMux
    port map (
            O => \N__66033\,
            I => \N__65987\
        );

    \I__14894\ : CascadeMux
    port map (
            O => \N__66032\,
            I => \N__65984\
        );

    \I__14893\ : CascadeMux
    port map (
            O => \N__66031\,
            I => \N__65980\
        );

    \I__14892\ : CascadeMux
    port map (
            O => \N__66030\,
            I => \N__65976\
        );

    \I__14891\ : CascadeMux
    port map (
            O => \N__66029\,
            I => \N__65972\
        );

    \I__14890\ : CascadeMux
    port map (
            O => \N__66028\,
            I => \N__65969\
        );

    \I__14889\ : LocalMux
    port map (
            O => \N__66025\,
            I => \N__65966\
        );

    \I__14888\ : InMux
    port map (
            O => \N__66022\,
            I => \N__65963\
        );

    \I__14887\ : Span4Mux_h
    port map (
            O => \N__66019\,
            I => \N__65958\
        );

    \I__14886\ : LocalMux
    port map (
            O => \N__66016\,
            I => \N__65958\
        );

    \I__14885\ : LocalMux
    port map (
            O => \N__66013\,
            I => \N__65955\
        );

    \I__14884\ : CascadeMux
    port map (
            O => \N__66012\,
            I => \N__65952\
        );

    \I__14883\ : Span4Mux_h
    port map (
            O => \N__66005\,
            I => \N__65941\
        );

    \I__14882\ : Span4Mux_h
    port map (
            O => \N__66002\,
            I => \N__65941\
        );

    \I__14881\ : Span4Mux_h
    port map (
            O => \N__65999\,
            I => \N__65941\
        );

    \I__14880\ : LocalMux
    port map (
            O => \N__65996\,
            I => \N__65941\
        );

    \I__14879\ : LocalMux
    port map (
            O => \N__65993\,
            I => \N__65941\
        );

    \I__14878\ : InMux
    port map (
            O => \N__65990\,
            I => \N__65938\
        );

    \I__14877\ : Span4Mux_v
    port map (
            O => \N__65987\,
            I => \N__65935\
        );

    \I__14876\ : InMux
    port map (
            O => \N__65984\,
            I => \N__65928\
        );

    \I__14875\ : InMux
    port map (
            O => \N__65983\,
            I => \N__65928\
        );

    \I__14874\ : InMux
    port map (
            O => \N__65980\,
            I => \N__65928\
        );

    \I__14873\ : InMux
    port map (
            O => \N__65979\,
            I => \N__65917\
        );

    \I__14872\ : InMux
    port map (
            O => \N__65976\,
            I => \N__65917\
        );

    \I__14871\ : InMux
    port map (
            O => \N__65975\,
            I => \N__65917\
        );

    \I__14870\ : InMux
    port map (
            O => \N__65972\,
            I => \N__65917\
        );

    \I__14869\ : InMux
    port map (
            O => \N__65969\,
            I => \N__65917\
        );

    \I__14868\ : Span4Mux_h
    port map (
            O => \N__65966\,
            I => \N__65914\
        );

    \I__14867\ : LocalMux
    port map (
            O => \N__65963\,
            I => \N__65911\
        );

    \I__14866\ : Sp12to4
    port map (
            O => \N__65958\,
            I => \N__65908\
        );

    \I__14865\ : Span4Mux_v
    port map (
            O => \N__65955\,
            I => \N__65905\
        );

    \I__14864\ : InMux
    port map (
            O => \N__65952\,
            I => \N__65902\
        );

    \I__14863\ : Span4Mux_v
    port map (
            O => \N__65941\,
            I => \N__65897\
        );

    \I__14862\ : LocalMux
    port map (
            O => \N__65938\,
            I => \N__65897\
        );

    \I__14861\ : Span4Mux_h
    port map (
            O => \N__65935\,
            I => \N__65890\
        );

    \I__14860\ : LocalMux
    port map (
            O => \N__65928\,
            I => \N__65890\
        );

    \I__14859\ : LocalMux
    port map (
            O => \N__65917\,
            I => \N__65890\
        );

    \I__14858\ : Span4Mux_v
    port map (
            O => \N__65914\,
            I => \N__65887\
        );

    \I__14857\ : Span4Mux_v
    port map (
            O => \N__65911\,
            I => \N__65884\
        );

    \I__14856\ : Span12Mux_s10_v
    port map (
            O => \N__65908\,
            I => \N__65877\
        );

    \I__14855\ : Sp12to4
    port map (
            O => \N__65905\,
            I => \N__65877\
        );

    \I__14854\ : LocalMux
    port map (
            O => \N__65902\,
            I => \N__65877\
        );

    \I__14853\ : Span4Mux_h
    port map (
            O => \N__65897\,
            I => \N__65872\
        );

    \I__14852\ : Span4Mux_h
    port map (
            O => \N__65890\,
            I => \N__65872\
        );

    \I__14851\ : Odrv4
    port map (
            O => \N__65887\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n132\
        );

    \I__14850\ : Odrv4
    port map (
            O => \N__65884\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n132\
        );

    \I__14849\ : Odrv12
    port map (
            O => \N__65877\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n132\
        );

    \I__14848\ : Odrv4
    port map (
            O => \N__65872\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n132\
        );

    \I__14847\ : InMux
    port map (
            O => \N__65863\,
            I => \N__65860\
        );

    \I__14846\ : LocalMux
    port map (
            O => \N__65860\,
            I => \N__65857\
        );

    \I__14845\ : Odrv12
    port map (
            O => \N__65857\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n562\
        );

    \I__14844\ : InMux
    port map (
            O => \N__65854\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18273\
        );

    \I__14843\ : InMux
    port map (
            O => \N__65851\,
            I => \N__65848\
        );

    \I__14842\ : LocalMux
    port map (
            O => \N__65848\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n565\
        );

    \I__14841\ : CascadeMux
    port map (
            O => \N__65845\,
            I => \N__65840\
        );

    \I__14840\ : CascadeMux
    port map (
            O => \N__65844\,
            I => \N__65836\
        );

    \I__14839\ : CascadeMux
    port map (
            O => \N__65843\,
            I => \N__65833\
        );

    \I__14838\ : InMux
    port map (
            O => \N__65840\,
            I => \N__65825\
        );

    \I__14837\ : CascadeMux
    port map (
            O => \N__65839\,
            I => \N__65822\
        );

    \I__14836\ : InMux
    port map (
            O => \N__65836\,
            I => \N__65819\
        );

    \I__14835\ : InMux
    port map (
            O => \N__65833\,
            I => \N__65816\
        );

    \I__14834\ : CascadeMux
    port map (
            O => \N__65832\,
            I => \N__65813\
        );

    \I__14833\ : CascadeMux
    port map (
            O => \N__65831\,
            I => \N__65810\
        );

    \I__14832\ : CascadeMux
    port map (
            O => \N__65830\,
            I => \N__65804\
        );

    \I__14831\ : CascadeMux
    port map (
            O => \N__65829\,
            I => \N__65801\
        );

    \I__14830\ : CascadeMux
    port map (
            O => \N__65828\,
            I => \N__65798\
        );

    \I__14829\ : LocalMux
    port map (
            O => \N__65825\,
            I => \N__65795\
        );

    \I__14828\ : InMux
    port map (
            O => \N__65822\,
            I => \N__65792\
        );

    \I__14827\ : LocalMux
    port map (
            O => \N__65819\,
            I => \N__65786\
        );

    \I__14826\ : LocalMux
    port map (
            O => \N__65816\,
            I => \N__65786\
        );

    \I__14825\ : InMux
    port map (
            O => \N__65813\,
            I => \N__65783\
        );

    \I__14824\ : InMux
    port map (
            O => \N__65810\,
            I => \N__65780\
        );

    \I__14823\ : CascadeMux
    port map (
            O => \N__65809\,
            I => \N__65777\
        );

    \I__14822\ : CascadeMux
    port map (
            O => \N__65808\,
            I => \N__65773\
        );

    \I__14821\ : CascadeMux
    port map (
            O => \N__65807\,
            I => \N__65770\
        );

    \I__14820\ : InMux
    port map (
            O => \N__65804\,
            I => \N__65767\
        );

    \I__14819\ : InMux
    port map (
            O => \N__65801\,
            I => \N__65764\
        );

    \I__14818\ : InMux
    port map (
            O => \N__65798\,
            I => \N__65761\
        );

    \I__14817\ : Span4Mux_v
    port map (
            O => \N__65795\,
            I => \N__65756\
        );

    \I__14816\ : LocalMux
    port map (
            O => \N__65792\,
            I => \N__65756\
        );

    \I__14815\ : CascadeMux
    port map (
            O => \N__65791\,
            I => \N__65753\
        );

    \I__14814\ : Span4Mux_v
    port map (
            O => \N__65786\,
            I => \N__65746\
        );

    \I__14813\ : LocalMux
    port map (
            O => \N__65783\,
            I => \N__65746\
        );

    \I__14812\ : LocalMux
    port map (
            O => \N__65780\,
            I => \N__65746\
        );

    \I__14811\ : InMux
    port map (
            O => \N__65777\,
            I => \N__65743\
        );

    \I__14810\ : CascadeMux
    port map (
            O => \N__65776\,
            I => \N__65740\
        );

    \I__14809\ : InMux
    port map (
            O => \N__65773\,
            I => \N__65731\
        );

    \I__14808\ : InMux
    port map (
            O => \N__65770\,
            I => \N__65728\
        );

    \I__14807\ : LocalMux
    port map (
            O => \N__65767\,
            I => \N__65725\
        );

    \I__14806\ : LocalMux
    port map (
            O => \N__65764\,
            I => \N__65718\
        );

    \I__14805\ : LocalMux
    port map (
            O => \N__65761\,
            I => \N__65718\
        );

    \I__14804\ : Span4Mux_h
    port map (
            O => \N__65756\,
            I => \N__65718\
        );

    \I__14803\ : InMux
    port map (
            O => \N__65753\,
            I => \N__65715\
        );

    \I__14802\ : Span4Mux_h
    port map (
            O => \N__65746\,
            I => \N__65710\
        );

    \I__14801\ : LocalMux
    port map (
            O => \N__65743\,
            I => \N__65710\
        );

    \I__14800\ : InMux
    port map (
            O => \N__65740\,
            I => \N__65707\
        );

    \I__14799\ : InMux
    port map (
            O => \N__65739\,
            I => \N__65704\
        );

    \I__14798\ : CascadeMux
    port map (
            O => \N__65738\,
            I => \N__65701\
        );

    \I__14797\ : CascadeMux
    port map (
            O => \N__65737\,
            I => \N__65698\
        );

    \I__14796\ : CascadeMux
    port map (
            O => \N__65736\,
            I => \N__65694\
        );

    \I__14795\ : CascadeMux
    port map (
            O => \N__65735\,
            I => \N__65691\
        );

    \I__14794\ : CascadeMux
    port map (
            O => \N__65734\,
            I => \N__65688\
        );

    \I__14793\ : LocalMux
    port map (
            O => \N__65731\,
            I => \N__65683\
        );

    \I__14792\ : LocalMux
    port map (
            O => \N__65728\,
            I => \N__65683\
        );

    \I__14791\ : Span4Mux_h
    port map (
            O => \N__65725\,
            I => \N__65680\
        );

    \I__14790\ : Span4Mux_v
    port map (
            O => \N__65718\,
            I => \N__65675\
        );

    \I__14789\ : LocalMux
    port map (
            O => \N__65715\,
            I => \N__65675\
        );

    \I__14788\ : Span4Mux_v
    port map (
            O => \N__65710\,
            I => \N__65670\
        );

    \I__14787\ : LocalMux
    port map (
            O => \N__65707\,
            I => \N__65670\
        );

    \I__14786\ : LocalMux
    port map (
            O => \N__65704\,
            I => \N__65667\
        );

    \I__14785\ : InMux
    port map (
            O => \N__65701\,
            I => \N__65662\
        );

    \I__14784\ : InMux
    port map (
            O => \N__65698\,
            I => \N__65662\
        );

    \I__14783\ : InMux
    port map (
            O => \N__65697\,
            I => \N__65653\
        );

    \I__14782\ : InMux
    port map (
            O => \N__65694\,
            I => \N__65653\
        );

    \I__14781\ : InMux
    port map (
            O => \N__65691\,
            I => \N__65653\
        );

    \I__14780\ : InMux
    port map (
            O => \N__65688\,
            I => \N__65653\
        );

    \I__14779\ : Span4Mux_v
    port map (
            O => \N__65683\,
            I => \N__65648\
        );

    \I__14778\ : Span4Mux_h
    port map (
            O => \N__65680\,
            I => \N__65648\
        );

    \I__14777\ : Span4Mux_h
    port map (
            O => \N__65675\,
            I => \N__65645\
        );

    \I__14776\ : Span4Mux_v
    port map (
            O => \N__65670\,
            I => \N__65636\
        );

    \I__14775\ : Span4Mux_h
    port map (
            O => \N__65667\,
            I => \N__65636\
        );

    \I__14774\ : LocalMux
    port map (
            O => \N__65662\,
            I => \N__65636\
        );

    \I__14773\ : LocalMux
    port map (
            O => \N__65653\,
            I => \N__65636\
        );

    \I__14772\ : Odrv4
    port map (
            O => \N__65648\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n135\
        );

    \I__14771\ : Odrv4
    port map (
            O => \N__65645\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n135\
        );

    \I__14770\ : Odrv4
    port map (
            O => \N__65636\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n135\
        );

    \I__14769\ : InMux
    port map (
            O => \N__65629\,
            I => \N__65626\
        );

    \I__14768\ : LocalMux
    port map (
            O => \N__65626\,
            I => \N__65623\
        );

    \I__14767\ : Odrv4
    port map (
            O => \N__65623\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n611\
        );

    \I__14766\ : InMux
    port map (
            O => \N__65620\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18274\
        );

    \I__14765\ : InMux
    port map (
            O => \N__65617\,
            I => \N__65614\
        );

    \I__14764\ : LocalMux
    port map (
            O => \N__65614\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n614\
        );

    \I__14763\ : CascadeMux
    port map (
            O => \N__65611\,
            I => \N__65606\
        );

    \I__14762\ : CascadeMux
    port map (
            O => \N__65610\,
            I => \N__65603\
        );

    \I__14761\ : CascadeMux
    port map (
            O => \N__65609\,
            I => \N__65597\
        );

    \I__14760\ : InMux
    port map (
            O => \N__65606\,
            I => \N__65592\
        );

    \I__14759\ : InMux
    port map (
            O => \N__65603\,
            I => \N__65589\
        );

    \I__14758\ : CascadeMux
    port map (
            O => \N__65602\,
            I => \N__65586\
        );

    \I__14757\ : CascadeMux
    port map (
            O => \N__65601\,
            I => \N__65583\
        );

    \I__14756\ : CascadeMux
    port map (
            O => \N__65600\,
            I => \N__65577\
        );

    \I__14755\ : InMux
    port map (
            O => \N__65597\,
            I => \N__65574\
        );

    \I__14754\ : CascadeMux
    port map (
            O => \N__65596\,
            I => \N__65571\
        );

    \I__14753\ : InMux
    port map (
            O => \N__65595\,
            I => \N__65567\
        );

    \I__14752\ : LocalMux
    port map (
            O => \N__65592\,
            I => \N__65562\
        );

    \I__14751\ : LocalMux
    port map (
            O => \N__65589\,
            I => \N__65562\
        );

    \I__14750\ : InMux
    port map (
            O => \N__65586\,
            I => \N__65559\
        );

    \I__14749\ : InMux
    port map (
            O => \N__65583\,
            I => \N__65556\
        );

    \I__14748\ : CascadeMux
    port map (
            O => \N__65582\,
            I => \N__65553\
        );

    \I__14747\ : CascadeMux
    port map (
            O => \N__65581\,
            I => \N__65550\
        );

    \I__14746\ : CascadeMux
    port map (
            O => \N__65580\,
            I => \N__65547\
        );

    \I__14745\ : InMux
    port map (
            O => \N__65577\,
            I => \N__65543\
        );

    \I__14744\ : LocalMux
    port map (
            O => \N__65574\,
            I => \N__65540\
        );

    \I__14743\ : InMux
    port map (
            O => \N__65571\,
            I => \N__65537\
        );

    \I__14742\ : CascadeMux
    port map (
            O => \N__65570\,
            I => \N__65534\
        );

    \I__14741\ : LocalMux
    port map (
            O => \N__65567\,
            I => \N__65531\
        );

    \I__14740\ : Span4Mux_v
    port map (
            O => \N__65562\,
            I => \N__65524\
        );

    \I__14739\ : LocalMux
    port map (
            O => \N__65559\,
            I => \N__65524\
        );

    \I__14738\ : LocalMux
    port map (
            O => \N__65556\,
            I => \N__65524\
        );

    \I__14737\ : InMux
    port map (
            O => \N__65553\,
            I => \N__65521\
        );

    \I__14736\ : InMux
    port map (
            O => \N__65550\,
            I => \N__65518\
        );

    \I__14735\ : InMux
    port map (
            O => \N__65547\,
            I => \N__65515\
        );

    \I__14734\ : CascadeMux
    port map (
            O => \N__65546\,
            I => \N__65512\
        );

    \I__14733\ : LocalMux
    port map (
            O => \N__65543\,
            I => \N__65504\
        );

    \I__14732\ : Span4Mux_h
    port map (
            O => \N__65540\,
            I => \N__65499\
        );

    \I__14731\ : LocalMux
    port map (
            O => \N__65537\,
            I => \N__65499\
        );

    \I__14730\ : InMux
    port map (
            O => \N__65534\,
            I => \N__65496\
        );

    \I__14729\ : Span4Mux_v
    port map (
            O => \N__65531\,
            I => \N__65493\
        );

    \I__14728\ : Span4Mux_h
    port map (
            O => \N__65524\,
            I => \N__65483\
        );

    \I__14727\ : LocalMux
    port map (
            O => \N__65521\,
            I => \N__65483\
        );

    \I__14726\ : LocalMux
    port map (
            O => \N__65518\,
            I => \N__65483\
        );

    \I__14725\ : LocalMux
    port map (
            O => \N__65515\,
            I => \N__65483\
        );

    \I__14724\ : InMux
    port map (
            O => \N__65512\,
            I => \N__65480\
        );

    \I__14723\ : InMux
    port map (
            O => \N__65511\,
            I => \N__65477\
        );

    \I__14722\ : InMux
    port map (
            O => \N__65510\,
            I => \N__65468\
        );

    \I__14721\ : InMux
    port map (
            O => \N__65509\,
            I => \N__65468\
        );

    \I__14720\ : InMux
    port map (
            O => \N__65508\,
            I => \N__65468\
        );

    \I__14719\ : InMux
    port map (
            O => \N__65507\,
            I => \N__65468\
        );

    \I__14718\ : Span4Mux_h
    port map (
            O => \N__65504\,
            I => \N__65464\
        );

    \I__14717\ : Span4Mux_v
    port map (
            O => \N__65499\,
            I => \N__65459\
        );

    \I__14716\ : LocalMux
    port map (
            O => \N__65496\,
            I => \N__65459\
        );

    \I__14715\ : Span4Mux_h
    port map (
            O => \N__65493\,
            I => \N__65456\
        );

    \I__14714\ : InMux
    port map (
            O => \N__65492\,
            I => \N__65453\
        );

    \I__14713\ : Span4Mux_v
    port map (
            O => \N__65483\,
            I => \N__65448\
        );

    \I__14712\ : LocalMux
    port map (
            O => \N__65480\,
            I => \N__65448\
        );

    \I__14711\ : LocalMux
    port map (
            O => \N__65477\,
            I => \N__65445\
        );

    \I__14710\ : LocalMux
    port map (
            O => \N__65468\,
            I => \N__65442\
        );

    \I__14709\ : InMux
    port map (
            O => \N__65467\,
            I => \N__65439\
        );

    \I__14708\ : Span4Mux_v
    port map (
            O => \N__65464\,
            I => \N__65432\
        );

    \I__14707\ : Span4Mux_h
    port map (
            O => \N__65459\,
            I => \N__65432\
        );

    \I__14706\ : Sp12to4
    port map (
            O => \N__65456\,
            I => \N__65427\
        );

    \I__14705\ : LocalMux
    port map (
            O => \N__65453\,
            I => \N__65427\
        );

    \I__14704\ : Span4Mux_v
    port map (
            O => \N__65448\,
            I => \N__65418\
        );

    \I__14703\ : Span4Mux_v
    port map (
            O => \N__65445\,
            I => \N__65418\
        );

    \I__14702\ : Span4Mux_v
    port map (
            O => \N__65442\,
            I => \N__65418\
        );

    \I__14701\ : LocalMux
    port map (
            O => \N__65439\,
            I => \N__65418\
        );

    \I__14700\ : InMux
    port map (
            O => \N__65438\,
            I => \N__65413\
        );

    \I__14699\ : InMux
    port map (
            O => \N__65437\,
            I => \N__65413\
        );

    \I__14698\ : Odrv4
    port map (
            O => \N__65432\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n138\
        );

    \I__14697\ : Odrv12
    port map (
            O => \N__65427\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n138\
        );

    \I__14696\ : Odrv4
    port map (
            O => \N__65418\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n138\
        );

    \I__14695\ : LocalMux
    port map (
            O => \N__65413\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n138\
        );

    \I__14694\ : CascadeMux
    port map (
            O => \N__65404\,
            I => \N__65401\
        );

    \I__14693\ : InMux
    port map (
            O => \N__65401\,
            I => \N__65398\
        );

    \I__14692\ : LocalMux
    port map (
            O => \N__65398\,
            I => \N__65395\
        );

    \I__14691\ : Odrv4
    port map (
            O => \N__65395\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n660\
        );

    \I__14690\ : InMux
    port map (
            O => \N__65392\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18275\
        );

    \I__14689\ : InMux
    port map (
            O => \N__65389\,
            I => \N__65381\
        );

    \I__14688\ : InMux
    port map (
            O => \N__65388\,
            I => \N__65378\
        );

    \I__14687\ : InMux
    port map (
            O => \N__65387\,
            I => \N__65375\
        );

    \I__14686\ : CascadeMux
    port map (
            O => \N__65386\,
            I => \N__65371\
        );

    \I__14685\ : InMux
    port map (
            O => \N__65385\,
            I => \N__65368\
        );

    \I__14684\ : InMux
    port map (
            O => \N__65384\,
            I => \N__65365\
        );

    \I__14683\ : LocalMux
    port map (
            O => \N__65381\,
            I => \N__65362\
        );

    \I__14682\ : LocalMux
    port map (
            O => \N__65378\,
            I => \N__65356\
        );

    \I__14681\ : LocalMux
    port map (
            O => \N__65375\,
            I => \N__65356\
        );

    \I__14680\ : InMux
    port map (
            O => \N__65374\,
            I => \N__65353\
        );

    \I__14679\ : InMux
    port map (
            O => \N__65371\,
            I => \N__65349\
        );

    \I__14678\ : LocalMux
    port map (
            O => \N__65368\,
            I => \N__65343\
        );

    \I__14677\ : LocalMux
    port map (
            O => \N__65365\,
            I => \N__65343\
        );

    \I__14676\ : Span4Mux_v
    port map (
            O => \N__65362\,
            I => \N__65338\
        );

    \I__14675\ : InMux
    port map (
            O => \N__65361\,
            I => \N__65335\
        );

    \I__14674\ : Span4Mux_h
    port map (
            O => \N__65356\,
            I => \N__65330\
        );

    \I__14673\ : LocalMux
    port map (
            O => \N__65353\,
            I => \N__65330\
        );

    \I__14672\ : InMux
    port map (
            O => \N__65352\,
            I => \N__65327\
        );

    \I__14671\ : LocalMux
    port map (
            O => \N__65349\,
            I => \N__65324\
        );

    \I__14670\ : InMux
    port map (
            O => \N__65348\,
            I => \N__65321\
        );

    \I__14669\ : Span4Mux_h
    port map (
            O => \N__65343\,
            I => \N__65317\
        );

    \I__14668\ : InMux
    port map (
            O => \N__65342\,
            I => \N__65314\
        );

    \I__14667\ : InMux
    port map (
            O => \N__65341\,
            I => \N__65310\
        );

    \I__14666\ : Span4Mux_h
    port map (
            O => \N__65338\,
            I => \N__65301\
        );

    \I__14665\ : LocalMux
    port map (
            O => \N__65335\,
            I => \N__65301\
        );

    \I__14664\ : Span4Mux_h
    port map (
            O => \N__65330\,
            I => \N__65301\
        );

    \I__14663\ : LocalMux
    port map (
            O => \N__65327\,
            I => \N__65301\
        );

    \I__14662\ : Span4Mux_v
    port map (
            O => \N__65324\,
            I => \N__65296\
        );

    \I__14661\ : LocalMux
    port map (
            O => \N__65321\,
            I => \N__65296\
        );

    \I__14660\ : InMux
    port map (
            O => \N__65320\,
            I => \N__65293\
        );

    \I__14659\ : Span4Mux_v
    port map (
            O => \N__65317\,
            I => \N__65288\
        );

    \I__14658\ : LocalMux
    port map (
            O => \N__65314\,
            I => \N__65288\
        );

    \I__14657\ : InMux
    port map (
            O => \N__65313\,
            I => \N__65285\
        );

    \I__14656\ : LocalMux
    port map (
            O => \N__65310\,
            I => \N__65281\
        );

    \I__14655\ : Span4Mux_v
    port map (
            O => \N__65301\,
            I => \N__65274\
        );

    \I__14654\ : Span4Mux_v
    port map (
            O => \N__65296\,
            I => \N__65274\
        );

    \I__14653\ : LocalMux
    port map (
            O => \N__65293\,
            I => \N__65274\
        );

    \I__14652\ : Span4Mux_h
    port map (
            O => \N__65288\,
            I => \N__65271\
        );

    \I__14651\ : LocalMux
    port map (
            O => \N__65285\,
            I => \N__65268\
        );

    \I__14650\ : InMux
    port map (
            O => \N__65284\,
            I => \N__65265\
        );

    \I__14649\ : Span4Mux_h
    port map (
            O => \N__65281\,
            I => \N__65261\
        );

    \I__14648\ : Span4Mux_h
    port map (
            O => \N__65274\,
            I => \N__65258\
        );

    \I__14647\ : Span4Mux_h
    port map (
            O => \N__65271\,
            I => \N__65251\
        );

    \I__14646\ : Span4Mux_v
    port map (
            O => \N__65268\,
            I => \N__65251\
        );

    \I__14645\ : LocalMux
    port map (
            O => \N__65265\,
            I => \N__65251\
        );

    \I__14644\ : CascadeMux
    port map (
            O => \N__65264\,
            I => \N__65248\
        );

    \I__14643\ : Sp12to4
    port map (
            O => \N__65261\,
            I => \N__65245\
        );

    \I__14642\ : Span4Mux_v
    port map (
            O => \N__65258\,
            I => \N__65242\
        );

    \I__14641\ : Span4Mux_h
    port map (
            O => \N__65251\,
            I => \N__65239\
        );

    \I__14640\ : InMux
    port map (
            O => \N__65248\,
            I => \N__65236\
        );

    \I__14639\ : Odrv12
    port map (
            O => \N__65245\,
            I => n141_adj_2421
        );

    \I__14638\ : Odrv4
    port map (
            O => \N__65242\,
            I => n141_adj_2421
        );

    \I__14637\ : Odrv4
    port map (
            O => \N__65239\,
            I => n141_adj_2421
        );

    \I__14636\ : LocalMux
    port map (
            O => \N__65236\,
            I => n141_adj_2421
        );

    \I__14635\ : CascadeMux
    port map (
            O => \N__65227\,
            I => \N__65224\
        );

    \I__14634\ : InMux
    port map (
            O => \N__65224\,
            I => \N__65221\
        );

    \I__14633\ : LocalMux
    port map (
            O => \N__65221\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n663\
        );

    \I__14632\ : CascadeMux
    port map (
            O => \N__65218\,
            I => \N__65215\
        );

    \I__14631\ : InMux
    port map (
            O => \N__65215\,
            I => \N__65212\
        );

    \I__14630\ : LocalMux
    port map (
            O => \N__65212\,
            I => \N__65209\
        );

    \I__14629\ : Odrv12
    port map (
            O => \N__65209\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n709\
        );

    \I__14628\ : InMux
    port map (
            O => \N__65206\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18276\
        );

    \I__14627\ : InMux
    port map (
            O => \N__65203\,
            I => \N__65198\
        );

    \I__14626\ : InMux
    port map (
            O => \N__65202\,
            I => \N__65195\
        );

    \I__14625\ : InMux
    port map (
            O => \N__65201\,
            I => \N__65189\
        );

    \I__14624\ : LocalMux
    port map (
            O => \N__65198\,
            I => \N__65185\
        );

    \I__14623\ : LocalMux
    port map (
            O => \N__65195\,
            I => \N__65182\
        );

    \I__14622\ : InMux
    port map (
            O => \N__65194\,
            I => \N__65179\
        );

    \I__14621\ : InMux
    port map (
            O => \N__65193\,
            I => \N__65175\
        );

    \I__14620\ : InMux
    port map (
            O => \N__65192\,
            I => \N__65172\
        );

    \I__14619\ : LocalMux
    port map (
            O => \N__65189\,
            I => \N__65166\
        );

    \I__14618\ : CascadeMux
    port map (
            O => \N__65188\,
            I => \N__65163\
        );

    \I__14617\ : Span4Mux_v
    port map (
            O => \N__65185\,
            I => \N__65156\
        );

    \I__14616\ : Span4Mux_h
    port map (
            O => \N__65182\,
            I => \N__65156\
        );

    \I__14615\ : LocalMux
    port map (
            O => \N__65179\,
            I => \N__65156\
        );

    \I__14614\ : CascadeMux
    port map (
            O => \N__65178\,
            I => \N__65153\
        );

    \I__14613\ : LocalMux
    port map (
            O => \N__65175\,
            I => \N__65149\
        );

    \I__14612\ : LocalMux
    port map (
            O => \N__65172\,
            I => \N__65146\
        );

    \I__14611\ : InMux
    port map (
            O => \N__65171\,
            I => \N__65143\
        );

    \I__14610\ : InMux
    port map (
            O => \N__65170\,
            I => \N__65140\
        );

    \I__14609\ : CascadeMux
    port map (
            O => \N__65169\,
            I => \N__65136\
        );

    \I__14608\ : Span4Mux_v
    port map (
            O => \N__65166\,
            I => \N__65132\
        );

    \I__14607\ : InMux
    port map (
            O => \N__65163\,
            I => \N__65129\
        );

    \I__14606\ : Span4Mux_v
    port map (
            O => \N__65156\,
            I => \N__65126\
        );

    \I__14605\ : InMux
    port map (
            O => \N__65153\,
            I => \N__65123\
        );

    \I__14604\ : CascadeMux
    port map (
            O => \N__65152\,
            I => \N__65120\
        );

    \I__14603\ : Span4Mux_h
    port map (
            O => \N__65149\,
            I => \N__65109\
        );

    \I__14602\ : Span4Mux_v
    port map (
            O => \N__65146\,
            I => \N__65109\
        );

    \I__14601\ : LocalMux
    port map (
            O => \N__65143\,
            I => \N__65109\
        );

    \I__14600\ : LocalMux
    port map (
            O => \N__65140\,
            I => \N__65109\
        );

    \I__14599\ : InMux
    port map (
            O => \N__65139\,
            I => \N__65106\
        );

    \I__14598\ : InMux
    port map (
            O => \N__65136\,
            I => \N__65103\
        );

    \I__14597\ : InMux
    port map (
            O => \N__65135\,
            I => \N__65100\
        );

    \I__14596\ : Span4Mux_h
    port map (
            O => \N__65132\,
            I => \N__65095\
        );

    \I__14595\ : LocalMux
    port map (
            O => \N__65129\,
            I => \N__65095\
        );

    \I__14594\ : Span4Mux_h
    port map (
            O => \N__65126\,
            I => \N__65090\
        );

    \I__14593\ : LocalMux
    port map (
            O => \N__65123\,
            I => \N__65090\
        );

    \I__14592\ : InMux
    port map (
            O => \N__65120\,
            I => \N__65087\
        );

    \I__14591\ : InMux
    port map (
            O => \N__65119\,
            I => \N__65082\
        );

    \I__14590\ : InMux
    port map (
            O => \N__65118\,
            I => \N__65082\
        );

    \I__14589\ : Span4Mux_v
    port map (
            O => \N__65109\,
            I => \N__65077\
        );

    \I__14588\ : LocalMux
    port map (
            O => \N__65106\,
            I => \N__65077\
        );

    \I__14587\ : LocalMux
    port map (
            O => \N__65103\,
            I => \N__65072\
        );

    \I__14586\ : LocalMux
    port map (
            O => \N__65100\,
            I => \N__65072\
        );

    \I__14585\ : Span4Mux_v
    port map (
            O => \N__65095\,
            I => \N__65065\
        );

    \I__14584\ : Span4Mux_h
    port map (
            O => \N__65090\,
            I => \N__65065\
        );

    \I__14583\ : LocalMux
    port map (
            O => \N__65087\,
            I => \N__65065\
        );

    \I__14582\ : LocalMux
    port map (
            O => \N__65082\,
            I => \N__65062\
        );

    \I__14581\ : Span4Mux_v
    port map (
            O => \N__65077\,
            I => \N__65058\
        );

    \I__14580\ : Span12Mux_v
    port map (
            O => \N__65072\,
            I => \N__65055\
        );

    \I__14579\ : Span4Mux_v
    port map (
            O => \N__65065\,
            I => \N__65050\
        );

    \I__14578\ : Span4Mux_h
    port map (
            O => \N__65062\,
            I => \N__65050\
        );

    \I__14577\ : InMux
    port map (
            O => \N__65061\,
            I => \N__65047\
        );

    \I__14576\ : Odrv4
    port map (
            O => \N__65058\,
            I => n146_adj_2423
        );

    \I__14575\ : Odrv12
    port map (
            O => \N__65055\,
            I => n146_adj_2423
        );

    \I__14574\ : Odrv4
    port map (
            O => \N__65050\,
            I => n146_adj_2423
        );

    \I__14573\ : LocalMux
    port map (
            O => \N__65047\,
            I => n146_adj_2423
        );

    \I__14572\ : CascadeMux
    port map (
            O => \N__65038\,
            I => \N__65035\
        );

    \I__14571\ : InMux
    port map (
            O => \N__65035\,
            I => \N__65032\
        );

    \I__14570\ : LocalMux
    port map (
            O => \N__65032\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n712\
        );

    \I__14569\ : InMux
    port map (
            O => \N__65029\,
            I => \N__65026\
        );

    \I__14568\ : LocalMux
    port map (
            O => \N__65026\,
            I => \N__65023\
        );

    \I__14567\ : Span12Mux_h
    port map (
            O => \N__65023\,
            I => \N__65020\
        );

    \I__14566\ : Odrv12
    port map (
            O => \N__65020\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n766\
        );

    \I__14565\ : CascadeMux
    port map (
            O => \N__65017\,
            I => \N__65001\
        );

    \I__14564\ : CascadeMux
    port map (
            O => \N__65016\,
            I => \N__64998\
        );

    \I__14563\ : CascadeMux
    port map (
            O => \N__65015\,
            I => \N__64995\
        );

    \I__14562\ : CascadeMux
    port map (
            O => \N__65014\,
            I => \N__64992\
        );

    \I__14561\ : CascadeMux
    port map (
            O => \N__65013\,
            I => \N__64989\
        );

    \I__14560\ : CascadeMux
    port map (
            O => \N__65012\,
            I => \N__64986\
        );

    \I__14559\ : CascadeMux
    port map (
            O => \N__65011\,
            I => \N__64983\
        );

    \I__14558\ : CascadeMux
    port map (
            O => \N__65010\,
            I => \N__64980\
        );

    \I__14557\ : CascadeMux
    port map (
            O => \N__65009\,
            I => \N__64977\
        );

    \I__14556\ : CascadeMux
    port map (
            O => \N__65008\,
            I => \N__64974\
        );

    \I__14555\ : CascadeMux
    port map (
            O => \N__65007\,
            I => \N__64971\
        );

    \I__14554\ : CascadeMux
    port map (
            O => \N__65006\,
            I => \N__64968\
        );

    \I__14553\ : CascadeMux
    port map (
            O => \N__65005\,
            I => \N__64965\
        );

    \I__14552\ : CascadeMux
    port map (
            O => \N__65004\,
            I => \N__64961\
        );

    \I__14551\ : InMux
    port map (
            O => \N__65001\,
            I => \N__64957\
        );

    \I__14550\ : InMux
    port map (
            O => \N__64998\,
            I => \N__64948\
        );

    \I__14549\ : InMux
    port map (
            O => \N__64995\,
            I => \N__64948\
        );

    \I__14548\ : InMux
    port map (
            O => \N__64992\,
            I => \N__64948\
        );

    \I__14547\ : InMux
    port map (
            O => \N__64989\,
            I => \N__64940\
        );

    \I__14546\ : InMux
    port map (
            O => \N__64986\,
            I => \N__64940\
        );

    \I__14545\ : InMux
    port map (
            O => \N__64983\,
            I => \N__64940\
        );

    \I__14544\ : InMux
    port map (
            O => \N__64980\,
            I => \N__64933\
        );

    \I__14543\ : InMux
    port map (
            O => \N__64977\,
            I => \N__64933\
        );

    \I__14542\ : InMux
    port map (
            O => \N__64974\,
            I => \N__64933\
        );

    \I__14541\ : InMux
    port map (
            O => \N__64971\,
            I => \N__64922\
        );

    \I__14540\ : InMux
    port map (
            O => \N__64968\,
            I => \N__64922\
        );

    \I__14539\ : InMux
    port map (
            O => \N__64965\,
            I => \N__64922\
        );

    \I__14538\ : InMux
    port map (
            O => \N__64964\,
            I => \N__64922\
        );

    \I__14537\ : InMux
    port map (
            O => \N__64961\,
            I => \N__64922\
        );

    \I__14536\ : InMux
    port map (
            O => \N__64960\,
            I => \N__64918\
        );

    \I__14535\ : LocalMux
    port map (
            O => \N__64957\,
            I => \N__64915\
        );

    \I__14534\ : InMux
    port map (
            O => \N__64956\,
            I => \N__64911\
        );

    \I__14533\ : CascadeMux
    port map (
            O => \N__64955\,
            I => \N__64907\
        );

    \I__14532\ : LocalMux
    port map (
            O => \N__64948\,
            I => \N__64904\
        );

    \I__14531\ : InMux
    port map (
            O => \N__64947\,
            I => \N__64901\
        );

    \I__14530\ : LocalMux
    port map (
            O => \N__64940\,
            I => \N__64892\
        );

    \I__14529\ : LocalMux
    port map (
            O => \N__64933\,
            I => \N__64892\
        );

    \I__14528\ : LocalMux
    port map (
            O => \N__64922\,
            I => \N__64892\
        );

    \I__14527\ : InMux
    port map (
            O => \N__64921\,
            I => \N__64889\
        );

    \I__14526\ : LocalMux
    port map (
            O => \N__64918\,
            I => \N__64884\
        );

    \I__14525\ : Span4Mux_v
    port map (
            O => \N__64915\,
            I => \N__64881\
        );

    \I__14524\ : InMux
    port map (
            O => \N__64914\,
            I => \N__64878\
        );

    \I__14523\ : LocalMux
    port map (
            O => \N__64911\,
            I => \N__64875\
        );

    \I__14522\ : InMux
    port map (
            O => \N__64910\,
            I => \N__64872\
        );

    \I__14521\ : InMux
    port map (
            O => \N__64907\,
            I => \N__64869\
        );

    \I__14520\ : Span4Mux_v
    port map (
            O => \N__64904\,
            I => \N__64864\
        );

    \I__14519\ : LocalMux
    port map (
            O => \N__64901\,
            I => \N__64864\
        );

    \I__14518\ : CascadeMux
    port map (
            O => \N__64900\,
            I => \N__64859\
        );

    \I__14517\ : InMux
    port map (
            O => \N__64899\,
            I => \N__64856\
        );

    \I__14516\ : Span4Mux_v
    port map (
            O => \N__64892\,
            I => \N__64851\
        );

    \I__14515\ : LocalMux
    port map (
            O => \N__64889\,
            I => \N__64851\
        );

    \I__14514\ : InMux
    port map (
            O => \N__64888\,
            I => \N__64848\
        );

    \I__14513\ : CascadeMux
    port map (
            O => \N__64887\,
            I => \N__64845\
        );

    \I__14512\ : Span4Mux_v
    port map (
            O => \N__64884\,
            I => \N__64837\
        );

    \I__14511\ : Span4Mux_h
    port map (
            O => \N__64881\,
            I => \N__64837\
        );

    \I__14510\ : LocalMux
    port map (
            O => \N__64878\,
            I => \N__64837\
        );

    \I__14509\ : Span4Mux_v
    port map (
            O => \N__64875\,
            I => \N__64832\
        );

    \I__14508\ : LocalMux
    port map (
            O => \N__64872\,
            I => \N__64832\
        );

    \I__14507\ : LocalMux
    port map (
            O => \N__64869\,
            I => \N__64829\
        );

    \I__14506\ : Span4Mux_v
    port map (
            O => \N__64864\,
            I => \N__64826\
        );

    \I__14505\ : InMux
    port map (
            O => \N__64863\,
            I => \N__64823\
        );

    \I__14504\ : InMux
    port map (
            O => \N__64862\,
            I => \N__64820\
        );

    \I__14503\ : InMux
    port map (
            O => \N__64859\,
            I => \N__64817\
        );

    \I__14502\ : LocalMux
    port map (
            O => \N__64856\,
            I => \N__64810\
        );

    \I__14501\ : Span4Mux_h
    port map (
            O => \N__64851\,
            I => \N__64810\
        );

    \I__14500\ : LocalMux
    port map (
            O => \N__64848\,
            I => \N__64810\
        );

    \I__14499\ : InMux
    port map (
            O => \N__64845\,
            I => \N__64807\
        );

    \I__14498\ : CascadeMux
    port map (
            O => \N__64844\,
            I => \N__64804\
        );

    \I__14497\ : Span4Mux_v
    port map (
            O => \N__64837\,
            I => \N__64801\
        );

    \I__14496\ : Span4Mux_v
    port map (
            O => \N__64832\,
            I => \N__64798\
        );

    \I__14495\ : Span4Mux_v
    port map (
            O => \N__64829\,
            I => \N__64787\
        );

    \I__14494\ : Span4Mux_h
    port map (
            O => \N__64826\,
            I => \N__64787\
        );

    \I__14493\ : LocalMux
    port map (
            O => \N__64823\,
            I => \N__64787\
        );

    \I__14492\ : LocalMux
    port map (
            O => \N__64820\,
            I => \N__64787\
        );

    \I__14491\ : LocalMux
    port map (
            O => \N__64817\,
            I => \N__64787\
        );

    \I__14490\ : Span4Mux_v
    port map (
            O => \N__64810\,
            I => \N__64782\
        );

    \I__14489\ : LocalMux
    port map (
            O => \N__64807\,
            I => \N__64782\
        );

    \I__14488\ : InMux
    port map (
            O => \N__64804\,
            I => \N__64779\
        );

    \I__14487\ : Span4Mux_v
    port map (
            O => \N__64801\,
            I => \N__64776\
        );

    \I__14486\ : Span4Mux_h
    port map (
            O => \N__64798\,
            I => \N__64771\
        );

    \I__14485\ : Span4Mux_v
    port map (
            O => \N__64787\,
            I => \N__64771\
        );

    \I__14484\ : Span4Mux_v
    port map (
            O => \N__64782\,
            I => \N__64766\
        );

    \I__14483\ : LocalMux
    port map (
            O => \N__64779\,
            I => \N__64766\
        );

    \I__14482\ : Odrv4
    port map (
            O => \N__64776\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n102\
        );

    \I__14481\ : Odrv4
    port map (
            O => \N__64771\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n102\
        );

    \I__14480\ : Odrv4
    port map (
            O => \N__64766\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n102\
        );

    \I__14479\ : CascadeMux
    port map (
            O => \N__64759\,
            I => \N__64755\
        );

    \I__14478\ : CascadeMux
    port map (
            O => \N__64758\,
            I => \N__64750\
        );

    \I__14477\ : InMux
    port map (
            O => \N__64755\,
            I => \N__64744\
        );

    \I__14476\ : CascadeMux
    port map (
            O => \N__64754\,
            I => \N__64741\
        );

    \I__14475\ : CascadeMux
    port map (
            O => \N__64753\,
            I => \N__64738\
        );

    \I__14474\ : InMux
    port map (
            O => \N__64750\,
            I => \N__64735\
        );

    \I__14473\ : CascadeMux
    port map (
            O => \N__64749\,
            I => \N__64731\
        );

    \I__14472\ : CascadeMux
    port map (
            O => \N__64748\,
            I => \N__64728\
        );

    \I__14471\ : InMux
    port map (
            O => \N__64747\,
            I => \N__64723\
        );

    \I__14470\ : LocalMux
    port map (
            O => \N__64744\,
            I => \N__64720\
        );

    \I__14469\ : InMux
    port map (
            O => \N__64741\,
            I => \N__64717\
        );

    \I__14468\ : InMux
    port map (
            O => \N__64738\,
            I => \N__64714\
        );

    \I__14467\ : LocalMux
    port map (
            O => \N__64735\,
            I => \N__64709\
        );

    \I__14466\ : CascadeMux
    port map (
            O => \N__64734\,
            I => \N__64706\
        );

    \I__14465\ : InMux
    port map (
            O => \N__64731\,
            I => \N__64703\
        );

    \I__14464\ : InMux
    port map (
            O => \N__64728\,
            I => \N__64700\
        );

    \I__14463\ : CascadeMux
    port map (
            O => \N__64727\,
            I => \N__64697\
        );

    \I__14462\ : CascadeMux
    port map (
            O => \N__64726\,
            I => \N__64694\
        );

    \I__14461\ : LocalMux
    port map (
            O => \N__64723\,
            I => \N__64690\
        );

    \I__14460\ : Span4Mux_v
    port map (
            O => \N__64720\,
            I => \N__64683\
        );

    \I__14459\ : LocalMux
    port map (
            O => \N__64717\,
            I => \N__64683\
        );

    \I__14458\ : LocalMux
    port map (
            O => \N__64714\,
            I => \N__64683\
        );

    \I__14457\ : InMux
    port map (
            O => \N__64713\,
            I => \N__64680\
        );

    \I__14456\ : InMux
    port map (
            O => \N__64712\,
            I => \N__64677\
        );

    \I__14455\ : Span4Mux_v
    port map (
            O => \N__64709\,
            I => \N__64674\
        );

    \I__14454\ : InMux
    port map (
            O => \N__64706\,
            I => \N__64671\
        );

    \I__14453\ : LocalMux
    port map (
            O => \N__64703\,
            I => \N__64666\
        );

    \I__14452\ : LocalMux
    port map (
            O => \N__64700\,
            I => \N__64666\
        );

    \I__14451\ : InMux
    port map (
            O => \N__64697\,
            I => \N__64663\
        );

    \I__14450\ : InMux
    port map (
            O => \N__64694\,
            I => \N__64660\
        );

    \I__14449\ : CascadeMux
    port map (
            O => \N__64693\,
            I => \N__64657\
        );

    \I__14448\ : Span4Mux_v
    port map (
            O => \N__64690\,
            I => \N__64648\
        );

    \I__14447\ : Span4Mux_h
    port map (
            O => \N__64683\,
            I => \N__64648\
        );

    \I__14446\ : LocalMux
    port map (
            O => \N__64680\,
            I => \N__64648\
        );

    \I__14445\ : LocalMux
    port map (
            O => \N__64677\,
            I => \N__64648\
        );

    \I__14444\ : Span4Mux_h
    port map (
            O => \N__64674\,
            I => \N__64633\
        );

    \I__14443\ : LocalMux
    port map (
            O => \N__64671\,
            I => \N__64633\
        );

    \I__14442\ : Span4Mux_v
    port map (
            O => \N__64666\,
            I => \N__64625\
        );

    \I__14441\ : LocalMux
    port map (
            O => \N__64663\,
            I => \N__64625\
        );

    \I__14440\ : LocalMux
    port map (
            O => \N__64660\,
            I => \N__64625\
        );

    \I__14439\ : InMux
    port map (
            O => \N__64657\,
            I => \N__64622\
        );

    \I__14438\ : Span4Mux_v
    port map (
            O => \N__64648\,
            I => \N__64619\
        );

    \I__14437\ : CascadeMux
    port map (
            O => \N__64647\,
            I => \N__64616\
        );

    \I__14436\ : CascadeMux
    port map (
            O => \N__64646\,
            I => \N__64613\
        );

    \I__14435\ : CascadeMux
    port map (
            O => \N__64645\,
            I => \N__64609\
        );

    \I__14434\ : CascadeMux
    port map (
            O => \N__64644\,
            I => \N__64606\
        );

    \I__14433\ : CascadeMux
    port map (
            O => \N__64643\,
            I => \N__64603\
        );

    \I__14432\ : CascadeMux
    port map (
            O => \N__64642\,
            I => \N__64600\
        );

    \I__14431\ : CascadeMux
    port map (
            O => \N__64641\,
            I => \N__64596\
        );

    \I__14430\ : CascadeMux
    port map (
            O => \N__64640\,
            I => \N__64593\
        );

    \I__14429\ : CascadeMux
    port map (
            O => \N__64639\,
            I => \N__64589\
        );

    \I__14428\ : CascadeMux
    port map (
            O => \N__64638\,
            I => \N__64585\
        );

    \I__14427\ : Span4Mux_v
    port map (
            O => \N__64633\,
            I => \N__64582\
        );

    \I__14426\ : InMux
    port map (
            O => \N__64632\,
            I => \N__64579\
        );

    \I__14425\ : Span4Mux_h
    port map (
            O => \N__64625\,
            I => \N__64576\
        );

    \I__14424\ : LocalMux
    port map (
            O => \N__64622\,
            I => \N__64573\
        );

    \I__14423\ : Span4Mux_h
    port map (
            O => \N__64619\,
            I => \N__64570\
        );

    \I__14422\ : InMux
    port map (
            O => \N__64616\,
            I => \N__64565\
        );

    \I__14421\ : InMux
    port map (
            O => \N__64613\,
            I => \N__64565\
        );

    \I__14420\ : InMux
    port map (
            O => \N__64612\,
            I => \N__64556\
        );

    \I__14419\ : InMux
    port map (
            O => \N__64609\,
            I => \N__64556\
        );

    \I__14418\ : InMux
    port map (
            O => \N__64606\,
            I => \N__64556\
        );

    \I__14417\ : InMux
    port map (
            O => \N__64603\,
            I => \N__64556\
        );

    \I__14416\ : InMux
    port map (
            O => \N__64600\,
            I => \N__64549\
        );

    \I__14415\ : InMux
    port map (
            O => \N__64599\,
            I => \N__64549\
        );

    \I__14414\ : InMux
    port map (
            O => \N__64596\,
            I => \N__64549\
        );

    \I__14413\ : InMux
    port map (
            O => \N__64593\,
            I => \N__64538\
        );

    \I__14412\ : InMux
    port map (
            O => \N__64592\,
            I => \N__64538\
        );

    \I__14411\ : InMux
    port map (
            O => \N__64589\,
            I => \N__64538\
        );

    \I__14410\ : InMux
    port map (
            O => \N__64588\,
            I => \N__64538\
        );

    \I__14409\ : InMux
    port map (
            O => \N__64585\,
            I => \N__64538\
        );

    \I__14408\ : Sp12to4
    port map (
            O => \N__64582\,
            I => \N__64533\
        );

    \I__14407\ : LocalMux
    port map (
            O => \N__64579\,
            I => \N__64533\
        );

    \I__14406\ : Span4Mux_v
    port map (
            O => \N__64576\,
            I => \N__64528\
        );

    \I__14405\ : Span4Mux_h
    port map (
            O => \N__64573\,
            I => \N__64528\
        );

    \I__14404\ : Sp12to4
    port map (
            O => \N__64570\,
            I => \N__64519\
        );

    \I__14403\ : LocalMux
    port map (
            O => \N__64565\,
            I => \N__64519\
        );

    \I__14402\ : LocalMux
    port map (
            O => \N__64556\,
            I => \N__64519\
        );

    \I__14401\ : LocalMux
    port map (
            O => \N__64549\,
            I => \N__64519\
        );

    \I__14400\ : LocalMux
    port map (
            O => \N__64538\,
            I => \N__64516\
        );

    \I__14399\ : Odrv12
    port map (
            O => \N__64533\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0\
        );

    \I__14398\ : Odrv4
    port map (
            O => \N__64528\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0\
        );

    \I__14397\ : Odrv12
    port map (
            O => \N__64519\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0\
        );

    \I__14396\ : Odrv4
    port map (
            O => \N__64516\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0\
        );

    \I__14395\ : InMux
    port map (
            O => \N__64507\,
            I => \N__64504\
        );

    \I__14394\ : LocalMux
    port map (
            O => \N__64504\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n75\
        );

    \I__14393\ : CascadeMux
    port map (
            O => \N__64501\,
            I => \N__64498\
        );

    \I__14392\ : InMux
    port map (
            O => \N__64498\,
            I => \N__64493\
        );

    \I__14391\ : CascadeMux
    port map (
            O => \N__64497\,
            I => \N__64490\
        );

    \I__14390\ : CascadeMux
    port map (
            O => \N__64496\,
            I => \N__64485\
        );

    \I__14389\ : LocalMux
    port map (
            O => \N__64493\,
            I => \N__64482\
        );

    \I__14388\ : InMux
    port map (
            O => \N__64490\,
            I => \N__64479\
        );

    \I__14387\ : CascadeMux
    port map (
            O => \N__64489\,
            I => \N__64475\
        );

    \I__14386\ : CascadeMux
    port map (
            O => \N__64488\,
            I => \N__64472\
        );

    \I__14385\ : InMux
    port map (
            O => \N__64485\,
            I => \N__64467\
        );

    \I__14384\ : Span4Mux_h
    port map (
            O => \N__64482\,
            I => \N__64461\
        );

    \I__14383\ : LocalMux
    port map (
            O => \N__64479\,
            I => \N__64461\
        );

    \I__14382\ : InMux
    port map (
            O => \N__64478\,
            I => \N__64458\
        );

    \I__14381\ : InMux
    port map (
            O => \N__64475\,
            I => \N__64455\
        );

    \I__14380\ : InMux
    port map (
            O => \N__64472\,
            I => \N__64447\
        );

    \I__14379\ : InMux
    port map (
            O => \N__64471\,
            I => \N__64444\
        );

    \I__14378\ : CascadeMux
    port map (
            O => \N__64470\,
            I => \N__64441\
        );

    \I__14377\ : LocalMux
    port map (
            O => \N__64467\,
            I => \N__64434\
        );

    \I__14376\ : CascadeMux
    port map (
            O => \N__64466\,
            I => \N__64431\
        );

    \I__14375\ : Span4Mux_v
    port map (
            O => \N__64461\,
            I => \N__64426\
        );

    \I__14374\ : LocalMux
    port map (
            O => \N__64458\,
            I => \N__64426\
        );

    \I__14373\ : LocalMux
    port map (
            O => \N__64455\,
            I => \N__64423\
        );

    \I__14372\ : InMux
    port map (
            O => \N__64454\,
            I => \N__64420\
        );

    \I__14371\ : InMux
    port map (
            O => \N__64453\,
            I => \N__64417\
        );

    \I__14370\ : CascadeMux
    port map (
            O => \N__64452\,
            I => \N__64414\
        );

    \I__14369\ : CascadeMux
    port map (
            O => \N__64451\,
            I => \N__64411\
        );

    \I__14368\ : CascadeMux
    port map (
            O => \N__64450\,
            I => \N__64408\
        );

    \I__14367\ : LocalMux
    port map (
            O => \N__64447\,
            I => \N__64403\
        );

    \I__14366\ : LocalMux
    port map (
            O => \N__64444\,
            I => \N__64403\
        );

    \I__14365\ : InMux
    port map (
            O => \N__64441\,
            I => \N__64400\
        );

    \I__14364\ : InMux
    port map (
            O => \N__64440\,
            I => \N__64397\
        );

    \I__14363\ : CascadeMux
    port map (
            O => \N__64439\,
            I => \N__64393\
        );

    \I__14362\ : CascadeMux
    port map (
            O => \N__64438\,
            I => \N__64389\
        );

    \I__14361\ : CascadeMux
    port map (
            O => \N__64437\,
            I => \N__64385\
        );

    \I__14360\ : Span4Mux_v
    port map (
            O => \N__64434\,
            I => \N__64378\
        );

    \I__14359\ : InMux
    port map (
            O => \N__64431\,
            I => \N__64375\
        );

    \I__14358\ : Span4Mux_v
    port map (
            O => \N__64426\,
            I => \N__64368\
        );

    \I__14357\ : Span4Mux_v
    port map (
            O => \N__64423\,
            I => \N__64368\
        );

    \I__14356\ : LocalMux
    port map (
            O => \N__64420\,
            I => \N__64368\
        );

    \I__14355\ : LocalMux
    port map (
            O => \N__64417\,
            I => \N__64365\
        );

    \I__14354\ : InMux
    port map (
            O => \N__64414\,
            I => \N__64362\
        );

    \I__14353\ : InMux
    port map (
            O => \N__64411\,
            I => \N__64359\
        );

    \I__14352\ : InMux
    port map (
            O => \N__64408\,
            I => \N__64356\
        );

    \I__14351\ : Span4Mux_v
    port map (
            O => \N__64403\,
            I => \N__64349\
        );

    \I__14350\ : LocalMux
    port map (
            O => \N__64400\,
            I => \N__64349\
        );

    \I__14349\ : LocalMux
    port map (
            O => \N__64397\,
            I => \N__64349\
        );

    \I__14348\ : InMux
    port map (
            O => \N__64396\,
            I => \N__64336\
        );

    \I__14347\ : InMux
    port map (
            O => \N__64393\,
            I => \N__64336\
        );

    \I__14346\ : InMux
    port map (
            O => \N__64392\,
            I => \N__64336\
        );

    \I__14345\ : InMux
    port map (
            O => \N__64389\,
            I => \N__64336\
        );

    \I__14344\ : InMux
    port map (
            O => \N__64388\,
            I => \N__64336\
        );

    \I__14343\ : InMux
    port map (
            O => \N__64385\,
            I => \N__64336\
        );

    \I__14342\ : CascadeMux
    port map (
            O => \N__64384\,
            I => \N__64332\
        );

    \I__14341\ : CascadeMux
    port map (
            O => \N__64383\,
            I => \N__64328\
        );

    \I__14340\ : CascadeMux
    port map (
            O => \N__64382\,
            I => \N__64324\
        );

    \I__14339\ : CascadeMux
    port map (
            O => \N__64381\,
            I => \N__64320\
        );

    \I__14338\ : Span4Mux_h
    port map (
            O => \N__64378\,
            I => \N__64315\
        );

    \I__14337\ : LocalMux
    port map (
            O => \N__64375\,
            I => \N__64315\
        );

    \I__14336\ : Span4Mux_h
    port map (
            O => \N__64368\,
            I => \N__64308\
        );

    \I__14335\ : Span4Mux_h
    port map (
            O => \N__64365\,
            I => \N__64308\
        );

    \I__14334\ : LocalMux
    port map (
            O => \N__64362\,
            I => \N__64308\
        );

    \I__14333\ : LocalMux
    port map (
            O => \N__64359\,
            I => \N__64303\
        );

    \I__14332\ : LocalMux
    port map (
            O => \N__64356\,
            I => \N__64303\
        );

    \I__14331\ : Span4Mux_h
    port map (
            O => \N__64349\,
            I => \N__64298\
        );

    \I__14330\ : LocalMux
    port map (
            O => \N__64336\,
            I => \N__64298\
        );

    \I__14329\ : InMux
    port map (
            O => \N__64335\,
            I => \N__64281\
        );

    \I__14328\ : InMux
    port map (
            O => \N__64332\,
            I => \N__64281\
        );

    \I__14327\ : InMux
    port map (
            O => \N__64331\,
            I => \N__64281\
        );

    \I__14326\ : InMux
    port map (
            O => \N__64328\,
            I => \N__64281\
        );

    \I__14325\ : InMux
    port map (
            O => \N__64327\,
            I => \N__64281\
        );

    \I__14324\ : InMux
    port map (
            O => \N__64324\,
            I => \N__64281\
        );

    \I__14323\ : InMux
    port map (
            O => \N__64323\,
            I => \N__64281\
        );

    \I__14322\ : InMux
    port map (
            O => \N__64320\,
            I => \N__64281\
        );

    \I__14321\ : Span4Mux_v
    port map (
            O => \N__64315\,
            I => \N__64278\
        );

    \I__14320\ : Span4Mux_v
    port map (
            O => \N__64308\,
            I => \N__64275\
        );

    \I__14319\ : Span12Mux_h
    port map (
            O => \N__64303\,
            I => \N__64268\
        );

    \I__14318\ : Sp12to4
    port map (
            O => \N__64298\,
            I => \N__64268\
        );

    \I__14317\ : LocalMux
    port map (
            O => \N__64281\,
            I => \N__64268\
        );

    \I__14316\ : Odrv4
    port map (
            O => \N__64278\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n105\
        );

    \I__14315\ : Odrv4
    port map (
            O => \N__64275\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n105\
        );

    \I__14314\ : Odrv12
    port map (
            O => \N__64268\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n105\
        );

    \I__14313\ : InMux
    port map (
            O => \N__64261\,
            I => \N__64258\
        );

    \I__14312\ : LocalMux
    port map (
            O => \N__64258\,
            I => \N__64255\
        );

    \I__14311\ : Odrv12
    port map (
            O => \N__64255\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n121\
        );

    \I__14310\ : InMux
    port map (
            O => \N__64252\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18264\
        );

    \I__14309\ : InMux
    port map (
            O => \N__64249\,
            I => \N__64246\
        );

    \I__14308\ : LocalMux
    port map (
            O => \N__64246\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n124\
        );

    \I__14307\ : CascadeMux
    port map (
            O => \N__64243\,
            I => \N__64227\
        );

    \I__14306\ : CascadeMux
    port map (
            O => \N__64242\,
            I => \N__64224\
        );

    \I__14305\ : CascadeMux
    port map (
            O => \N__64241\,
            I => \N__64221\
        );

    \I__14304\ : CascadeMux
    port map (
            O => \N__64240\,
            I => \N__64216\
        );

    \I__14303\ : CascadeMux
    port map (
            O => \N__64239\,
            I => \N__64212\
        );

    \I__14302\ : CascadeMux
    port map (
            O => \N__64238\,
            I => \N__64208\
        );

    \I__14301\ : CascadeMux
    port map (
            O => \N__64237\,
            I => \N__64204\
        );

    \I__14300\ : CascadeMux
    port map (
            O => \N__64236\,
            I => \N__64201\
        );

    \I__14299\ : CascadeMux
    port map (
            O => \N__64235\,
            I => \N__64197\
        );

    \I__14298\ : CascadeMux
    port map (
            O => \N__64234\,
            I => \N__64193\
        );

    \I__14297\ : CascadeMux
    port map (
            O => \N__64233\,
            I => \N__64189\
        );

    \I__14296\ : CascadeMux
    port map (
            O => \N__64232\,
            I => \N__64186\
        );

    \I__14295\ : CascadeMux
    port map (
            O => \N__64231\,
            I => \N__64183\
        );

    \I__14294\ : CascadeMux
    port map (
            O => \N__64230\,
            I => \N__64179\
        );

    \I__14293\ : InMux
    port map (
            O => \N__64227\,
            I => \N__64175\
        );

    \I__14292\ : InMux
    port map (
            O => \N__64224\,
            I => \N__64172\
        );

    \I__14291\ : InMux
    port map (
            O => \N__64221\,
            I => \N__64169\
        );

    \I__14290\ : CascadeMux
    port map (
            O => \N__64220\,
            I => \N__64166\
        );

    \I__14289\ : InMux
    port map (
            O => \N__64219\,
            I => \N__64149\
        );

    \I__14288\ : InMux
    port map (
            O => \N__64216\,
            I => \N__64149\
        );

    \I__14287\ : InMux
    port map (
            O => \N__64215\,
            I => \N__64149\
        );

    \I__14286\ : InMux
    port map (
            O => \N__64212\,
            I => \N__64149\
        );

    \I__14285\ : InMux
    port map (
            O => \N__64211\,
            I => \N__64149\
        );

    \I__14284\ : InMux
    port map (
            O => \N__64208\,
            I => \N__64149\
        );

    \I__14283\ : InMux
    port map (
            O => \N__64207\,
            I => \N__64149\
        );

    \I__14282\ : InMux
    port map (
            O => \N__64204\,
            I => \N__64149\
        );

    \I__14281\ : InMux
    port map (
            O => \N__64201\,
            I => \N__64146\
        );

    \I__14280\ : InMux
    port map (
            O => \N__64200\,
            I => \N__64133\
        );

    \I__14279\ : InMux
    port map (
            O => \N__64197\,
            I => \N__64133\
        );

    \I__14278\ : InMux
    port map (
            O => \N__64196\,
            I => \N__64133\
        );

    \I__14277\ : InMux
    port map (
            O => \N__64193\,
            I => \N__64133\
        );

    \I__14276\ : InMux
    port map (
            O => \N__64192\,
            I => \N__64133\
        );

    \I__14275\ : InMux
    port map (
            O => \N__64189\,
            I => \N__64133\
        );

    \I__14274\ : InMux
    port map (
            O => \N__64186\,
            I => \N__64129\
        );

    \I__14273\ : InMux
    port map (
            O => \N__64183\,
            I => \N__64126\
        );

    \I__14272\ : InMux
    port map (
            O => \N__64182\,
            I => \N__64123\
        );

    \I__14271\ : InMux
    port map (
            O => \N__64179\,
            I => \N__64120\
        );

    \I__14270\ : CascadeMux
    port map (
            O => \N__64178\,
            I => \N__64117\
        );

    \I__14269\ : LocalMux
    port map (
            O => \N__64175\,
            I => \N__64112\
        );

    \I__14268\ : LocalMux
    port map (
            O => \N__64172\,
            I => \N__64112\
        );

    \I__14267\ : LocalMux
    port map (
            O => \N__64169\,
            I => \N__64108\
        );

    \I__14266\ : InMux
    port map (
            O => \N__64166\,
            I => \N__64105\
        );

    \I__14265\ : LocalMux
    port map (
            O => \N__64149\,
            I => \N__64102\
        );

    \I__14264\ : LocalMux
    port map (
            O => \N__64146\,
            I => \N__64098\
        );

    \I__14263\ : LocalMux
    port map (
            O => \N__64133\,
            I => \N__64095\
        );

    \I__14262\ : InMux
    port map (
            O => \N__64132\,
            I => \N__64092\
        );

    \I__14261\ : LocalMux
    port map (
            O => \N__64129\,
            I => \N__64081\
        );

    \I__14260\ : LocalMux
    port map (
            O => \N__64126\,
            I => \N__64081\
        );

    \I__14259\ : LocalMux
    port map (
            O => \N__64123\,
            I => \N__64081\
        );

    \I__14258\ : LocalMux
    port map (
            O => \N__64120\,
            I => \N__64081\
        );

    \I__14257\ : InMux
    port map (
            O => \N__64117\,
            I => \N__64078\
        );

    \I__14256\ : Span4Mux_v
    port map (
            O => \N__64112\,
            I => \N__64075\
        );

    \I__14255\ : InMux
    port map (
            O => \N__64111\,
            I => \N__64072\
        );

    \I__14254\ : Span4Mux_h
    port map (
            O => \N__64108\,
            I => \N__64067\
        );

    \I__14253\ : LocalMux
    port map (
            O => \N__64105\,
            I => \N__64067\
        );

    \I__14252\ : Span4Mux_v
    port map (
            O => \N__64102\,
            I => \N__64064\
        );

    \I__14251\ : InMux
    port map (
            O => \N__64101\,
            I => \N__64061\
        );

    \I__14250\ : Span4Mux_v
    port map (
            O => \N__64098\,
            I => \N__64054\
        );

    \I__14249\ : Span4Mux_h
    port map (
            O => \N__64095\,
            I => \N__64054\
        );

    \I__14248\ : LocalMux
    port map (
            O => \N__64092\,
            I => \N__64054\
        );

    \I__14247\ : InMux
    port map (
            O => \N__64091\,
            I => \N__64051\
        );

    \I__14246\ : CascadeMux
    port map (
            O => \N__64090\,
            I => \N__64048\
        );

    \I__14245\ : Span4Mux_v
    port map (
            O => \N__64081\,
            I => \N__64043\
        );

    \I__14244\ : LocalMux
    port map (
            O => \N__64078\,
            I => \N__64043\
        );

    \I__14243\ : Span4Mux_h
    port map (
            O => \N__64075\,
            I => \N__64038\
        );

    \I__14242\ : LocalMux
    port map (
            O => \N__64072\,
            I => \N__64038\
        );

    \I__14241\ : Span4Mux_v
    port map (
            O => \N__64067\,
            I => \N__64031\
        );

    \I__14240\ : Span4Mux_h
    port map (
            O => \N__64064\,
            I => \N__64031\
        );

    \I__14239\ : LocalMux
    port map (
            O => \N__64061\,
            I => \N__64031\
        );

    \I__14238\ : Span4Mux_h
    port map (
            O => \N__64054\,
            I => \N__64026\
        );

    \I__14237\ : LocalMux
    port map (
            O => \N__64051\,
            I => \N__64026\
        );

    \I__14236\ : InMux
    port map (
            O => \N__64048\,
            I => \N__64023\
        );

    \I__14235\ : Span4Mux_v
    port map (
            O => \N__64043\,
            I => \N__64020\
        );

    \I__14234\ : Span4Mux_v
    port map (
            O => \N__64038\,
            I => \N__64017\
        );

    \I__14233\ : Span4Mux_h
    port map (
            O => \N__64031\,
            I => \N__64014\
        );

    \I__14232\ : Sp12to4
    port map (
            O => \N__64026\,
            I => \N__64009\
        );

    \I__14231\ : LocalMux
    port map (
            O => \N__64023\,
            I => \N__64009\
        );

    \I__14230\ : Odrv4
    port map (
            O => \N__64020\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n108\
        );

    \I__14229\ : Odrv4
    port map (
            O => \N__64017\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n108\
        );

    \I__14228\ : Odrv4
    port map (
            O => \N__64014\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n108\
        );

    \I__14227\ : Odrv12
    port map (
            O => \N__64009\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n108\
        );

    \I__14226\ : InMux
    port map (
            O => \N__64000\,
            I => \N__63997\
        );

    \I__14225\ : LocalMux
    port map (
            O => \N__63997\,
            I => \N__63994\
        );

    \I__14224\ : Odrv4
    port map (
            O => \N__63994\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n170\
        );

    \I__14223\ : InMux
    port map (
            O => \N__63991\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18265\
        );

    \I__14222\ : InMux
    port map (
            O => \N__63988\,
            I => \N__63985\
        );

    \I__14221\ : LocalMux
    port map (
            O => \N__63985\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n173\
        );

    \I__14220\ : CascadeMux
    port map (
            O => \N__63982\,
            I => \N__63976\
        );

    \I__14219\ : CascadeMux
    port map (
            O => \N__63981\,
            I => \N__63971\
        );

    \I__14218\ : CascadeMux
    port map (
            O => \N__63980\,
            I => \N__63968\
        );

    \I__14217\ : CascadeMux
    port map (
            O => \N__63979\,
            I => \N__63964\
        );

    \I__14216\ : InMux
    port map (
            O => \N__63976\,
            I => \N__63959\
        );

    \I__14215\ : InMux
    port map (
            O => \N__63975\,
            I => \N__63956\
        );

    \I__14214\ : CascadeMux
    port map (
            O => \N__63974\,
            I => \N__63952\
        );

    \I__14213\ : InMux
    port map (
            O => \N__63971\,
            I => \N__63943\
        );

    \I__14212\ : InMux
    port map (
            O => \N__63968\,
            I => \N__63940\
        );

    \I__14211\ : CascadeMux
    port map (
            O => \N__63967\,
            I => \N__63937\
        );

    \I__14210\ : InMux
    port map (
            O => \N__63964\,
            I => \N__63933\
        );

    \I__14209\ : CascadeMux
    port map (
            O => \N__63963\,
            I => \N__63930\
        );

    \I__14208\ : CascadeMux
    port map (
            O => \N__63962\,
            I => \N__63926\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__63959\,
            I => \N__63921\
        );

    \I__14206\ : LocalMux
    port map (
            O => \N__63956\,
            I => \N__63921\
        );

    \I__14205\ : CascadeMux
    port map (
            O => \N__63955\,
            I => \N__63918\
        );

    \I__14204\ : InMux
    port map (
            O => \N__63952\,
            I => \N__63915\
        );

    \I__14203\ : CascadeMux
    port map (
            O => \N__63951\,
            I => \N__63912\
        );

    \I__14202\ : CascadeMux
    port map (
            O => \N__63950\,
            I => \N__63909\
        );

    \I__14201\ : CascadeMux
    port map (
            O => \N__63949\,
            I => \N__63906\
        );

    \I__14200\ : CascadeMux
    port map (
            O => \N__63948\,
            I => \N__63903\
        );

    \I__14199\ : CascadeMux
    port map (
            O => \N__63947\,
            I => \N__63900\
        );

    \I__14198\ : CascadeMux
    port map (
            O => \N__63946\,
            I => \N__63897\
        );

    \I__14197\ : LocalMux
    port map (
            O => \N__63943\,
            I => \N__63885\
        );

    \I__14196\ : LocalMux
    port map (
            O => \N__63940\,
            I => \N__63882\
        );

    \I__14195\ : InMux
    port map (
            O => \N__63937\,
            I => \N__63879\
        );

    \I__14194\ : CascadeMux
    port map (
            O => \N__63936\,
            I => \N__63876\
        );

    \I__14193\ : LocalMux
    port map (
            O => \N__63933\,
            I => \N__63872\
        );

    \I__14192\ : InMux
    port map (
            O => \N__63930\,
            I => \N__63869\
        );

    \I__14191\ : CascadeMux
    port map (
            O => \N__63929\,
            I => \N__63866\
        );

    \I__14190\ : InMux
    port map (
            O => \N__63926\,
            I => \N__63863\
        );

    \I__14189\ : Span4Mux_h
    port map (
            O => \N__63921\,
            I => \N__63859\
        );

    \I__14188\ : InMux
    port map (
            O => \N__63918\,
            I => \N__63856\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__63915\,
            I => \N__63853\
        );

    \I__14186\ : InMux
    port map (
            O => \N__63912\,
            I => \N__63846\
        );

    \I__14185\ : InMux
    port map (
            O => \N__63909\,
            I => \N__63846\
        );

    \I__14184\ : InMux
    port map (
            O => \N__63906\,
            I => \N__63846\
        );

    \I__14183\ : InMux
    port map (
            O => \N__63903\,
            I => \N__63839\
        );

    \I__14182\ : InMux
    port map (
            O => \N__63900\,
            I => \N__63839\
        );

    \I__14181\ : InMux
    port map (
            O => \N__63897\,
            I => \N__63839\
        );

    \I__14180\ : CascadeMux
    port map (
            O => \N__63896\,
            I => \N__63836\
        );

    \I__14179\ : CascadeMux
    port map (
            O => \N__63895\,
            I => \N__63833\
        );

    \I__14178\ : CascadeMux
    port map (
            O => \N__63894\,
            I => \N__63830\
        );

    \I__14177\ : CascadeMux
    port map (
            O => \N__63893\,
            I => \N__63827\
        );

    \I__14176\ : CascadeMux
    port map (
            O => \N__63892\,
            I => \N__63824\
        );

    \I__14175\ : CascadeMux
    port map (
            O => \N__63891\,
            I => \N__63821\
        );

    \I__14174\ : CascadeMux
    port map (
            O => \N__63890\,
            I => \N__63818\
        );

    \I__14173\ : CascadeMux
    port map (
            O => \N__63889\,
            I => \N__63815\
        );

    \I__14172\ : CascadeMux
    port map (
            O => \N__63888\,
            I => \N__63812\
        );

    \I__14171\ : Span4Mux_v
    port map (
            O => \N__63885\,
            I => \N__63805\
        );

    \I__14170\ : Span4Mux_h
    port map (
            O => \N__63882\,
            I => \N__63805\
        );

    \I__14169\ : LocalMux
    port map (
            O => \N__63879\,
            I => \N__63805\
        );

    \I__14168\ : InMux
    port map (
            O => \N__63876\,
            I => \N__63802\
        );

    \I__14167\ : InMux
    port map (
            O => \N__63875\,
            I => \N__63799\
        );

    \I__14166\ : Span4Mux_v
    port map (
            O => \N__63872\,
            I => \N__63794\
        );

    \I__14165\ : LocalMux
    port map (
            O => \N__63869\,
            I => \N__63794\
        );

    \I__14164\ : InMux
    port map (
            O => \N__63866\,
            I => \N__63791\
        );

    \I__14163\ : LocalMux
    port map (
            O => \N__63863\,
            I => \N__63788\
        );

    \I__14162\ : InMux
    port map (
            O => \N__63862\,
            I => \N__63785\
        );

    \I__14161\ : Span4Mux_v
    port map (
            O => \N__63859\,
            I => \N__63780\
        );

    \I__14160\ : LocalMux
    port map (
            O => \N__63856\,
            I => \N__63780\
        );

    \I__14159\ : Span4Mux_v
    port map (
            O => \N__63853\,
            I => \N__63777\
        );

    \I__14158\ : LocalMux
    port map (
            O => \N__63846\,
            I => \N__63772\
        );

    \I__14157\ : LocalMux
    port map (
            O => \N__63839\,
            I => \N__63772\
        );

    \I__14156\ : InMux
    port map (
            O => \N__63836\,
            I => \N__63763\
        );

    \I__14155\ : InMux
    port map (
            O => \N__63833\,
            I => \N__63763\
        );

    \I__14154\ : InMux
    port map (
            O => \N__63830\,
            I => \N__63763\
        );

    \I__14153\ : InMux
    port map (
            O => \N__63827\,
            I => \N__63763\
        );

    \I__14152\ : InMux
    port map (
            O => \N__63824\,
            I => \N__63754\
        );

    \I__14151\ : InMux
    port map (
            O => \N__63821\,
            I => \N__63754\
        );

    \I__14150\ : InMux
    port map (
            O => \N__63818\,
            I => \N__63754\
        );

    \I__14149\ : InMux
    port map (
            O => \N__63815\,
            I => \N__63754\
        );

    \I__14148\ : InMux
    port map (
            O => \N__63812\,
            I => \N__63751\
        );

    \I__14147\ : Span4Mux_v
    port map (
            O => \N__63805\,
            I => \N__63746\
        );

    \I__14146\ : LocalMux
    port map (
            O => \N__63802\,
            I => \N__63746\
        );

    \I__14145\ : LocalMux
    port map (
            O => \N__63799\,
            I => \N__63739\
        );

    \I__14144\ : Span4Mux_h
    port map (
            O => \N__63794\,
            I => \N__63739\
        );

    \I__14143\ : LocalMux
    port map (
            O => \N__63791\,
            I => \N__63739\
        );

    \I__14142\ : Span4Mux_h
    port map (
            O => \N__63788\,
            I => \N__63734\
        );

    \I__14141\ : LocalMux
    port map (
            O => \N__63785\,
            I => \N__63734\
        );

    \I__14140\ : Span4Mux_h
    port map (
            O => \N__63780\,
            I => \N__63731\
        );

    \I__14139\ : Sp12to4
    port map (
            O => \N__63777\,
            I => \N__63720\
        );

    \I__14138\ : Span12Mux_s9_v
    port map (
            O => \N__63772\,
            I => \N__63720\
        );

    \I__14137\ : LocalMux
    port map (
            O => \N__63763\,
            I => \N__63720\
        );

    \I__14136\ : LocalMux
    port map (
            O => \N__63754\,
            I => \N__63720\
        );

    \I__14135\ : LocalMux
    port map (
            O => \N__63751\,
            I => \N__63720\
        );

    \I__14134\ : Span4Mux_h
    port map (
            O => \N__63746\,
            I => \N__63715\
        );

    \I__14133\ : Span4Mux_h
    port map (
            O => \N__63739\,
            I => \N__63715\
        );

    \I__14132\ : Odrv4
    port map (
            O => \N__63734\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n111\
        );

    \I__14131\ : Odrv4
    port map (
            O => \N__63731\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n111\
        );

    \I__14130\ : Odrv12
    port map (
            O => \N__63720\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n111\
        );

    \I__14129\ : Odrv4
    port map (
            O => \N__63715\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n111\
        );

    \I__14128\ : InMux
    port map (
            O => \N__63706\,
            I => \N__63703\
        );

    \I__14127\ : LocalMux
    port map (
            O => \N__63703\,
            I => \N__63700\
        );

    \I__14126\ : Odrv12
    port map (
            O => \N__63700\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n219\
        );

    \I__14125\ : InMux
    port map (
            O => \N__63697\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18266\
        );

    \I__14124\ : InMux
    port map (
            O => \N__63694\,
            I => \N__63691\
        );

    \I__14123\ : LocalMux
    port map (
            O => \N__63691\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n222\
        );

    \I__14122\ : CascadeMux
    port map (
            O => \N__63688\,
            I => \N__63683\
        );

    \I__14121\ : CascadeMux
    port map (
            O => \N__63687\,
            I => \N__63679\
        );

    \I__14120\ : CascadeMux
    port map (
            O => \N__63686\,
            I => \N__63676\
        );

    \I__14119\ : InMux
    port map (
            O => \N__63683\,
            I => \N__63673\
        );

    \I__14118\ : CascadeMux
    port map (
            O => \N__63682\,
            I => \N__63670\
        );

    \I__14117\ : InMux
    port map (
            O => \N__63679\,
            I => \N__63665\
        );

    \I__14116\ : InMux
    port map (
            O => \N__63676\,
            I => \N__63662\
        );

    \I__14115\ : LocalMux
    port map (
            O => \N__63673\,
            I => \N__63659\
        );

    \I__14114\ : InMux
    port map (
            O => \N__63670\,
            I => \N__63656\
        );

    \I__14113\ : CascadeMux
    port map (
            O => \N__63669\,
            I => \N__63652\
        );

    \I__14112\ : CascadeMux
    port map (
            O => \N__63668\,
            I => \N__63649\
        );

    \I__14111\ : LocalMux
    port map (
            O => \N__63665\,
            I => \N__63644\
        );

    \I__14110\ : LocalMux
    port map (
            O => \N__63662\,
            I => \N__63641\
        );

    \I__14109\ : Span4Mux_v
    port map (
            O => \N__63659\,
            I => \N__63636\
        );

    \I__14108\ : LocalMux
    port map (
            O => \N__63656\,
            I => \N__63636\
        );

    \I__14107\ : CascadeMux
    port map (
            O => \N__63655\,
            I => \N__63627\
        );

    \I__14106\ : InMux
    port map (
            O => \N__63652\,
            I => \N__63619\
        );

    \I__14105\ : InMux
    port map (
            O => \N__63649\,
            I => \N__63616\
        );

    \I__14104\ : CascadeMux
    port map (
            O => \N__63648\,
            I => \N__63613\
        );

    \I__14103\ : CascadeMux
    port map (
            O => \N__63647\,
            I => \N__63610\
        );

    \I__14102\ : Span4Mux_v
    port map (
            O => \N__63644\,
            I => \N__63600\
        );

    \I__14101\ : Span4Mux_v
    port map (
            O => \N__63641\,
            I => \N__63600\
        );

    \I__14100\ : Span4Mux_v
    port map (
            O => \N__63636\,
            I => \N__63600\
        );

    \I__14099\ : CascadeMux
    port map (
            O => \N__63635\,
            I => \N__63596\
        );

    \I__14098\ : CascadeMux
    port map (
            O => \N__63634\,
            I => \N__63592\
        );

    \I__14097\ : CascadeMux
    port map (
            O => \N__63633\,
            I => \N__63588\
        );

    \I__14096\ : CascadeMux
    port map (
            O => \N__63632\,
            I => \N__63584\
        );

    \I__14095\ : CascadeMux
    port map (
            O => \N__63631\,
            I => \N__63581\
        );

    \I__14094\ : InMux
    port map (
            O => \N__63630\,
            I => \N__63578\
        );

    \I__14093\ : InMux
    port map (
            O => \N__63627\,
            I => \N__63575\
        );

    \I__14092\ : CascadeMux
    port map (
            O => \N__63626\,
            I => \N__63572\
        );

    \I__14091\ : CascadeMux
    port map (
            O => \N__63625\,
            I => \N__63569\
        );

    \I__14090\ : CascadeMux
    port map (
            O => \N__63624\,
            I => \N__63566\
        );

    \I__14089\ : CascadeMux
    port map (
            O => \N__63623\,
            I => \N__63562\
        );

    \I__14088\ : CascadeMux
    port map (
            O => \N__63622\,
            I => \N__63558\
        );

    \I__14087\ : LocalMux
    port map (
            O => \N__63619\,
            I => \N__63553\
        );

    \I__14086\ : LocalMux
    port map (
            O => \N__63616\,
            I => \N__63553\
        );

    \I__14085\ : InMux
    port map (
            O => \N__63613\,
            I => \N__63550\
        );

    \I__14084\ : InMux
    port map (
            O => \N__63610\,
            I => \N__63547\
        );

    \I__14083\ : CascadeMux
    port map (
            O => \N__63609\,
            I => \N__63544\
        );

    \I__14082\ : CascadeMux
    port map (
            O => \N__63608\,
            I => \N__63541\
        );

    \I__14081\ : InMux
    port map (
            O => \N__63607\,
            I => \N__63538\
        );

    \I__14080\ : Span4Mux_h
    port map (
            O => \N__63600\,
            I => \N__63535\
        );

    \I__14079\ : InMux
    port map (
            O => \N__63599\,
            I => \N__63518\
        );

    \I__14078\ : InMux
    port map (
            O => \N__63596\,
            I => \N__63518\
        );

    \I__14077\ : InMux
    port map (
            O => \N__63595\,
            I => \N__63518\
        );

    \I__14076\ : InMux
    port map (
            O => \N__63592\,
            I => \N__63518\
        );

    \I__14075\ : InMux
    port map (
            O => \N__63591\,
            I => \N__63518\
        );

    \I__14074\ : InMux
    port map (
            O => \N__63588\,
            I => \N__63518\
        );

    \I__14073\ : InMux
    port map (
            O => \N__63587\,
            I => \N__63518\
        );

    \I__14072\ : InMux
    port map (
            O => \N__63584\,
            I => \N__63518\
        );

    \I__14071\ : InMux
    port map (
            O => \N__63581\,
            I => \N__63515\
        );

    \I__14070\ : LocalMux
    port map (
            O => \N__63578\,
            I => \N__63510\
        );

    \I__14069\ : LocalMux
    port map (
            O => \N__63575\,
            I => \N__63510\
        );

    \I__14068\ : InMux
    port map (
            O => \N__63572\,
            I => \N__63507\
        );

    \I__14067\ : InMux
    port map (
            O => \N__63569\,
            I => \N__63504\
        );

    \I__14066\ : InMux
    port map (
            O => \N__63566\,
            I => \N__63493\
        );

    \I__14065\ : InMux
    port map (
            O => \N__63565\,
            I => \N__63493\
        );

    \I__14064\ : InMux
    port map (
            O => \N__63562\,
            I => \N__63493\
        );

    \I__14063\ : InMux
    port map (
            O => \N__63561\,
            I => \N__63493\
        );

    \I__14062\ : InMux
    port map (
            O => \N__63558\,
            I => \N__63493\
        );

    \I__14061\ : Span4Mux_v
    port map (
            O => \N__63553\,
            I => \N__63488\
        );

    \I__14060\ : LocalMux
    port map (
            O => \N__63550\,
            I => \N__63488\
        );

    \I__14059\ : LocalMux
    port map (
            O => \N__63547\,
            I => \N__63485\
        );

    \I__14058\ : InMux
    port map (
            O => \N__63544\,
            I => \N__63482\
        );

    \I__14057\ : InMux
    port map (
            O => \N__63541\,
            I => \N__63479\
        );

    \I__14056\ : LocalMux
    port map (
            O => \N__63538\,
            I => \N__63472\
        );

    \I__14055\ : Sp12to4
    port map (
            O => \N__63535\,
            I => \N__63472\
        );

    \I__14054\ : LocalMux
    port map (
            O => \N__63518\,
            I => \N__63472\
        );

    \I__14053\ : LocalMux
    port map (
            O => \N__63515\,
            I => \N__63469\
        );

    \I__14052\ : Span4Mux_h
    port map (
            O => \N__63510\,
            I => \N__63464\
        );

    \I__14051\ : LocalMux
    port map (
            O => \N__63507\,
            I => \N__63464\
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__63504\,
            I => \N__63457\
        );

    \I__14049\ : LocalMux
    port map (
            O => \N__63493\,
            I => \N__63457\
        );

    \I__14048\ : Span4Mux_h
    port map (
            O => \N__63488\,
            I => \N__63457\
        );

    \I__14047\ : Span4Mux_h
    port map (
            O => \N__63485\,
            I => \N__63454\
        );

    \I__14046\ : LocalMux
    port map (
            O => \N__63482\,
            I => \N__63451\
        );

    \I__14045\ : LocalMux
    port map (
            O => \N__63479\,
            I => \N__63448\
        );

    \I__14044\ : Span12Mux_h
    port map (
            O => \N__63472\,
            I => \N__63443\
        );

    \I__14043\ : Span12Mux_h
    port map (
            O => \N__63469\,
            I => \N__63443\
        );

    \I__14042\ : Span4Mux_v
    port map (
            O => \N__63464\,
            I => \N__63438\
        );

    \I__14041\ : Span4Mux_h
    port map (
            O => \N__63457\,
            I => \N__63438\
        );

    \I__14040\ : Span4Mux_v
    port map (
            O => \N__63454\,
            I => \N__63433\
        );

    \I__14039\ : Span4Mux_h
    port map (
            O => \N__63451\,
            I => \N__63433\
        );

    \I__14038\ : Odrv12
    port map (
            O => \N__63448\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n114\
        );

    \I__14037\ : Odrv12
    port map (
            O => \N__63443\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n114\
        );

    \I__14036\ : Odrv4
    port map (
            O => \N__63438\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n114\
        );

    \I__14035\ : Odrv4
    port map (
            O => \N__63433\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n114\
        );

    \I__14034\ : InMux
    port map (
            O => \N__63424\,
            I => \N__63421\
        );

    \I__14033\ : LocalMux
    port map (
            O => \N__63421\,
            I => \N__63418\
        );

    \I__14032\ : Odrv4
    port map (
            O => \N__63418\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n268\
        );

    \I__14031\ : InMux
    port map (
            O => \N__63415\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18267\
        );

    \I__14030\ : InMux
    port map (
            O => \N__63412\,
            I => \N__63409\
        );

    \I__14029\ : LocalMux
    port map (
            O => \N__63409\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n271\
        );

    \I__14028\ : CascadeMux
    port map (
            O => \N__63406\,
            I => \N__63402\
        );

    \I__14027\ : CascadeMux
    port map (
            O => \N__63405\,
            I => \N__63396\
        );

    \I__14026\ : InMux
    port map (
            O => \N__63402\,
            I => \N__63393\
        );

    \I__14025\ : CascadeMux
    port map (
            O => \N__63401\,
            I => \N__63390\
        );

    \I__14024\ : CascadeMux
    port map (
            O => \N__63400\,
            I => \N__63386\
        );

    \I__14023\ : CascadeMux
    port map (
            O => \N__63399\,
            I => \N__63379\
        );

    \I__14022\ : InMux
    port map (
            O => \N__63396\,
            I => \N__63374\
        );

    \I__14021\ : LocalMux
    port map (
            O => \N__63393\,
            I => \N__63371\
        );

    \I__14020\ : InMux
    port map (
            O => \N__63390\,
            I => \N__63368\
        );

    \I__14019\ : CascadeMux
    port map (
            O => \N__63389\,
            I => \N__63365\
        );

    \I__14018\ : InMux
    port map (
            O => \N__63386\,
            I => \N__63362\
        );

    \I__14017\ : CascadeMux
    port map (
            O => \N__63385\,
            I => \N__63355\
        );

    \I__14016\ : CascadeMux
    port map (
            O => \N__63384\,
            I => \N__63352\
        );

    \I__14015\ : CascadeMux
    port map (
            O => \N__63383\,
            I => \N__63349\
        );

    \I__14014\ : CascadeMux
    port map (
            O => \N__63382\,
            I => \N__63346\
        );

    \I__14013\ : InMux
    port map (
            O => \N__63379\,
            I => \N__63343\
        );

    \I__14012\ : CascadeMux
    port map (
            O => \N__63378\,
            I => \N__63340\
        );

    \I__14011\ : CascadeMux
    port map (
            O => \N__63377\,
            I => \N__63337\
        );

    \I__14010\ : LocalMux
    port map (
            O => \N__63374\,
            I => \N__63329\
        );

    \I__14009\ : Span4Mux_v
    port map (
            O => \N__63371\,
            I => \N__63329\
        );

    \I__14008\ : LocalMux
    port map (
            O => \N__63368\,
            I => \N__63329\
        );

    \I__14007\ : InMux
    port map (
            O => \N__63365\,
            I => \N__63326\
        );

    \I__14006\ : LocalMux
    port map (
            O => \N__63362\,
            I => \N__63323\
        );

    \I__14005\ : CascadeMux
    port map (
            O => \N__63361\,
            I => \N__63320\
        );

    \I__14004\ : CascadeMux
    port map (
            O => \N__63360\,
            I => \N__63316\
        );

    \I__14003\ : CascadeMux
    port map (
            O => \N__63359\,
            I => \N__63312\
        );

    \I__14002\ : CascadeMux
    port map (
            O => \N__63358\,
            I => \N__63308\
        );

    \I__14001\ : InMux
    port map (
            O => \N__63355\,
            I => \N__63305\
        );

    \I__14000\ : InMux
    port map (
            O => \N__63352\,
            I => \N__63302\
        );

    \I__13999\ : InMux
    port map (
            O => \N__63349\,
            I => \N__63299\
        );

    \I__13998\ : InMux
    port map (
            O => \N__63346\,
            I => \N__63296\
        );

    \I__13997\ : LocalMux
    port map (
            O => \N__63343\,
            I => \N__63293\
        );

    \I__13996\ : InMux
    port map (
            O => \N__63340\,
            I => \N__63290\
        );

    \I__13995\ : InMux
    port map (
            O => \N__63337\,
            I => \N__63287\
        );

    \I__13994\ : CascadeMux
    port map (
            O => \N__63336\,
            I => \N__63281\
        );

    \I__13993\ : Span4Mux_h
    port map (
            O => \N__63329\,
            I => \N__63274\
        );

    \I__13992\ : LocalMux
    port map (
            O => \N__63326\,
            I => \N__63274\
        );

    \I__13991\ : Span4Mux_h
    port map (
            O => \N__63323\,
            I => \N__63271\
        );

    \I__13990\ : InMux
    port map (
            O => \N__63320\,
            I => \N__63268\
        );

    \I__13989\ : InMux
    port map (
            O => \N__63319\,
            I => \N__63255\
        );

    \I__13988\ : InMux
    port map (
            O => \N__63316\,
            I => \N__63255\
        );

    \I__13987\ : InMux
    port map (
            O => \N__63315\,
            I => \N__63255\
        );

    \I__13986\ : InMux
    port map (
            O => \N__63312\,
            I => \N__63255\
        );

    \I__13985\ : InMux
    port map (
            O => \N__63311\,
            I => \N__63255\
        );

    \I__13984\ : InMux
    port map (
            O => \N__63308\,
            I => \N__63255\
        );

    \I__13983\ : LocalMux
    port map (
            O => \N__63305\,
            I => \N__63252\
        );

    \I__13982\ : LocalMux
    port map (
            O => \N__63302\,
            I => \N__63247\
        );

    \I__13981\ : LocalMux
    port map (
            O => \N__63299\,
            I => \N__63247\
        );

    \I__13980\ : LocalMux
    port map (
            O => \N__63296\,
            I => \N__63238\
        );

    \I__13979\ : Span4Mux_h
    port map (
            O => \N__63293\,
            I => \N__63238\
        );

    \I__13978\ : LocalMux
    port map (
            O => \N__63290\,
            I => \N__63238\
        );

    \I__13977\ : LocalMux
    port map (
            O => \N__63287\,
            I => \N__63238\
        );

    \I__13976\ : CascadeMux
    port map (
            O => \N__63286\,
            I => \N__63234\
        );

    \I__13975\ : CascadeMux
    port map (
            O => \N__63285\,
            I => \N__63230\
        );

    \I__13974\ : CascadeMux
    port map (
            O => \N__63284\,
            I => \N__63226\
        );

    \I__13973\ : InMux
    port map (
            O => \N__63281\,
            I => \N__63221\
        );

    \I__13972\ : InMux
    port map (
            O => \N__63280\,
            I => \N__63221\
        );

    \I__13971\ : CascadeMux
    port map (
            O => \N__63279\,
            I => \N__63218\
        );

    \I__13970\ : Span4Mux_h
    port map (
            O => \N__63274\,
            I => \N__63215\
        );

    \I__13969\ : Span4Mux_v
    port map (
            O => \N__63271\,
            I => \N__63210\
        );

    \I__13968\ : LocalMux
    port map (
            O => \N__63268\,
            I => \N__63210\
        );

    \I__13967\ : LocalMux
    port map (
            O => \N__63255\,
            I => \N__63207\
        );

    \I__13966\ : Span4Mux_v
    port map (
            O => \N__63252\,
            I => \N__63200\
        );

    \I__13965\ : Span4Mux_h
    port map (
            O => \N__63247\,
            I => \N__63200\
        );

    \I__13964\ : Span4Mux_v
    port map (
            O => \N__63238\,
            I => \N__63200\
        );

    \I__13963\ : InMux
    port map (
            O => \N__63237\,
            I => \N__63187\
        );

    \I__13962\ : InMux
    port map (
            O => \N__63234\,
            I => \N__63187\
        );

    \I__13961\ : InMux
    port map (
            O => \N__63233\,
            I => \N__63187\
        );

    \I__13960\ : InMux
    port map (
            O => \N__63230\,
            I => \N__63187\
        );

    \I__13959\ : InMux
    port map (
            O => \N__63229\,
            I => \N__63187\
        );

    \I__13958\ : InMux
    port map (
            O => \N__63226\,
            I => \N__63187\
        );

    \I__13957\ : LocalMux
    port map (
            O => \N__63221\,
            I => \N__63184\
        );

    \I__13956\ : InMux
    port map (
            O => \N__63218\,
            I => \N__63181\
        );

    \I__13955\ : Span4Mux_v
    port map (
            O => \N__63215\,
            I => \N__63177\
        );

    \I__13954\ : Span4Mux_v
    port map (
            O => \N__63210\,
            I => \N__63174\
        );

    \I__13953\ : Span4Mux_v
    port map (
            O => \N__63207\,
            I => \N__63167\
        );

    \I__13952\ : Span4Mux_h
    port map (
            O => \N__63200\,
            I => \N__63167\
        );

    \I__13951\ : LocalMux
    port map (
            O => \N__63187\,
            I => \N__63167\
        );

    \I__13950\ : Span4Mux_h
    port map (
            O => \N__63184\,
            I => \N__63162\
        );

    \I__13949\ : LocalMux
    port map (
            O => \N__63181\,
            I => \N__63162\
        );

    \I__13948\ : InMux
    port map (
            O => \N__63180\,
            I => \N__63159\
        );

    \I__13947\ : Odrv4
    port map (
            O => \N__63177\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\
        );

    \I__13946\ : Odrv4
    port map (
            O => \N__63174\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\
        );

    \I__13945\ : Odrv4
    port map (
            O => \N__63167\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\
        );

    \I__13944\ : Odrv4
    port map (
            O => \N__63162\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\
        );

    \I__13943\ : LocalMux
    port map (
            O => \N__63159\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\
        );

    \I__13942\ : InMux
    port map (
            O => \N__63148\,
            I => \N__63145\
        );

    \I__13941\ : LocalMux
    port map (
            O => \N__63145\,
            I => \N__63142\
        );

    \I__13940\ : Odrv4
    port map (
            O => \N__63142\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n317\
        );

    \I__13939\ : InMux
    port map (
            O => \N__63139\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18268\
        );

    \I__13938\ : CascadeMux
    port map (
            O => \N__63136\,
            I => \N__63128\
        );

    \I__13937\ : CascadeMux
    port map (
            O => \N__63135\,
            I => \N__63124\
        );

    \I__13936\ : CascadeMux
    port map (
            O => \N__63134\,
            I => \N__63121\
        );

    \I__13935\ : CascadeMux
    port map (
            O => \N__63133\,
            I => \N__63118\
        );

    \I__13934\ : CascadeMux
    port map (
            O => \N__63132\,
            I => \N__63115\
        );

    \I__13933\ : CascadeMux
    port map (
            O => \N__63131\,
            I => \N__63106\
        );

    \I__13932\ : InMux
    port map (
            O => \N__63128\,
            I => \N__63103\
        );

    \I__13931\ : CascadeMux
    port map (
            O => \N__63127\,
            I => \N__63100\
        );

    \I__13930\ : InMux
    port map (
            O => \N__63124\,
            I => \N__63084\
        );

    \I__13929\ : InMux
    port map (
            O => \N__63121\,
            I => \N__63084\
        );

    \I__13928\ : InMux
    port map (
            O => \N__63118\,
            I => \N__63084\
        );

    \I__13927\ : InMux
    port map (
            O => \N__63115\,
            I => \N__63084\
        );

    \I__13926\ : CascadeMux
    port map (
            O => \N__63114\,
            I => \N__63081\
        );

    \I__13925\ : CascadeMux
    port map (
            O => \N__63113\,
            I => \N__63078\
        );

    \I__13924\ : CascadeMux
    port map (
            O => \N__63112\,
            I => \N__63075\
        );

    \I__13923\ : CascadeMux
    port map (
            O => \N__63111\,
            I => \N__63072\
        );

    \I__13922\ : InMux
    port map (
            O => \N__63110\,
            I => \N__63069\
        );

    \I__13921\ : CascadeMux
    port map (
            O => \N__63109\,
            I => \N__63066\
        );

    \I__13920\ : InMux
    port map (
            O => \N__63106\,
            I => \N__63062\
        );

    \I__13919\ : LocalMux
    port map (
            O => \N__63103\,
            I => \N__63059\
        );

    \I__13918\ : InMux
    port map (
            O => \N__63100\,
            I => \N__63056\
        );

    \I__13917\ : CascadeMux
    port map (
            O => \N__63099\,
            I => \N__63053\
        );

    \I__13916\ : CascadeMux
    port map (
            O => \N__63098\,
            I => \N__63049\
        );

    \I__13915\ : CascadeMux
    port map (
            O => \N__63097\,
            I => \N__63045\
        );

    \I__13914\ : CascadeMux
    port map (
            O => \N__63096\,
            I => \N__63041\
        );

    \I__13913\ : CascadeMux
    port map (
            O => \N__63095\,
            I => \N__63038\
        );

    \I__13912\ : InMux
    port map (
            O => \N__63094\,
            I => \N__63035\
        );

    \I__13911\ : InMux
    port map (
            O => \N__63093\,
            I => \N__63032\
        );

    \I__13910\ : LocalMux
    port map (
            O => \N__63084\,
            I => \N__63028\
        );

    \I__13909\ : InMux
    port map (
            O => \N__63081\,
            I => \N__63019\
        );

    \I__13908\ : InMux
    port map (
            O => \N__63078\,
            I => \N__63019\
        );

    \I__13907\ : InMux
    port map (
            O => \N__63075\,
            I => \N__63019\
        );

    \I__13906\ : InMux
    port map (
            O => \N__63072\,
            I => \N__63019\
        );

    \I__13905\ : LocalMux
    port map (
            O => \N__63069\,
            I => \N__63016\
        );

    \I__13904\ : InMux
    port map (
            O => \N__63066\,
            I => \N__63013\
        );

    \I__13903\ : CascadeMux
    port map (
            O => \N__63065\,
            I => \N__63010\
        );

    \I__13902\ : LocalMux
    port map (
            O => \N__63062\,
            I => \N__63003\
        );

    \I__13901\ : Span4Mux_v
    port map (
            O => \N__63059\,
            I => \N__63003\
        );

    \I__13900\ : LocalMux
    port map (
            O => \N__63056\,
            I => \N__63003\
        );

    \I__13899\ : InMux
    port map (
            O => \N__63053\,
            I => \N__63000\
        );

    \I__13898\ : InMux
    port map (
            O => \N__63052\,
            I => \N__62986\
        );

    \I__13897\ : InMux
    port map (
            O => \N__63049\,
            I => \N__62986\
        );

    \I__13896\ : InMux
    port map (
            O => \N__63048\,
            I => \N__62986\
        );

    \I__13895\ : InMux
    port map (
            O => \N__63045\,
            I => \N__62986\
        );

    \I__13894\ : InMux
    port map (
            O => \N__63044\,
            I => \N__62986\
        );

    \I__13893\ : InMux
    port map (
            O => \N__63041\,
            I => \N__62986\
        );

    \I__13892\ : InMux
    port map (
            O => \N__63038\,
            I => \N__62983\
        );

    \I__13891\ : LocalMux
    port map (
            O => \N__63035\,
            I => \N__62978\
        );

    \I__13890\ : LocalMux
    port map (
            O => \N__63032\,
            I => \N__62978\
        );

    \I__13889\ : CascadeMux
    port map (
            O => \N__63031\,
            I => \N__62975\
        );

    \I__13888\ : Span4Mux_v
    port map (
            O => \N__63028\,
            I => \N__62971\
        );

    \I__13887\ : LocalMux
    port map (
            O => \N__63019\,
            I => \N__62968\
        );

    \I__13886\ : Span4Mux_h
    port map (
            O => \N__63016\,
            I => \N__62963\
        );

    \I__13885\ : LocalMux
    port map (
            O => \N__63013\,
            I => \N__62963\
        );

    \I__13884\ : InMux
    port map (
            O => \N__63010\,
            I => \N__62960\
        );

    \I__13883\ : Span4Mux_h
    port map (
            O => \N__63003\,
            I => \N__62954\
        );

    \I__13882\ : LocalMux
    port map (
            O => \N__63000\,
            I => \N__62954\
        );

    \I__13881\ : InMux
    port map (
            O => \N__62999\,
            I => \N__62951\
        );

    \I__13880\ : LocalMux
    port map (
            O => \N__62986\,
            I => \N__62948\
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__62983\,
            I => \N__62945\
        );

    \I__13878\ : Span4Mux_v
    port map (
            O => \N__62978\,
            I => \N__62942\
        );

    \I__13877\ : InMux
    port map (
            O => \N__62975\,
            I => \N__62939\
        );

    \I__13876\ : CascadeMux
    port map (
            O => \N__62974\,
            I => \N__62935\
        );

    \I__13875\ : Span4Mux_h
    port map (
            O => \N__62971\,
            I => \N__62930\
        );

    \I__13874\ : Span4Mux_v
    port map (
            O => \N__62968\,
            I => \N__62930\
        );

    \I__13873\ : Span4Mux_v
    port map (
            O => \N__62963\,
            I => \N__62925\
        );

    \I__13872\ : LocalMux
    port map (
            O => \N__62960\,
            I => \N__62925\
        );

    \I__13871\ : CascadeMux
    port map (
            O => \N__62959\,
            I => \N__62922\
        );

    \I__13870\ : Span4Mux_v
    port map (
            O => \N__62954\,
            I => \N__62919\
        );

    \I__13869\ : LocalMux
    port map (
            O => \N__62951\,
            I => \N__62916\
        );

    \I__13868\ : Span4Mux_v
    port map (
            O => \N__62948\,
            I => \N__62913\
        );

    \I__13867\ : Span4Mux_v
    port map (
            O => \N__62945\,
            I => \N__62906\
        );

    \I__13866\ : Span4Mux_h
    port map (
            O => \N__62942\,
            I => \N__62906\
        );

    \I__13865\ : LocalMux
    port map (
            O => \N__62939\,
            I => \N__62906\
        );

    \I__13864\ : InMux
    port map (
            O => \N__62938\,
            I => \N__62903\
        );

    \I__13863\ : InMux
    port map (
            O => \N__62935\,
            I => \N__62900\
        );

    \I__13862\ : Span4Mux_h
    port map (
            O => \N__62930\,
            I => \N__62895\
        );

    \I__13861\ : Span4Mux_v
    port map (
            O => \N__62925\,
            I => \N__62895\
        );

    \I__13860\ : InMux
    port map (
            O => \N__62922\,
            I => \N__62892\
        );

    \I__13859\ : Span4Mux_h
    port map (
            O => \N__62919\,
            I => \N__62887\
        );

    \I__13858\ : Span4Mux_v
    port map (
            O => \N__62916\,
            I => \N__62887\
        );

    \I__13857\ : Span4Mux_h
    port map (
            O => \N__62913\,
            I => \N__62882\
        );

    \I__13856\ : Span4Mux_h
    port map (
            O => \N__62906\,
            I => \N__62882\
        );

    \I__13855\ : LocalMux
    port map (
            O => \N__62903\,
            I => \N__62879\
        );

    \I__13854\ : LocalMux
    port map (
            O => \N__62900\,
            I => \N__62872\
        );

    \I__13853\ : Span4Mux_h
    port map (
            O => \N__62895\,
            I => \N__62872\
        );

    \I__13852\ : LocalMux
    port map (
            O => \N__62892\,
            I => \N__62872\
        );

    \I__13851\ : Span4Mux_v
    port map (
            O => \N__62887\,
            I => \N__62869\
        );

    \I__13850\ : Span4Mux_v
    port map (
            O => \N__62882\,
            I => \N__62866\
        );

    \I__13849\ : Span4Mux_h
    port map (
            O => \N__62879\,
            I => \N__62861\
        );

    \I__13848\ : Span4Mux_v
    port map (
            O => \N__62872\,
            I => \N__62861\
        );

    \I__13847\ : Odrv4
    port map (
            O => \N__62869\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n120\
        );

    \I__13846\ : Odrv4
    port map (
            O => \N__62866\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n120\
        );

    \I__13845\ : Odrv4
    port map (
            O => \N__62861\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n120\
        );

    \I__13844\ : CascadeMux
    port map (
            O => \N__62854\,
            I => \N__62851\
        );

    \I__13843\ : InMux
    port map (
            O => \N__62851\,
            I => \N__62848\
        );

    \I__13842\ : LocalMux
    port map (
            O => \N__62848\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n320\
        );

    \I__13841\ : InMux
    port map (
            O => \N__62845\,
            I => \N__62842\
        );

    \I__13840\ : LocalMux
    port map (
            O => \N__62842\,
            I => \N__62839\
        );

    \I__13839\ : Odrv4
    port map (
            O => \N__62839\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n366\
        );

    \I__13838\ : InMux
    port map (
            O => \N__62836\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18269\
        );

    \I__13837\ : InMux
    port map (
            O => \N__62833\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18255\
        );

    \I__13836\ : InMux
    port map (
            O => \N__62830\,
            I => \N__62827\
        );

    \I__13835\ : LocalMux
    port map (
            O => \N__62827\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n461\
        );

    \I__13834\ : InMux
    port map (
            O => \N__62824\,
            I => \bfn_23_26_0_\
        );

    \I__13833\ : InMux
    port map (
            O => \N__62821\,
            I => \N__62818\
        );

    \I__13832\ : LocalMux
    port map (
            O => \N__62818\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n510\
        );

    \I__13831\ : InMux
    port map (
            O => \N__62815\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18257\
        );

    \I__13830\ : InMux
    port map (
            O => \N__62812\,
            I => \N__62809\
        );

    \I__13829\ : LocalMux
    port map (
            O => \N__62809\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n559\
        );

    \I__13828\ : InMux
    port map (
            O => \N__62806\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18258\
        );

    \I__13827\ : InMux
    port map (
            O => \N__62803\,
            I => \N__62800\
        );

    \I__13826\ : LocalMux
    port map (
            O => \N__62800\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n608\
        );

    \I__13825\ : InMux
    port map (
            O => \N__62797\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18259\
        );

    \I__13824\ : CascadeMux
    port map (
            O => \N__62794\,
            I => \N__62791\
        );

    \I__13823\ : InMux
    port map (
            O => \N__62791\,
            I => \N__62788\
        );

    \I__13822\ : LocalMux
    port map (
            O => \N__62788\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n657\
        );

    \I__13821\ : InMux
    port map (
            O => \N__62785\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18260\
        );

    \I__13820\ : CascadeMux
    port map (
            O => \N__62782\,
            I => \N__62779\
        );

    \I__13819\ : InMux
    port map (
            O => \N__62779\,
            I => \N__62776\
        );

    \I__13818\ : LocalMux
    port map (
            O => \N__62776\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n706\
        );

    \I__13817\ : InMux
    port map (
            O => \N__62773\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18261\
        );

    \I__13816\ : InMux
    port map (
            O => \N__62770\,
            I => \N__62767\
        );

    \I__13815\ : LocalMux
    port map (
            O => \N__62767\,
            I => \N__62764\
        );

    \I__13814\ : Span4Mux_v
    port map (
            O => \N__62764\,
            I => \N__62761\
        );

    \I__13813\ : Span4Mux_h
    port map (
            O => \N__62761\,
            I => \N__62758\
        );

    \I__13812\ : Odrv4
    port map (
            O => \N__62758\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n762\
        );

    \I__13811\ : InMux
    port map (
            O => \N__62755\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18262\
        );

    \I__13810\ : InMux
    port map (
            O => \N__62752\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763\
        );

    \I__13809\ : CascadeMux
    port map (
            O => \N__62749\,
            I => \N__62746\
        );

    \I__13808\ : InMux
    port map (
            O => \N__62746\,
            I => \N__62743\
        );

    \I__13807\ : LocalMux
    port map (
            O => \N__62743\,
            I => \N__62740\
        );

    \I__13806\ : Span4Mux_h
    port map (
            O => \N__62740\,
            I => \N__62737\
        );

    \I__13805\ : Span4Mux_v
    port map (
            O => \N__62737\,
            I => \N__62734\
        );

    \I__13804\ : Odrv4
    port map (
            O => \N__62734\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_CO\
        );

    \I__13803\ : InMux
    port map (
            O => \N__62731\,
            I => \N__62728\
        );

    \I__13802\ : LocalMux
    port map (
            O => \N__62728\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19755\
        );

    \I__13801\ : InMux
    port map (
            O => \N__62725\,
            I => \N__62722\
        );

    \I__13800\ : LocalMux
    port map (
            O => \N__62722\,
            I => \N__62718\
        );

    \I__13799\ : InMux
    port map (
            O => \N__62721\,
            I => \N__62715\
        );

    \I__13798\ : Span4Mux_h
    port map (
            O => \N__62718\,
            I => \N__62711\
        );

    \I__13797\ : LocalMux
    port map (
            O => \N__62715\,
            I => \N__62708\
        );

    \I__13796\ : InMux
    port map (
            O => \N__62714\,
            I => \N__62705\
        );

    \I__13795\ : Odrv4
    port map (
            O => \N__62711\,
            I => \Add_add_temp_11_adj_2409\
        );

    \I__13794\ : Odrv4
    port map (
            O => \N__62708\,
            I => \Add_add_temp_11_adj_2409\
        );

    \I__13793\ : LocalMux
    port map (
            O => \N__62705\,
            I => \Add_add_temp_11_adj_2409\
        );

    \I__13792\ : CascadeMux
    port map (
            O => \N__62698\,
            I => \N__62694\
        );

    \I__13791\ : InMux
    port map (
            O => \N__62697\,
            I => \N__62691\
        );

    \I__13790\ : InMux
    port map (
            O => \N__62694\,
            I => \N__62688\
        );

    \I__13789\ : LocalMux
    port map (
            O => \N__62691\,
            I => \N__62684\
        );

    \I__13788\ : LocalMux
    port map (
            O => \N__62688\,
            I => \N__62681\
        );

    \I__13787\ : InMux
    port map (
            O => \N__62687\,
            I => \N__62678\
        );

    \I__13786\ : Odrv12
    port map (
            O => \N__62684\,
            I => \Add_add_temp_9_adj_2411\
        );

    \I__13785\ : Odrv4
    port map (
            O => \N__62681\,
            I => \Add_add_temp_9_adj_2411\
        );

    \I__13784\ : LocalMux
    port map (
            O => \N__62678\,
            I => \Add_add_temp_9_adj_2411\
        );

    \I__13783\ : InMux
    port map (
            O => \N__62671\,
            I => \N__62668\
        );

    \I__13782\ : LocalMux
    port map (
            O => \N__62668\,
            I => \N__62664\
        );

    \I__13781\ : InMux
    port map (
            O => \N__62667\,
            I => \N__62661\
        );

    \I__13780\ : Span4Mux_v
    port map (
            O => \N__62664\,
            I => \N__62655\
        );

    \I__13779\ : LocalMux
    port map (
            O => \N__62661\,
            I => \N__62655\
        );

    \I__13778\ : InMux
    port map (
            O => \N__62660\,
            I => \N__62652\
        );

    \I__13777\ : Odrv4
    port map (
            O => \N__62655\,
            I => \Add_add_temp_10_adj_2410\
        );

    \I__13776\ : LocalMux
    port map (
            O => \N__62652\,
            I => \Add_add_temp_10_adj_2410\
        );

    \I__13775\ : InMux
    port map (
            O => \N__62647\,
            I => \N__62644\
        );

    \I__13774\ : LocalMux
    port map (
            O => \N__62644\,
            I => \N__62641\
        );

    \I__13773\ : Span4Mux_h
    port map (
            O => \N__62641\,
            I => \N__62638\
        );

    \I__13772\ : Odrv4
    port map (
            O => \N__62638\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20718\
        );

    \I__13771\ : InMux
    port map (
            O => \N__62635\,
            I => \N__62632\
        );

    \I__13770\ : LocalMux
    port map (
            O => \N__62632\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n72\
        );

    \I__13769\ : InMux
    port map (
            O => \N__62629\,
            I => \N__62626\
        );

    \I__13768\ : LocalMux
    port map (
            O => \N__62626\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n118\
        );

    \I__13767\ : InMux
    port map (
            O => \N__62623\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18249\
        );

    \I__13766\ : InMux
    port map (
            O => \N__62620\,
            I => \N__62617\
        );

    \I__13765\ : LocalMux
    port map (
            O => \N__62617\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n167\
        );

    \I__13764\ : InMux
    port map (
            O => \N__62614\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18250\
        );

    \I__13763\ : InMux
    port map (
            O => \N__62611\,
            I => \N__62608\
        );

    \I__13762\ : LocalMux
    port map (
            O => \N__62608\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n216\
        );

    \I__13761\ : InMux
    port map (
            O => \N__62605\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18251\
        );

    \I__13760\ : InMux
    port map (
            O => \N__62602\,
            I => \N__62599\
        );

    \I__13759\ : LocalMux
    port map (
            O => \N__62599\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n265\
        );

    \I__13758\ : InMux
    port map (
            O => \N__62596\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18252\
        );

    \I__13757\ : InMux
    port map (
            O => \N__62593\,
            I => \N__62590\
        );

    \I__13756\ : LocalMux
    port map (
            O => \N__62590\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n314\
        );

    \I__13755\ : InMux
    port map (
            O => \N__62587\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18253\
        );

    \I__13754\ : InMux
    port map (
            O => \N__62584\,
            I => \N__62581\
        );

    \I__13753\ : LocalMux
    port map (
            O => \N__62581\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n363\
        );

    \I__13752\ : InMux
    port map (
            O => \N__62578\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18254\
        );

    \I__13751\ : InMux
    port map (
            O => \N__62575\,
            I => \N__62572\
        );

    \I__13750\ : LocalMux
    port map (
            O => \N__62572\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n412\
        );

    \I__13749\ : InMux
    port map (
            O => \N__62569\,
            I => \N__62566\
        );

    \I__13748\ : LocalMux
    port map (
            O => \N__62566\,
            I => \N__62561\
        );

    \I__13747\ : InMux
    port map (
            O => \N__62565\,
            I => \N__62556\
        );

    \I__13746\ : InMux
    port map (
            O => \N__62564\,
            I => \N__62556\
        );

    \I__13745\ : Odrv12
    port map (
            O => \N__62561\,
            I => \Add_add_temp_5\
        );

    \I__13744\ : LocalMux
    port map (
            O => \N__62556\,
            I => \Add_add_temp_5\
        );

    \I__13743\ : InMux
    port map (
            O => \N__62551\,
            I => \N__62548\
        );

    \I__13742\ : LocalMux
    port map (
            O => \N__62548\,
            I => \N__62544\
        );

    \I__13741\ : InMux
    port map (
            O => \N__62547\,
            I => \N__62541\
        );

    \I__13740\ : Odrv4
    port map (
            O => \N__62544\,
            I => \Add_add_temp_4\
        );

    \I__13739\ : LocalMux
    port map (
            O => \N__62541\,
            I => \Add_add_temp_4\
        );

    \I__13738\ : InMux
    port map (
            O => \N__62536\,
            I => \N__62531\
        );

    \I__13737\ : InMux
    port map (
            O => \N__62535\,
            I => \N__62528\
        );

    \I__13736\ : InMux
    port map (
            O => \N__62534\,
            I => \N__62525\
        );

    \I__13735\ : LocalMux
    port map (
            O => \N__62531\,
            I => \Add_add_temp_8\
        );

    \I__13734\ : LocalMux
    port map (
            O => \N__62528\,
            I => \Add_add_temp_8\
        );

    \I__13733\ : LocalMux
    port map (
            O => \N__62525\,
            I => \Add_add_temp_8\
        );

    \I__13732\ : InMux
    port map (
            O => \N__62518\,
            I => \N__62513\
        );

    \I__13731\ : CascadeMux
    port map (
            O => \N__62517\,
            I => \N__62510\
        );

    \I__13730\ : InMux
    port map (
            O => \N__62516\,
            I => \N__62507\
        );

    \I__13729\ : LocalMux
    port map (
            O => \N__62513\,
            I => \N__62504\
        );

    \I__13728\ : InMux
    port map (
            O => \N__62510\,
            I => \N__62501\
        );

    \I__13727\ : LocalMux
    port map (
            O => \N__62507\,
            I => \Add_add_temp_7\
        );

    \I__13726\ : Odrv4
    port map (
            O => \N__62504\,
            I => \Add_add_temp_7\
        );

    \I__13725\ : LocalMux
    port map (
            O => \N__62501\,
            I => \Add_add_temp_7\
        );

    \I__13724\ : CascadeMux
    port map (
            O => \N__62494\,
            I => \N__62491\
        );

    \I__13723\ : InMux
    port map (
            O => \N__62491\,
            I => \N__62487\
        );

    \I__13722\ : InMux
    port map (
            O => \N__62490\,
            I => \N__62484\
        );

    \I__13721\ : LocalMux
    port map (
            O => \N__62487\,
            I => \N__62480\
        );

    \I__13720\ : LocalMux
    port map (
            O => \N__62484\,
            I => \N__62477\
        );

    \I__13719\ : InMux
    port map (
            O => \N__62483\,
            I => \N__62474\
        );

    \I__13718\ : Odrv4
    port map (
            O => \N__62480\,
            I => \Add_add_temp_6\
        );

    \I__13717\ : Odrv12
    port map (
            O => \N__62477\,
            I => \Add_add_temp_6\
        );

    \I__13716\ : LocalMux
    port map (
            O => \N__62474\,
            I => \Add_add_temp_6\
        );

    \I__13715\ : InMux
    port map (
            O => \N__62467\,
            I => \N__62464\
        );

    \I__13714\ : LocalMux
    port map (
            O => \N__62464\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20712\
        );

    \I__13713\ : InMux
    port map (
            O => \N__62461\,
            I => \N__62456\
        );

    \I__13712\ : InMux
    port map (
            O => \N__62460\,
            I => \N__62453\
        );

    \I__13711\ : InMux
    port map (
            O => \N__62459\,
            I => \N__62450\
        );

    \I__13710\ : LocalMux
    port map (
            O => \N__62456\,
            I => \Add_add_temp_9\
        );

    \I__13709\ : LocalMux
    port map (
            O => \N__62453\,
            I => \Add_add_temp_9\
        );

    \I__13708\ : LocalMux
    port map (
            O => \N__62450\,
            I => \Add_add_temp_9\
        );

    \I__13707\ : InMux
    port map (
            O => \N__62443\,
            I => \N__62440\
        );

    \I__13706\ : LocalMux
    port map (
            O => \N__62440\,
            I => \N__62437\
        );

    \I__13705\ : Span4Mux_v
    port map (
            O => \N__62437\,
            I => \N__62432\
        );

    \I__13704\ : InMux
    port map (
            O => \N__62436\,
            I => \N__62429\
        );

    \I__13703\ : InMux
    port map (
            O => \N__62435\,
            I => \N__62426\
        );

    \I__13702\ : Odrv4
    port map (
            O => \N__62432\,
            I => \Add_add_temp_11\
        );

    \I__13701\ : LocalMux
    port map (
            O => \N__62429\,
            I => \Add_add_temp_11\
        );

    \I__13700\ : LocalMux
    port map (
            O => \N__62426\,
            I => \Add_add_temp_11\
        );

    \I__13699\ : CascadeMux
    port map (
            O => \N__62419\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19777_cascade_\
        );

    \I__13698\ : InMux
    port map (
            O => \N__62416\,
            I => \N__62412\
        );

    \I__13697\ : InMux
    port map (
            O => \N__62415\,
            I => \N__62408\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__62412\,
            I => \N__62405\
        );

    \I__13695\ : InMux
    port map (
            O => \N__62411\,
            I => \N__62402\
        );

    \I__13694\ : LocalMux
    port map (
            O => \N__62408\,
            I => \Add_add_temp_10\
        );

    \I__13693\ : Odrv4
    port map (
            O => \N__62405\,
            I => \Add_add_temp_10\
        );

    \I__13692\ : LocalMux
    port map (
            O => \N__62402\,
            I => \Add_add_temp_10\
        );

    \I__13691\ : InMux
    port map (
            O => \N__62395\,
            I => \N__62392\
        );

    \I__13690\ : LocalMux
    port map (
            O => \N__62392\,
            I => \N__62389\
        );

    \I__13689\ : Span4Mux_h
    port map (
            O => \N__62389\,
            I => \N__62384\
        );

    \I__13688\ : InMux
    port map (
            O => \N__62388\,
            I => \N__62381\
        );

    \I__13687\ : InMux
    port map (
            O => \N__62387\,
            I => \N__62378\
        );

    \I__13686\ : Odrv4
    port map (
            O => \N__62384\,
            I => \Add_add_temp_14\
        );

    \I__13685\ : LocalMux
    port map (
            O => \N__62381\,
            I => \Add_add_temp_14\
        );

    \I__13684\ : LocalMux
    port map (
            O => \N__62378\,
            I => \Add_add_temp_14\
        );

    \I__13683\ : InMux
    port map (
            O => \N__62371\,
            I => \N__62368\
        );

    \I__13682\ : LocalMux
    port map (
            O => \N__62368\,
            I => \N__62363\
        );

    \I__13681\ : InMux
    port map (
            O => \N__62367\,
            I => \N__62360\
        );

    \I__13680\ : InMux
    port map (
            O => \N__62366\,
            I => \N__62357\
        );

    \I__13679\ : Odrv4
    port map (
            O => \N__62363\,
            I => \Add_add_temp_13\
        );

    \I__13678\ : LocalMux
    port map (
            O => \N__62360\,
            I => \Add_add_temp_13\
        );

    \I__13677\ : LocalMux
    port map (
            O => \N__62357\,
            I => \Add_add_temp_13\
        );

    \I__13676\ : CascadeMux
    port map (
            O => \N__62350\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20700_cascade_\
        );

    \I__13675\ : InMux
    port map (
            O => \N__62347\,
            I => \N__62344\
        );

    \I__13674\ : LocalMux
    port map (
            O => \N__62344\,
            I => \N__62341\
        );

    \I__13673\ : Span4Mux_v
    port map (
            O => \N__62341\,
            I => \N__62336\
        );

    \I__13672\ : InMux
    port map (
            O => \N__62340\,
            I => \N__62333\
        );

    \I__13671\ : InMux
    port map (
            O => \N__62339\,
            I => \N__62330\
        );

    \I__13670\ : Odrv4
    port map (
            O => \N__62336\,
            I => \Add_add_temp_12\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__62333\,
            I => \Add_add_temp_12\
        );

    \I__13668\ : LocalMux
    port map (
            O => \N__62330\,
            I => \Add_add_temp_12\
        );

    \I__13667\ : InMux
    port map (
            O => \N__62323\,
            I => \N__62320\
        );

    \I__13666\ : LocalMux
    port map (
            O => \N__62320\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15205\
        );

    \I__13665\ : InMux
    port map (
            O => \N__62317\,
            I => \N__62314\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__62314\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20670\
        );

    \I__13663\ : InMux
    port map (
            O => \N__62311\,
            I => \N__62308\
        );

    \I__13662\ : LocalMux
    port map (
            O => \N__62308\,
            I => \N__62304\
        );

    \I__13661\ : InMux
    port map (
            O => \N__62307\,
            I => \N__62301\
        );

    \I__13660\ : Span4Mux_h
    port map (
            O => \N__62304\,
            I => \N__62297\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__62301\,
            I => \N__62294\
        );

    \I__13658\ : InMux
    port map (
            O => \N__62300\,
            I => \N__62291\
        );

    \I__13657\ : Odrv4
    port map (
            O => \N__62297\,
            I => \Add_add_temp_20\
        );

    \I__13656\ : Odrv12
    port map (
            O => \N__62294\,
            I => \Add_add_temp_20\
        );

    \I__13655\ : LocalMux
    port map (
            O => \N__62291\,
            I => \Add_add_temp_20\
        );

    \I__13654\ : CascadeMux
    port map (
            O => \N__62284\,
            I => \N__62280\
        );

    \I__13653\ : InMux
    port map (
            O => \N__62283\,
            I => \N__62276\
        );

    \I__13652\ : InMux
    port map (
            O => \N__62280\,
            I => \N__62273\
        );

    \I__13651\ : CascadeMux
    port map (
            O => \N__62279\,
            I => \N__62270\
        );

    \I__13650\ : LocalMux
    port map (
            O => \N__62276\,
            I => \N__62267\
        );

    \I__13649\ : LocalMux
    port map (
            O => \N__62273\,
            I => \N__62264\
        );

    \I__13648\ : InMux
    port map (
            O => \N__62270\,
            I => \N__62261\
        );

    \I__13647\ : Odrv4
    port map (
            O => \N__62267\,
            I => \Add_add_temp_18\
        );

    \I__13646\ : Odrv4
    port map (
            O => \N__62264\,
            I => \Add_add_temp_18\
        );

    \I__13645\ : LocalMux
    port map (
            O => \N__62261\,
            I => \Add_add_temp_18\
        );

    \I__13644\ : InMux
    port map (
            O => \N__62254\,
            I => \N__62251\
        );

    \I__13643\ : LocalMux
    port map (
            O => \N__62251\,
            I => \N__62247\
        );

    \I__13642\ : InMux
    port map (
            O => \N__62250\,
            I => \N__62244\
        );

    \I__13641\ : Span4Mux_h
    port map (
            O => \N__62247\,
            I => \N__62238\
        );

    \I__13640\ : LocalMux
    port map (
            O => \N__62244\,
            I => \N__62238\
        );

    \I__13639\ : InMux
    port map (
            O => \N__62243\,
            I => \N__62235\
        );

    \I__13638\ : Odrv4
    port map (
            O => \N__62238\,
            I => \Add_add_temp_19\
        );

    \I__13637\ : LocalMux
    port map (
            O => \N__62235\,
            I => \Add_add_temp_19\
        );

    \I__13636\ : InMux
    port map (
            O => \N__62230\,
            I => \N__62227\
        );

    \I__13635\ : LocalMux
    port map (
            O => \N__62227\,
            I => \N__62223\
        );

    \I__13634\ : InMux
    port map (
            O => \N__62226\,
            I => \N__62220\
        );

    \I__13633\ : Span4Mux_v
    port map (
            O => \N__62223\,
            I => \N__62215\
        );

    \I__13632\ : LocalMux
    port map (
            O => \N__62220\,
            I => \N__62215\
        );

    \I__13631\ : Span4Mux_h
    port map (
            O => \N__62215\,
            I => \N__62211\
        );

    \I__13630\ : InMux
    port map (
            O => \N__62214\,
            I => \N__62208\
        );

    \I__13629\ : Odrv4
    port map (
            O => \N__62211\,
            I => \Add_add_temp_21\
        );

    \I__13628\ : LocalMux
    port map (
            O => \N__62208\,
            I => \Add_add_temp_21\
        );

    \I__13627\ : InMux
    port map (
            O => \N__62203\,
            I => \N__62199\
        );

    \I__13626\ : InMux
    port map (
            O => \N__62202\,
            I => \N__62196\
        );

    \I__13625\ : LocalMux
    port map (
            O => \N__62199\,
            I => \N__62191\
        );

    \I__13624\ : LocalMux
    port map (
            O => \N__62196\,
            I => \N__62191\
        );

    \I__13623\ : Span4Mux_h
    port map (
            O => \N__62191\,
            I => \N__62187\
        );

    \I__13622\ : InMux
    port map (
            O => \N__62190\,
            I => \N__62184\
        );

    \I__13621\ : Odrv4
    port map (
            O => \N__62187\,
            I => \Add_add_temp_23\
        );

    \I__13620\ : LocalMux
    port map (
            O => \N__62184\,
            I => \Add_add_temp_23\
        );

    \I__13619\ : CascadeMux
    port map (
            O => \N__62179\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19746_cascade_\
        );

    \I__13618\ : InMux
    port map (
            O => \N__62176\,
            I => \N__62172\
        );

    \I__13617\ : InMux
    port map (
            O => \N__62175\,
            I => \N__62169\
        );

    \I__13616\ : LocalMux
    port map (
            O => \N__62172\,
            I => \N__62166\
        );

    \I__13615\ : LocalMux
    port map (
            O => \N__62169\,
            I => \N__62160\
        );

    \I__13614\ : Sp12to4
    port map (
            O => \N__62166\,
            I => \N__62160\
        );

    \I__13613\ : InMux
    port map (
            O => \N__62165\,
            I => \N__62157\
        );

    \I__13612\ : Odrv12
    port map (
            O => \N__62160\,
            I => \Add_add_temp_22\
        );

    \I__13611\ : LocalMux
    port map (
            O => \N__62157\,
            I => \Add_add_temp_22\
        );

    \I__13610\ : InMux
    port map (
            O => \N__62152\,
            I => \N__62149\
        );

    \I__13609\ : LocalMux
    port map (
            O => \N__62149\,
            I => \N__62146\
        );

    \I__13608\ : Odrv4
    port map (
            O => \N__62146\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20656\
        );

    \I__13607\ : InMux
    port map (
            O => \N__62143\,
            I => \N__62139\
        );

    \I__13606\ : InMux
    port map (
            O => \N__62142\,
            I => \N__62136\
        );

    \I__13605\ : LocalMux
    port map (
            O => \N__62139\,
            I => \N__62131\
        );

    \I__13604\ : LocalMux
    port map (
            O => \N__62136\,
            I => \N__62131\
        );

    \I__13603\ : Span4Mux_v
    port map (
            O => \N__62131\,
            I => \N__62127\
        );

    \I__13602\ : InMux
    port map (
            O => \N__62130\,
            I => \N__62124\
        );

    \I__13601\ : Odrv4
    port map (
            O => \N__62127\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31\
        );

    \I__13600\ : LocalMux
    port map (
            O => \N__62124\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31\
        );

    \I__13599\ : ClkMux
    port map (
            O => \N__62119\,
            I => \N__62071\
        );

    \I__13598\ : ClkMux
    port map (
            O => \N__62118\,
            I => \N__62071\
        );

    \I__13597\ : ClkMux
    port map (
            O => \N__62117\,
            I => \N__62071\
        );

    \I__13596\ : ClkMux
    port map (
            O => \N__62116\,
            I => \N__62071\
        );

    \I__13595\ : ClkMux
    port map (
            O => \N__62115\,
            I => \N__62071\
        );

    \I__13594\ : ClkMux
    port map (
            O => \N__62114\,
            I => \N__62071\
        );

    \I__13593\ : ClkMux
    port map (
            O => \N__62113\,
            I => \N__62071\
        );

    \I__13592\ : ClkMux
    port map (
            O => \N__62112\,
            I => \N__62071\
        );

    \I__13591\ : ClkMux
    port map (
            O => \N__62111\,
            I => \N__62071\
        );

    \I__13590\ : ClkMux
    port map (
            O => \N__62110\,
            I => \N__62071\
        );

    \I__13589\ : ClkMux
    port map (
            O => \N__62109\,
            I => \N__62071\
        );

    \I__13588\ : ClkMux
    port map (
            O => \N__62108\,
            I => \N__62071\
        );

    \I__13587\ : ClkMux
    port map (
            O => \N__62107\,
            I => \N__62071\
        );

    \I__13586\ : ClkMux
    port map (
            O => \N__62106\,
            I => \N__62071\
        );

    \I__13585\ : ClkMux
    port map (
            O => \N__62105\,
            I => \N__62071\
        );

    \I__13584\ : ClkMux
    port map (
            O => \N__62104\,
            I => \N__62071\
        );

    \I__13583\ : GlobalMux
    port map (
            O => \N__62071\,
            I => \N__62068\
        );

    \I__13582\ : gio2CtrlBuf
    port map (
            O => \N__62068\,
            I => \pin3_clk_16mhz_N\
        );

    \I__13581\ : InMux
    port map (
            O => \N__62065\,
            I => \N__62061\
        );

    \I__13580\ : CascadeMux
    port map (
            O => \N__62064\,
            I => \N__62057\
        );

    \I__13579\ : LocalMux
    port map (
            O => \N__62061\,
            I => \N__62054\
        );

    \I__13578\ : InMux
    port map (
            O => \N__62060\,
            I => \N__62051\
        );

    \I__13577\ : InMux
    port map (
            O => \N__62057\,
            I => \N__62048\
        );

    \I__13576\ : Span4Mux_v
    port map (
            O => \N__62054\,
            I => \N__62045\
        );

    \I__13575\ : LocalMux
    port map (
            O => \N__62051\,
            I => \N__62040\
        );

    \I__13574\ : LocalMux
    port map (
            O => \N__62048\,
            I => \N__62040\
        );

    \I__13573\ : Odrv4
    port map (
            O => \N__62045\,
            I => \Add_add_temp_25\
        );

    \I__13572\ : Odrv12
    port map (
            O => \N__62040\,
            I => \Add_add_temp_25\
        );

    \I__13571\ : InMux
    port map (
            O => \N__62035\,
            I => \N__62032\
        );

    \I__13570\ : LocalMux
    port map (
            O => \N__62032\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_5\
        );

    \I__13569\ : InMux
    port map (
            O => \N__62029\,
            I => \N__61998\
        );

    \I__13568\ : InMux
    port map (
            O => \N__62028\,
            I => \N__61998\
        );

    \I__13567\ : InMux
    port map (
            O => \N__62027\,
            I => \N__61998\
        );

    \I__13566\ : InMux
    port map (
            O => \N__62026\,
            I => \N__61998\
        );

    \I__13565\ : InMux
    port map (
            O => \N__62025\,
            I => \N__61998\
        );

    \I__13564\ : InMux
    port map (
            O => \N__62024\,
            I => \N__61998\
        );

    \I__13563\ : InMux
    port map (
            O => \N__62023\,
            I => \N__61998\
        );

    \I__13562\ : InMux
    port map (
            O => \N__62022\,
            I => \N__61998\
        );

    \I__13561\ : InMux
    port map (
            O => \N__62021\,
            I => \N__61987\
        );

    \I__13560\ : InMux
    port map (
            O => \N__62020\,
            I => \N__61987\
        );

    \I__13559\ : InMux
    port map (
            O => \N__62019\,
            I => \N__61987\
        );

    \I__13558\ : InMux
    port map (
            O => \N__62018\,
            I => \N__61987\
        );

    \I__13557\ : InMux
    port map (
            O => \N__62017\,
            I => \N__61987\
        );

    \I__13556\ : CascadeMux
    port map (
            O => \N__62016\,
            I => \N__61982\
        );

    \I__13555\ : CascadeMux
    port map (
            O => \N__62015\,
            I => \N__61978\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__61998\,
            I => \N__61961\
        );

    \I__13553\ : LocalMux
    port map (
            O => \N__61987\,
            I => \N__61961\
        );

    \I__13552\ : InMux
    port map (
            O => \N__61986\,
            I => \N__61956\
        );

    \I__13551\ : InMux
    port map (
            O => \N__61985\,
            I => \N__61956\
        );

    \I__13550\ : InMux
    port map (
            O => \N__61982\,
            I => \N__61943\
        );

    \I__13549\ : InMux
    port map (
            O => \N__61981\,
            I => \N__61943\
        );

    \I__13548\ : InMux
    port map (
            O => \N__61978\,
            I => \N__61943\
        );

    \I__13547\ : InMux
    port map (
            O => \N__61977\,
            I => \N__61943\
        );

    \I__13546\ : InMux
    port map (
            O => \N__61976\,
            I => \N__61943\
        );

    \I__13545\ : InMux
    port map (
            O => \N__61975\,
            I => \N__61943\
        );

    \I__13544\ : InMux
    port map (
            O => \N__61974\,
            I => \N__61934\
        );

    \I__13543\ : InMux
    port map (
            O => \N__61973\,
            I => \N__61934\
        );

    \I__13542\ : InMux
    port map (
            O => \N__61972\,
            I => \N__61934\
        );

    \I__13541\ : InMux
    port map (
            O => \N__61971\,
            I => \N__61934\
        );

    \I__13540\ : InMux
    port map (
            O => \N__61970\,
            I => \N__61923\
        );

    \I__13539\ : InMux
    port map (
            O => \N__61969\,
            I => \N__61923\
        );

    \I__13538\ : InMux
    port map (
            O => \N__61968\,
            I => \N__61923\
        );

    \I__13537\ : InMux
    port map (
            O => \N__61967\,
            I => \N__61923\
        );

    \I__13536\ : InMux
    port map (
            O => \N__61966\,
            I => \N__61923\
        );

    \I__13535\ : Odrv4
    port map (
            O => \N__61961\,
            I => \Saturate_out1_31__N_267\
        );

    \I__13534\ : LocalMux
    port map (
            O => \N__61956\,
            I => \Saturate_out1_31__N_267\
        );

    \I__13533\ : LocalMux
    port map (
            O => \N__61943\,
            I => \Saturate_out1_31__N_267\
        );

    \I__13532\ : LocalMux
    port map (
            O => \N__61934\,
            I => \Saturate_out1_31__N_267\
        );

    \I__13531\ : LocalMux
    port map (
            O => \N__61923\,
            I => \Saturate_out1_31__N_267\
        );

    \I__13530\ : InMux
    port map (
            O => \N__61912\,
            I => \N__61878\
        );

    \I__13529\ : InMux
    port map (
            O => \N__61911\,
            I => \N__61878\
        );

    \I__13528\ : InMux
    port map (
            O => \N__61910\,
            I => \N__61869\
        );

    \I__13527\ : InMux
    port map (
            O => \N__61909\,
            I => \N__61869\
        );

    \I__13526\ : InMux
    port map (
            O => \N__61908\,
            I => \N__61869\
        );

    \I__13525\ : InMux
    port map (
            O => \N__61907\,
            I => \N__61869\
        );

    \I__13524\ : InMux
    port map (
            O => \N__61906\,
            I => \N__61856\
        );

    \I__13523\ : InMux
    port map (
            O => \N__61905\,
            I => \N__61856\
        );

    \I__13522\ : InMux
    port map (
            O => \N__61904\,
            I => \N__61856\
        );

    \I__13521\ : InMux
    port map (
            O => \N__61903\,
            I => \N__61856\
        );

    \I__13520\ : InMux
    port map (
            O => \N__61902\,
            I => \N__61856\
        );

    \I__13519\ : InMux
    port map (
            O => \N__61901\,
            I => \N__61856\
        );

    \I__13518\ : InMux
    port map (
            O => \N__61900\,
            I => \N__61839\
        );

    \I__13517\ : InMux
    port map (
            O => \N__61899\,
            I => \N__61839\
        );

    \I__13516\ : InMux
    port map (
            O => \N__61898\,
            I => \N__61839\
        );

    \I__13515\ : InMux
    port map (
            O => \N__61897\,
            I => \N__61839\
        );

    \I__13514\ : InMux
    port map (
            O => \N__61896\,
            I => \N__61839\
        );

    \I__13513\ : InMux
    port map (
            O => \N__61895\,
            I => \N__61839\
        );

    \I__13512\ : InMux
    port map (
            O => \N__61894\,
            I => \N__61839\
        );

    \I__13511\ : InMux
    port map (
            O => \N__61893\,
            I => \N__61839\
        );

    \I__13510\ : InMux
    port map (
            O => \N__61892\,
            I => \N__61834\
        );

    \I__13509\ : InMux
    port map (
            O => \N__61891\,
            I => \N__61834\
        );

    \I__13508\ : InMux
    port map (
            O => \N__61890\,
            I => \N__61827\
        );

    \I__13507\ : InMux
    port map (
            O => \N__61889\,
            I => \N__61827\
        );

    \I__13506\ : InMux
    port map (
            O => \N__61888\,
            I => \N__61827\
        );

    \I__13505\ : InMux
    port map (
            O => \N__61887\,
            I => \N__61822\
        );

    \I__13504\ : InMux
    port map (
            O => \N__61886\,
            I => \N__61822\
        );

    \I__13503\ : InMux
    port map (
            O => \N__61885\,
            I => \N__61815\
        );

    \I__13502\ : InMux
    port map (
            O => \N__61884\,
            I => \N__61815\
        );

    \I__13501\ : InMux
    port map (
            O => \N__61883\,
            I => \N__61815\
        );

    \I__13500\ : LocalMux
    port map (
            O => \N__61878\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13499\ : LocalMux
    port map (
            O => \N__61869\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__61856\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13497\ : LocalMux
    port map (
            O => \N__61839\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13496\ : LocalMux
    port map (
            O => \N__61834\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13495\ : LocalMux
    port map (
            O => \N__61827\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13494\ : LocalMux
    port map (
            O => \N__61822\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13493\ : LocalMux
    port map (
            O => \N__61815\,
            I => \Saturate_out1_31__N_266\
        );

    \I__13492\ : CascadeMux
    port map (
            O => \N__61798\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19723_cascade_\
        );

    \I__13491\ : CascadeMux
    port map (
            O => \N__61795\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20708_cascade_\
        );

    \I__13490\ : CascadeMux
    port map (
            O => \N__61792\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n22_adj_519_cascade_\
        );

    \I__13489\ : InMux
    port map (
            O => \N__61789\,
            I => \N__61786\
        );

    \I__13488\ : LocalMux
    port map (
            O => \N__61786\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20688\
        );

    \I__13487\ : InMux
    port map (
            O => \N__61783\,
            I => \N__61780\
        );

    \I__13486\ : LocalMux
    port map (
            O => \N__61780\,
            I => \N__61777\
        );

    \I__13485\ : Span4Mux_h
    port map (
            O => \N__61777\,
            I => \N__61772\
        );

    \I__13484\ : InMux
    port map (
            O => \N__61776\,
            I => \N__61767\
        );

    \I__13483\ : InMux
    port map (
            O => \N__61775\,
            I => \N__61767\
        );

    \I__13482\ : Odrv4
    port map (
            O => \N__61772\,
            I => \Add_add_temp_17\
        );

    \I__13481\ : LocalMux
    port map (
            O => \N__61767\,
            I => \Add_add_temp_17\
        );

    \I__13480\ : InMux
    port map (
            O => \N__61762\,
            I => \N__61759\
        );

    \I__13479\ : LocalMux
    port map (
            O => \N__61759\,
            I => \N__61755\
        );

    \I__13478\ : CascadeMux
    port map (
            O => \N__61758\,
            I => \N__61751\
        );

    \I__13477\ : Span4Mux_v
    port map (
            O => \N__61755\,
            I => \N__61748\
        );

    \I__13476\ : InMux
    port map (
            O => \N__61754\,
            I => \N__61743\
        );

    \I__13475\ : InMux
    port map (
            O => \N__61751\,
            I => \N__61743\
        );

    \I__13474\ : Odrv4
    port map (
            O => \N__61748\,
            I => \Add_add_temp_16\
        );

    \I__13473\ : LocalMux
    port map (
            O => \N__61743\,
            I => \Add_add_temp_16\
        );

    \I__13472\ : InMux
    port map (
            O => \N__61738\,
            I => \N__61735\
        );

    \I__13471\ : LocalMux
    port map (
            O => \N__61735\,
            I => \N__61732\
        );

    \I__13470\ : Span4Mux_h
    port map (
            O => \N__61732\,
            I => \N__61727\
        );

    \I__13469\ : InMux
    port map (
            O => \N__61731\,
            I => \N__61722\
        );

    \I__13468\ : InMux
    port map (
            O => \N__61730\,
            I => \N__61722\
        );

    \I__13467\ : Odrv4
    port map (
            O => \N__61727\,
            I => \Add_add_temp_15\
        );

    \I__13466\ : LocalMux
    port map (
            O => \N__61722\,
            I => \Add_add_temp_15\
        );

    \I__13465\ : InMux
    port map (
            O => \N__61717\,
            I => \N__61713\
        );

    \I__13464\ : CascadeMux
    port map (
            O => \N__61716\,
            I => \N__61709\
        );

    \I__13463\ : LocalMux
    port map (
            O => \N__61713\,
            I => \N__61706\
        );

    \I__13462\ : InMux
    port map (
            O => \N__61712\,
            I => \N__61703\
        );

    \I__13461\ : InMux
    port map (
            O => \N__61709\,
            I => \N__61700\
        );

    \I__13460\ : Span4Mux_v
    port map (
            O => \N__61706\,
            I => \N__61697\
        );

    \I__13459\ : LocalMux
    port map (
            O => \N__61703\,
            I => \N__61692\
        );

    \I__13458\ : LocalMux
    port map (
            O => \N__61700\,
            I => \N__61692\
        );

    \I__13457\ : Odrv4
    port map (
            O => \N__61697\,
            I => \Add_add_temp_31\
        );

    \I__13456\ : Odrv12
    port map (
            O => \N__61692\,
            I => \Add_add_temp_31\
        );

    \I__13455\ : InMux
    port map (
            O => \N__61687\,
            I => \N__61680\
        );

    \I__13454\ : InMux
    port map (
            O => \N__61686\,
            I => \N__61680\
        );

    \I__13453\ : InMux
    port map (
            O => \N__61685\,
            I => \N__61677\
        );

    \I__13452\ : LocalMux
    port map (
            O => \N__61680\,
            I => \N__61674\
        );

    \I__13451\ : LocalMux
    port map (
            O => \N__61677\,
            I => \N__61671\
        );

    \I__13450\ : Span4Mux_v
    port map (
            O => \N__61674\,
            I => \N__61668\
        );

    \I__13449\ : Span4Mux_v
    port map (
            O => \N__61671\,
            I => \N__61665\
        );

    \I__13448\ : Odrv4
    port map (
            O => \N__61668\,
            I => \Add_add_temp_32\
        );

    \I__13447\ : Odrv4
    port map (
            O => \N__61665\,
            I => \Add_add_temp_32\
        );

    \I__13446\ : CascadeMux
    port map (
            O => \N__61660\,
            I => \N__61657\
        );

    \I__13445\ : InMux
    port map (
            O => \N__61657\,
            I => \N__61650\
        );

    \I__13444\ : InMux
    port map (
            O => \N__61656\,
            I => \N__61650\
        );

    \I__13443\ : InMux
    port map (
            O => \N__61655\,
            I => \N__61647\
        );

    \I__13442\ : LocalMux
    port map (
            O => \N__61650\,
            I => \N__61642\
        );

    \I__13441\ : LocalMux
    port map (
            O => \N__61647\,
            I => \N__61642\
        );

    \I__13440\ : Span4Mux_v
    port map (
            O => \N__61642\,
            I => \N__61639\
        );

    \I__13439\ : Odrv4
    port map (
            O => \N__61639\,
            I => \Add_add_temp_30\
        );

    \I__13438\ : InMux
    port map (
            O => \N__61636\,
            I => \N__61633\
        );

    \I__13437\ : LocalMux
    port map (
            O => \N__61633\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20644\
        );

    \I__13436\ : InMux
    port map (
            O => \N__61630\,
            I => \N__61626\
        );

    \I__13435\ : InMux
    port map (
            O => \N__61629\,
            I => \N__61623\
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__61626\,
            I => \N__61619\
        );

    \I__13433\ : LocalMux
    port map (
            O => \N__61623\,
            I => \N__61616\
        );

    \I__13432\ : InMux
    port map (
            O => \N__61622\,
            I => \N__61613\
        );

    \I__13431\ : Span4Mux_v
    port map (
            O => \N__61619\,
            I => \N__61610\
        );

    \I__13430\ : Span12Mux_s10_h
    port map (
            O => \N__61616\,
            I => \N__61605\
        );

    \I__13429\ : LocalMux
    port map (
            O => \N__61613\,
            I => \N__61605\
        );

    \I__13428\ : Odrv4
    port map (
            O => \N__61610\,
            I => \Add_add_temp_34\
        );

    \I__13427\ : Odrv12
    port map (
            O => \N__61605\,
            I => \Add_add_temp_34\
        );

    \I__13426\ : CascadeMux
    port map (
            O => \N__61600\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n58_cascade_\
        );

    \I__13425\ : InMux
    port map (
            O => \N__61597\,
            I => \N__61593\
        );

    \I__13424\ : InMux
    port map (
            O => \N__61596\,
            I => \N__61589\
        );

    \I__13423\ : LocalMux
    port map (
            O => \N__61593\,
            I => \N__61586\
        );

    \I__13422\ : InMux
    port map (
            O => \N__61592\,
            I => \N__61583\
        );

    \I__13421\ : LocalMux
    port map (
            O => \N__61589\,
            I => \N__61580\
        );

    \I__13420\ : Span4Mux_v
    port map (
            O => \N__61586\,
            I => \N__61575\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__61583\,
            I => \N__61575\
        );

    \I__13418\ : Span4Mux_h
    port map (
            O => \N__61580\,
            I => \N__61570\
        );

    \I__13417\ : Span4Mux_h
    port map (
            O => \N__61575\,
            I => \N__61570\
        );

    \I__13416\ : Span4Mux_v
    port map (
            O => \N__61570\,
            I => \N__61567\
        );

    \I__13415\ : Odrv4
    port map (
            O => \N__61567\,
            I => \Add_add_temp_33\
        );

    \I__13414\ : CascadeMux
    port map (
            O => \N__61564\,
            I => \Saturate_out1_31__N_266_cascade_\
        );

    \I__13413\ : InMux
    port map (
            O => \N__61561\,
            I => \N__61558\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__61558\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_4\
        );

    \I__13411\ : InMux
    port map (
            O => \N__61555\,
            I => \N__61552\
        );

    \I__13410\ : LocalMux
    port map (
            O => \N__61552\,
            I => \N__61547\
        );

    \I__13409\ : InMux
    port map (
            O => \N__61551\,
            I => \N__61542\
        );

    \I__13408\ : InMux
    port map (
            O => \N__61550\,
            I => \N__61542\
        );

    \I__13407\ : Span4Mux_v
    port map (
            O => \N__61547\,
            I => \N__61539\
        );

    \I__13406\ : LocalMux
    port map (
            O => \N__61542\,
            I => \N__61536\
        );

    \I__13405\ : Odrv4
    port map (
            O => \N__61539\,
            I => \Add_add_temp_26\
        );

    \I__13404\ : Odrv12
    port map (
            O => \N__61536\,
            I => \Add_add_temp_26\
        );

    \I__13403\ : InMux
    port map (
            O => \N__61531\,
            I => \N__61526\
        );

    \I__13402\ : InMux
    port map (
            O => \N__61530\,
            I => \N__61521\
        );

    \I__13401\ : InMux
    port map (
            O => \N__61529\,
            I => \N__61521\
        );

    \I__13400\ : LocalMux
    port map (
            O => \N__61526\,
            I => \N__61516\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__61521\,
            I => \N__61516\
        );

    \I__13398\ : Span4Mux_v
    port map (
            O => \N__61516\,
            I => \N__61513\
        );

    \I__13397\ : Odrv4
    port map (
            O => \N__61513\,
            I => \Add_add_temp_27\
        );

    \I__13396\ : CascadeMux
    port map (
            O => \N__61510\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n22_cascade_\
        );

    \I__13395\ : CascadeMux
    port map (
            O => \N__61507\,
            I => \foc.dVoltage_13_cascade_\
        );

    \I__13394\ : CascadeMux
    port map (
            O => \N__61504\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20568_cascade_\
        );

    \I__13393\ : InMux
    port map (
            O => \N__61501\,
            I => \N__61498\
        );

    \I__13392\ : LocalMux
    port map (
            O => \N__61498\,
            I => \N__61495\
        );

    \I__13391\ : Odrv4
    port map (
            O => \N__61495\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20576\
        );

    \I__13390\ : InMux
    port map (
            O => \N__61492\,
            I => \N__61489\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__61489\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n14\
        );

    \I__13388\ : InMux
    port map (
            O => \N__61486\,
            I => \N__61483\
        );

    \I__13387\ : LocalMux
    port map (
            O => \N__61483\,
            I => \foc.dVoltage_6\
        );

    \I__13386\ : CascadeMux
    port map (
            O => \N__61480\,
            I => \N__61472\
        );

    \I__13385\ : CascadeMux
    port map (
            O => \N__61479\,
            I => \N__61466\
        );

    \I__13384\ : CascadeMux
    port map (
            O => \N__61478\,
            I => \N__61463\
        );

    \I__13383\ : InMux
    port map (
            O => \N__61477\,
            I => \N__61455\
        );

    \I__13382\ : CascadeMux
    port map (
            O => \N__61476\,
            I => \N__61451\
        );

    \I__13381\ : CascadeMux
    port map (
            O => \N__61475\,
            I => \N__61446\
        );

    \I__13380\ : InMux
    port map (
            O => \N__61472\,
            I => \N__61437\
        );

    \I__13379\ : InMux
    port map (
            O => \N__61471\,
            I => \N__61437\
        );

    \I__13378\ : InMux
    port map (
            O => \N__61470\,
            I => \N__61437\
        );

    \I__13377\ : InMux
    port map (
            O => \N__61469\,
            I => \N__61437\
        );

    \I__13376\ : InMux
    port map (
            O => \N__61466\,
            I => \N__61426\
        );

    \I__13375\ : InMux
    port map (
            O => \N__61463\,
            I => \N__61426\
        );

    \I__13374\ : InMux
    port map (
            O => \N__61462\,
            I => \N__61426\
        );

    \I__13373\ : InMux
    port map (
            O => \N__61461\,
            I => \N__61426\
        );

    \I__13372\ : InMux
    port map (
            O => \N__61460\,
            I => \N__61426\
        );

    \I__13371\ : InMux
    port map (
            O => \N__61459\,
            I => \N__61421\
        );

    \I__13370\ : InMux
    port map (
            O => \N__61458\,
            I => \N__61421\
        );

    \I__13369\ : LocalMux
    port map (
            O => \N__61455\,
            I => \N__61418\
        );

    \I__13368\ : InMux
    port map (
            O => \N__61454\,
            I => \N__61415\
        );

    \I__13367\ : InMux
    port map (
            O => \N__61451\,
            I => \N__61412\
        );

    \I__13366\ : InMux
    port map (
            O => \N__61450\,
            I => \N__61405\
        );

    \I__13365\ : InMux
    port map (
            O => \N__61449\,
            I => \N__61405\
        );

    \I__13364\ : InMux
    port map (
            O => \N__61446\,
            I => \N__61405\
        );

    \I__13363\ : LocalMux
    port map (
            O => \N__61437\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__61426\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13361\ : LocalMux
    port map (
            O => \N__61421\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13360\ : Odrv12
    port map (
            O => \N__61418\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13359\ : LocalMux
    port map (
            O => \N__61415\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13358\ : LocalMux
    port map (
            O => \N__61412\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__61405\,
            I => \foc.Out_31__N_332_adj_2312\
        );

    \I__13356\ : CascadeMux
    port map (
            O => \N__61390\,
            I => \N__61383\
        );

    \I__13355\ : InMux
    port map (
            O => \N__61389\,
            I => \N__61368\
        );

    \I__13354\ : InMux
    port map (
            O => \N__61388\,
            I => \N__61365\
        );

    \I__13353\ : InMux
    port map (
            O => \N__61387\,
            I => \N__61356\
        );

    \I__13352\ : InMux
    port map (
            O => \N__61386\,
            I => \N__61356\
        );

    \I__13351\ : InMux
    port map (
            O => \N__61383\,
            I => \N__61356\
        );

    \I__13350\ : InMux
    port map (
            O => \N__61382\,
            I => \N__61356\
        );

    \I__13349\ : InMux
    port map (
            O => \N__61381\,
            I => \N__61347\
        );

    \I__13348\ : InMux
    port map (
            O => \N__61380\,
            I => \N__61347\
        );

    \I__13347\ : InMux
    port map (
            O => \N__61379\,
            I => \N__61347\
        );

    \I__13346\ : InMux
    port map (
            O => \N__61378\,
            I => \N__61347\
        );

    \I__13345\ : InMux
    port map (
            O => \N__61377\,
            I => \N__61336\
        );

    \I__13344\ : InMux
    port map (
            O => \N__61376\,
            I => \N__61336\
        );

    \I__13343\ : InMux
    port map (
            O => \N__61375\,
            I => \N__61336\
        );

    \I__13342\ : InMux
    port map (
            O => \N__61374\,
            I => \N__61336\
        );

    \I__13341\ : InMux
    port map (
            O => \N__61373\,
            I => \N__61336\
        );

    \I__13340\ : InMux
    port map (
            O => \N__61372\,
            I => \N__61331\
        );

    \I__13339\ : InMux
    port map (
            O => \N__61371\,
            I => \N__61331\
        );

    \I__13338\ : LocalMux
    port map (
            O => \N__61368\,
            I => \foc.Out_31__N_333_adj_2310\
        );

    \I__13337\ : LocalMux
    port map (
            O => \N__61365\,
            I => \foc.Out_31__N_333_adj_2310\
        );

    \I__13336\ : LocalMux
    port map (
            O => \N__61356\,
            I => \foc.Out_31__N_333_adj_2310\
        );

    \I__13335\ : LocalMux
    port map (
            O => \N__61347\,
            I => \foc.Out_31__N_333_adj_2310\
        );

    \I__13334\ : LocalMux
    port map (
            O => \N__61336\,
            I => \foc.Out_31__N_333_adj_2310\
        );

    \I__13333\ : LocalMux
    port map (
            O => \N__61331\,
            I => \foc.Out_31__N_333_adj_2310\
        );

    \I__13332\ : InMux
    port map (
            O => \N__61318\,
            I => \N__61315\
        );

    \I__13331\ : LocalMux
    port map (
            O => \N__61315\,
            I => \foc.dVoltage_7\
        );

    \I__13330\ : InMux
    port map (
            O => \N__61312\,
            I => \N__61309\
        );

    \I__13329\ : LocalMux
    port map (
            O => \N__61309\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19747\
        );

    \I__13328\ : InMux
    port map (
            O => \N__61306\,
            I => \N__61303\
        );

    \I__13327\ : LocalMux
    port map (
            O => \N__61303\,
            I => \N__61300\
        );

    \I__13326\ : Span4Mux_v
    port map (
            O => \N__61300\,
            I => \N__61297\
        );

    \I__13325\ : Odrv4
    port map (
            O => \N__61297\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19858\
        );

    \I__13324\ : InMux
    port map (
            O => \N__61294\,
            I => \N__61291\
        );

    \I__13323\ : LocalMux
    port map (
            O => \N__61291\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19904\
        );

    \I__13322\ : InMux
    port map (
            O => \N__61288\,
            I => \N__61285\
        );

    \I__13321\ : LocalMux
    port map (
            O => \N__61285\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n446\
        );

    \I__13320\ : InMux
    port map (
            O => \N__61282\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17529\
        );

    \I__13319\ : InMux
    port map (
            O => \N__61279\,
            I => \N__61276\
        );

    \I__13318\ : LocalMux
    port map (
            O => \N__61276\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n495\
        );

    \I__13317\ : InMux
    port map (
            O => \N__61273\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17530\
        );

    \I__13316\ : InMux
    port map (
            O => \N__61270\,
            I => \N__61267\
        );

    \I__13315\ : LocalMux
    port map (
            O => \N__61267\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n544\
        );

    \I__13314\ : InMux
    port map (
            O => \N__61264\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17531\
        );

    \I__13313\ : InMux
    port map (
            O => \N__61261\,
            I => \N__61258\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__61258\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n593\
        );

    \I__13311\ : InMux
    port map (
            O => \N__61255\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17532\
        );

    \I__13310\ : InMux
    port map (
            O => \N__61252\,
            I => \N__61249\
        );

    \I__13309\ : LocalMux
    port map (
            O => \N__61249\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n642\
        );

    \I__13308\ : InMux
    port map (
            O => \N__61246\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17533\
        );

    \I__13307\ : InMux
    port map (
            O => \N__61243\,
            I => \N__61240\
        );

    \I__13306\ : LocalMux
    port map (
            O => \N__61240\,
            I => \N__61237\
        );

    \I__13305\ : Span4Mux_v
    port map (
            O => \N__61237\,
            I => \N__61233\
        );

    \I__13304\ : InMux
    port map (
            O => \N__61236\,
            I => \N__61230\
        );

    \I__13303\ : Span4Mux_h
    port map (
            O => \N__61233\,
            I => \N__61227\
        );

    \I__13302\ : LocalMux
    port map (
            O => \N__61230\,
            I => \N__61224\
        );

    \I__13301\ : Span4Mux_v
    port map (
            O => \N__61227\,
            I => \N__61221\
        );

    \I__13300\ : Span4Mux_v
    port map (
            O => \N__61224\,
            I => \N__61218\
        );

    \I__13299\ : Odrv4
    port map (
            O => \N__61221\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n737\
        );

    \I__13298\ : Odrv4
    port map (
            O => \N__61218\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n737\
        );

    \I__13297\ : CascadeMux
    port map (
            O => \N__61213\,
            I => \N__61210\
        );

    \I__13296\ : InMux
    port map (
            O => \N__61210\,
            I => \N__61207\
        );

    \I__13295\ : LocalMux
    port map (
            O => \N__61207\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n691_adj_440\
        );

    \I__13294\ : CascadeMux
    port map (
            O => \N__61204\,
            I => \N__61201\
        );

    \I__13293\ : InMux
    port map (
            O => \N__61201\,
            I => \N__61197\
        );

    \I__13292\ : InMux
    port map (
            O => \N__61200\,
            I => \N__61194\
        );

    \I__13291\ : LocalMux
    port map (
            O => \N__61197\,
            I => \N__61189\
        );

    \I__13290\ : LocalMux
    port map (
            O => \N__61194\,
            I => \N__61189\
        );

    \I__13289\ : Span4Mux_h
    port map (
            O => \N__61189\,
            I => \N__61186\
        );

    \I__13288\ : Odrv4
    port map (
            O => \N__61186\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n738\
        );

    \I__13287\ : InMux
    port map (
            O => \N__61183\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17534\
        );

    \I__13286\ : InMux
    port map (
            O => \N__61180\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n739\
        );

    \I__13285\ : CascadeMux
    port map (
            O => \N__61177\,
            I => \N__61174\
        );

    \I__13284\ : InMux
    port map (
            O => \N__61174\,
            I => \N__61171\
        );

    \I__13283\ : LocalMux
    port map (
            O => \N__61171\,
            I => \N__61168\
        );

    \I__13282\ : Span4Mux_v
    port map (
            O => \N__61168\,
            I => \N__61165\
        );

    \I__13281\ : Odrv4
    port map (
            O => \N__61165\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_CO\
        );

    \I__13280\ : InMux
    port map (
            O => \N__61162\,
            I => \N__61159\
        );

    \I__13279\ : LocalMux
    port map (
            O => \N__61159\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19932\
        );

    \I__13278\ : InMux
    port map (
            O => \N__61156\,
            I => \N__61153\
        );

    \I__13277\ : LocalMux
    port map (
            O => \N__61153\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20546\
        );

    \I__13276\ : CascadeMux
    port map (
            O => \N__61150\,
            I => \N__61147\
        );

    \I__13275\ : InMux
    port map (
            O => \N__61147\,
            I => \N__61144\
        );

    \I__13274\ : LocalMux
    port map (
            O => \N__61144\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n54\
        );

    \I__13273\ : InMux
    port map (
            O => \N__61141\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17521\
        );

    \I__13272\ : InMux
    port map (
            O => \N__61138\,
            I => \N__61135\
        );

    \I__13271\ : LocalMux
    port map (
            O => \N__61135\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n103\
        );

    \I__13270\ : InMux
    port map (
            O => \N__61132\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17522\
        );

    \I__13269\ : CascadeMux
    port map (
            O => \N__61129\,
            I => \N__61126\
        );

    \I__13268\ : InMux
    port map (
            O => \N__61126\,
            I => \N__61123\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__61123\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n152\
        );

    \I__13266\ : InMux
    port map (
            O => \N__61120\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17523\
        );

    \I__13265\ : InMux
    port map (
            O => \N__61117\,
            I => \N__61114\
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__61114\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n201\
        );

    \I__13263\ : InMux
    port map (
            O => \N__61111\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17524\
        );

    \I__13262\ : CascadeMux
    port map (
            O => \N__61108\,
            I => \N__61105\
        );

    \I__13261\ : InMux
    port map (
            O => \N__61105\,
            I => \N__61102\
        );

    \I__13260\ : LocalMux
    port map (
            O => \N__61102\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n250\
        );

    \I__13259\ : InMux
    port map (
            O => \N__61099\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17525\
        );

    \I__13258\ : InMux
    port map (
            O => \N__61096\,
            I => \N__61093\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__61093\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n299\
        );

    \I__13256\ : InMux
    port map (
            O => \N__61090\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17526\
        );

    \I__13255\ : CascadeMux
    port map (
            O => \N__61087\,
            I => \N__61084\
        );

    \I__13254\ : InMux
    port map (
            O => \N__61084\,
            I => \N__61081\
        );

    \I__13253\ : LocalMux
    port map (
            O => \N__61081\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n348\
        );

    \I__13252\ : InMux
    port map (
            O => \N__61078\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17527\
        );

    \I__13251\ : CascadeMux
    port map (
            O => \N__61075\,
            I => \N__61072\
        );

    \I__13250\ : InMux
    port map (
            O => \N__61072\,
            I => \N__61069\
        );

    \I__13249\ : LocalMux
    port map (
            O => \N__61069\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n397\
        );

    \I__13248\ : InMux
    port map (
            O => \N__61066\,
            I => \bfn_23_12_0_\
        );

    \I__13247\ : InMux
    port map (
            O => \N__61063\,
            I => \N__61060\
        );

    \I__13246\ : LocalMux
    port map (
            O => \N__61060\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n470_adj_594\
        );

    \I__13245\ : InMux
    port map (
            O => \N__61057\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18287\
        );

    \I__13244\ : InMux
    port map (
            O => \N__61054\,
            I => \N__61051\
        );

    \I__13243\ : LocalMux
    port map (
            O => \N__61051\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n519_adj_593\
        );

    \I__13242\ : InMux
    port map (
            O => \N__61048\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18288\
        );

    \I__13241\ : InMux
    port map (
            O => \N__61045\,
            I => \N__61042\
        );

    \I__13240\ : LocalMux
    port map (
            O => \N__61042\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n568_adj_592\
        );

    \I__13239\ : InMux
    port map (
            O => \N__61039\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18289\
        );

    \I__13238\ : InMux
    port map (
            O => \N__61036\,
            I => \N__61033\
        );

    \I__13237\ : LocalMux
    port map (
            O => \N__61033\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n617_adj_591\
        );

    \I__13236\ : InMux
    port map (
            O => \N__61030\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18290\
        );

    \I__13235\ : CascadeMux
    port map (
            O => \N__61027\,
            I => \N__61024\
        );

    \I__13234\ : InMux
    port map (
            O => \N__61024\,
            I => \N__61021\
        );

    \I__13233\ : LocalMux
    port map (
            O => \N__61021\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n666\
        );

    \I__13232\ : InMux
    port map (
            O => \N__61018\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18291\
        );

    \I__13231\ : CascadeMux
    port map (
            O => \N__61015\,
            I => \N__61012\
        );

    \I__13230\ : InMux
    port map (
            O => \N__61012\,
            I => \N__61009\
        );

    \I__13229\ : LocalMux
    port map (
            O => \N__61009\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n715\
        );

    \I__13228\ : InMux
    port map (
            O => \N__61006\,
            I => \N__61003\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__61003\,
            I => \N__61000\
        );

    \I__13226\ : Span4Mux_h
    port map (
            O => \N__61000\,
            I => \N__60997\
        );

    \I__13225\ : Span4Mux_v
    port map (
            O => \N__60997\,
            I => \N__60994\
        );

    \I__13224\ : Odrv4
    port map (
            O => \N__60994\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n770\
        );

    \I__13223\ : InMux
    port map (
            O => \N__60991\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18292\
        );

    \I__13222\ : InMux
    port map (
            O => \N__60988\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771\
        );

    \I__13221\ : CascadeMux
    port map (
            O => \N__60985\,
            I => \N__60982\
        );

    \I__13220\ : InMux
    port map (
            O => \N__60982\,
            I => \N__60979\
        );

    \I__13219\ : LocalMux
    port map (
            O => \N__60979\,
            I => \N__60976\
        );

    \I__13218\ : Span4Mux_h
    port map (
            O => \N__60976\,
            I => \N__60973\
        );

    \I__13217\ : Span4Mux_v
    port map (
            O => \N__60973\,
            I => \N__60970\
        );

    \I__13216\ : Odrv4
    port map (
            O => \N__60970\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_CO\
        );

    \I__13215\ : InMux
    port map (
            O => \N__60967\,
            I => \N__60963\
        );

    \I__13214\ : InMux
    port map (
            O => \N__60966\,
            I => \N__60960\
        );

    \I__13213\ : LocalMux
    port map (
            O => \N__60963\,
            I => \N__60946\
        );

    \I__13212\ : LocalMux
    port map (
            O => \N__60960\,
            I => \N__60946\
        );

    \I__13211\ : InMux
    port map (
            O => \N__60959\,
            I => \N__60943\
        );

    \I__13210\ : InMux
    port map (
            O => \N__60958\,
            I => \N__60940\
        );

    \I__13209\ : CascadeMux
    port map (
            O => \N__60957\,
            I => \N__60935\
        );

    \I__13208\ : CascadeMux
    port map (
            O => \N__60956\,
            I => \N__60931\
        );

    \I__13207\ : CascadeMux
    port map (
            O => \N__60955\,
            I => \N__60927\
        );

    \I__13206\ : CascadeMux
    port map (
            O => \N__60954\,
            I => \N__60923\
        );

    \I__13205\ : CascadeMux
    port map (
            O => \N__60953\,
            I => \N__60919\
        );

    \I__13204\ : CascadeMux
    port map (
            O => \N__60952\,
            I => \N__60915\
        );

    \I__13203\ : CascadeMux
    port map (
            O => \N__60951\,
            I => \N__60911\
        );

    \I__13202\ : Span4Mux_v
    port map (
            O => \N__60946\,
            I => \N__60904\
        );

    \I__13201\ : LocalMux
    port map (
            O => \N__60943\,
            I => \N__60904\
        );

    \I__13200\ : LocalMux
    port map (
            O => \N__60940\,
            I => \N__60904\
        );

    \I__13199\ : InMux
    port map (
            O => \N__60939\,
            I => \N__60899\
        );

    \I__13198\ : InMux
    port map (
            O => \N__60938\,
            I => \N__60886\
        );

    \I__13197\ : InMux
    port map (
            O => \N__60935\,
            I => \N__60886\
        );

    \I__13196\ : InMux
    port map (
            O => \N__60934\,
            I => \N__60886\
        );

    \I__13195\ : InMux
    port map (
            O => \N__60931\,
            I => \N__60886\
        );

    \I__13194\ : InMux
    port map (
            O => \N__60930\,
            I => \N__60886\
        );

    \I__13193\ : InMux
    port map (
            O => \N__60927\,
            I => \N__60886\
        );

    \I__13192\ : InMux
    port map (
            O => \N__60926\,
            I => \N__60869\
        );

    \I__13191\ : InMux
    port map (
            O => \N__60923\,
            I => \N__60869\
        );

    \I__13190\ : InMux
    port map (
            O => \N__60922\,
            I => \N__60869\
        );

    \I__13189\ : InMux
    port map (
            O => \N__60919\,
            I => \N__60869\
        );

    \I__13188\ : InMux
    port map (
            O => \N__60918\,
            I => \N__60869\
        );

    \I__13187\ : InMux
    port map (
            O => \N__60915\,
            I => \N__60869\
        );

    \I__13186\ : InMux
    port map (
            O => \N__60914\,
            I => \N__60869\
        );

    \I__13185\ : InMux
    port map (
            O => \N__60911\,
            I => \N__60869\
        );

    \I__13184\ : Span4Mux_v
    port map (
            O => \N__60904\,
            I => \N__60866\
        );

    \I__13183\ : InMux
    port map (
            O => \N__60903\,
            I => \N__60863\
        );

    \I__13182\ : InMux
    port map (
            O => \N__60902\,
            I => \N__60859\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__60899\,
            I => \N__60853\
        );

    \I__13180\ : LocalMux
    port map (
            O => \N__60886\,
            I => \N__60848\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__60869\,
            I => \N__60848\
        );

    \I__13178\ : Span4Mux_h
    port map (
            O => \N__60866\,
            I => \N__60843\
        );

    \I__13177\ : LocalMux
    port map (
            O => \N__60863\,
            I => \N__60843\
        );

    \I__13176\ : CascadeMux
    port map (
            O => \N__60862\,
            I => \N__60840\
        );

    \I__13175\ : LocalMux
    port map (
            O => \N__60859\,
            I => \N__60836\
        );

    \I__13174\ : InMux
    port map (
            O => \N__60858\,
            I => \N__60833\
        );

    \I__13173\ : InMux
    port map (
            O => \N__60857\,
            I => \N__60830\
        );

    \I__13172\ : InMux
    port map (
            O => \N__60856\,
            I => \N__60825\
        );

    \I__13171\ : Span4Mux_v
    port map (
            O => \N__60853\,
            I => \N__60822\
        );

    \I__13170\ : Span4Mux_v
    port map (
            O => \N__60848\,
            I => \N__60817\
        );

    \I__13169\ : Span4Mux_v
    port map (
            O => \N__60843\,
            I => \N__60817\
        );

    \I__13168\ : InMux
    port map (
            O => \N__60840\,
            I => \N__60814\
        );

    \I__13167\ : InMux
    port map (
            O => \N__60839\,
            I => \N__60811\
        );

    \I__13166\ : Span4Mux_h
    port map (
            O => \N__60836\,
            I => \N__60806\
        );

    \I__13165\ : LocalMux
    port map (
            O => \N__60833\,
            I => \N__60806\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__60830\,
            I => \N__60803\
        );

    \I__13163\ : InMux
    port map (
            O => \N__60829\,
            I => \N__60800\
        );

    \I__13162\ : InMux
    port map (
            O => \N__60828\,
            I => \N__60797\
        );

    \I__13161\ : LocalMux
    port map (
            O => \N__60825\,
            I => \N__60793\
        );

    \I__13160\ : Sp12to4
    port map (
            O => \N__60822\,
            I => \N__60786\
        );

    \I__13159\ : Sp12to4
    port map (
            O => \N__60817\,
            I => \N__60786\
        );

    \I__13158\ : LocalMux
    port map (
            O => \N__60814\,
            I => \N__60786\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__60811\,
            I => \N__60783\
        );

    \I__13156\ : Span4Mux_v
    port map (
            O => \N__60806\,
            I => \N__60774\
        );

    \I__13155\ : Span4Mux_h
    port map (
            O => \N__60803\,
            I => \N__60774\
        );

    \I__13154\ : LocalMux
    port map (
            O => \N__60800\,
            I => \N__60774\
        );

    \I__13153\ : LocalMux
    port map (
            O => \N__60797\,
            I => \N__60774\
        );

    \I__13152\ : InMux
    port map (
            O => \N__60796\,
            I => \N__60771\
        );

    \I__13151\ : Span4Mux_v
    port map (
            O => \N__60793\,
            I => \N__60768\
        );

    \I__13150\ : Span12Mux_h
    port map (
            O => \N__60786\,
            I => \N__60765\
        );

    \I__13149\ : Span4Mux_h
    port map (
            O => \N__60783\,
            I => \N__60762\
        );

    \I__13148\ : Span4Mux_v
    port map (
            O => \N__60774\,
            I => \N__60757\
        );

    \I__13147\ : LocalMux
    port map (
            O => \N__60771\,
            I => \N__60757\
        );

    \I__13146\ : Odrv4
    port map (
            O => \N__60768\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n102\
        );

    \I__13145\ : Odrv12
    port map (
            O => \N__60765\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n102\
        );

    \I__13144\ : Odrv4
    port map (
            O => \N__60762\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n102\
        );

    \I__13143\ : Odrv4
    port map (
            O => \N__60757\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n102\
        );

    \I__13142\ : InMux
    port map (
            O => \N__60748\,
            I => \N__60745\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__60745\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n78\
        );

    \I__13140\ : InMux
    port map (
            O => \N__60742\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18279\
        );

    \I__13139\ : InMux
    port map (
            O => \N__60739\,
            I => \N__60736\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__60736\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n127\
        );

    \I__13137\ : InMux
    port map (
            O => \N__60733\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18280\
        );

    \I__13136\ : InMux
    port map (
            O => \N__60730\,
            I => \N__60727\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__60727\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n176\
        );

    \I__13134\ : InMux
    port map (
            O => \N__60724\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18281\
        );

    \I__13133\ : InMux
    port map (
            O => \N__60721\,
            I => \N__60718\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__60718\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n225\
        );

    \I__13131\ : InMux
    port map (
            O => \N__60715\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18282\
        );

    \I__13130\ : InMux
    port map (
            O => \N__60712\,
            I => \N__60709\
        );

    \I__13129\ : LocalMux
    port map (
            O => \N__60709\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n274\
        );

    \I__13128\ : InMux
    port map (
            O => \N__60706\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18283\
        );

    \I__13127\ : InMux
    port map (
            O => \N__60703\,
            I => \N__60700\
        );

    \I__13126\ : LocalMux
    port map (
            O => \N__60700\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n323\
        );

    \I__13125\ : InMux
    port map (
            O => \N__60697\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18284\
        );

    \I__13124\ : CascadeMux
    port map (
            O => \N__60694\,
            I => \N__60691\
        );

    \I__13123\ : InMux
    port map (
            O => \N__60691\,
            I => \N__60688\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__60688\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n372_adj_596\
        );

    \I__13121\ : InMux
    port map (
            O => \N__60685\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18285\
        );

    \I__13120\ : InMux
    port map (
            O => \N__60682\,
            I => \N__60679\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__60679\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n421_adj_595\
        );

    \I__13118\ : InMux
    port map (
            O => \N__60676\,
            I => \bfn_22_29_0_\
        );

    \I__13117\ : InMux
    port map (
            O => \N__60673\,
            I => \N__60670\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__60670\,
            I => \N__60667\
        );

    \I__13115\ : Odrv12
    port map (
            O => \N__60667\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n458\
        );

    \I__13114\ : InMux
    port map (
            O => \N__60664\,
            I => \bfn_22_26_0_\
        );

    \I__13113\ : InMux
    port map (
            O => \N__60661\,
            I => \N__60658\
        );

    \I__13112\ : LocalMux
    port map (
            O => \N__60658\,
            I => \N__60655\
        );

    \I__13111\ : Odrv12
    port map (
            O => \N__60655\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n507\
        );

    \I__13110\ : InMux
    port map (
            O => \N__60652\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18242\
        );

    \I__13109\ : InMux
    port map (
            O => \N__60649\,
            I => \N__60646\
        );

    \I__13108\ : LocalMux
    port map (
            O => \N__60646\,
            I => \N__60643\
        );

    \I__13107\ : Odrv12
    port map (
            O => \N__60643\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n556\
        );

    \I__13106\ : InMux
    port map (
            O => \N__60640\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18243\
        );

    \I__13105\ : InMux
    port map (
            O => \N__60637\,
            I => \N__60634\
        );

    \I__13104\ : LocalMux
    port map (
            O => \N__60634\,
            I => \N__60631\
        );

    \I__13103\ : Odrv12
    port map (
            O => \N__60631\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n605\
        );

    \I__13102\ : InMux
    port map (
            O => \N__60628\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18244\
        );

    \I__13101\ : CascadeMux
    port map (
            O => \N__60625\,
            I => \N__60622\
        );

    \I__13100\ : InMux
    port map (
            O => \N__60622\,
            I => \N__60619\
        );

    \I__13099\ : LocalMux
    port map (
            O => \N__60619\,
            I => \N__60616\
        );

    \I__13098\ : Odrv12
    port map (
            O => \N__60616\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n654\
        );

    \I__13097\ : InMux
    port map (
            O => \N__60613\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18245\
        );

    \I__13096\ : CascadeMux
    port map (
            O => \N__60610\,
            I => \N__60607\
        );

    \I__13095\ : InMux
    port map (
            O => \N__60607\,
            I => \N__60604\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__60604\,
            I => \N__60601\
        );

    \I__13093\ : Odrv4
    port map (
            O => \N__60601\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n703\
        );

    \I__13092\ : InMux
    port map (
            O => \N__60598\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18246\
        );

    \I__13091\ : InMux
    port map (
            O => \N__60595\,
            I => \N__60592\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__60592\,
            I => \N__60589\
        );

    \I__13089\ : Span4Mux_v
    port map (
            O => \N__60589\,
            I => \N__60586\
        );

    \I__13088\ : Span4Mux_v
    port map (
            O => \N__60586\,
            I => \N__60583\
        );

    \I__13087\ : Odrv4
    port map (
            O => \N__60583\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n758\
        );

    \I__13086\ : InMux
    port map (
            O => \N__60580\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18247\
        );

    \I__13085\ : InMux
    port map (
            O => \N__60577\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759\
        );

    \I__13084\ : CascadeMux
    port map (
            O => \N__60574\,
            I => \N__60571\
        );

    \I__13083\ : InMux
    port map (
            O => \N__60571\,
            I => \N__60568\
        );

    \I__13082\ : LocalMux
    port map (
            O => \N__60568\,
            I => \N__60565\
        );

    \I__13081\ : Span12Mux_h
    port map (
            O => \N__60565\,
            I => \N__60562\
        );

    \I__13080\ : Odrv12
    port map (
            O => \N__60562\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_CO\
        );

    \I__13079\ : CascadeMux
    port map (
            O => \N__60559\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19761_cascade_\
        );

    \I__13078\ : InMux
    port map (
            O => \N__60556\,
            I => \N__60553\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__60553\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20704\
        );

    \I__13076\ : InMux
    port map (
            O => \N__60550\,
            I => \N__60547\
        );

    \I__13075\ : LocalMux
    port map (
            O => \N__60547\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n69\
        );

    \I__13074\ : InMux
    port map (
            O => \N__60544\,
            I => \N__60541\
        );

    \I__13073\ : LocalMux
    port map (
            O => \N__60541\,
            I => \N__60538\
        );

    \I__13072\ : Odrv12
    port map (
            O => \N__60538\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n115\
        );

    \I__13071\ : InMux
    port map (
            O => \N__60535\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18234\
        );

    \I__13070\ : InMux
    port map (
            O => \N__60532\,
            I => \N__60529\
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__60529\,
            I => \N__60526\
        );

    \I__13068\ : Odrv12
    port map (
            O => \N__60526\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n164\
        );

    \I__13067\ : InMux
    port map (
            O => \N__60523\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18235\
        );

    \I__13066\ : InMux
    port map (
            O => \N__60520\,
            I => \N__60517\
        );

    \I__13065\ : LocalMux
    port map (
            O => \N__60517\,
            I => \N__60514\
        );

    \I__13064\ : Odrv12
    port map (
            O => \N__60514\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n213\
        );

    \I__13063\ : InMux
    port map (
            O => \N__60511\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18236\
        );

    \I__13062\ : InMux
    port map (
            O => \N__60508\,
            I => \N__60505\
        );

    \I__13061\ : LocalMux
    port map (
            O => \N__60505\,
            I => \N__60502\
        );

    \I__13060\ : Odrv12
    port map (
            O => \N__60502\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n262\
        );

    \I__13059\ : InMux
    port map (
            O => \N__60499\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18237\
        );

    \I__13058\ : CascadeMux
    port map (
            O => \N__60496\,
            I => \N__60493\
        );

    \I__13057\ : InMux
    port map (
            O => \N__60493\,
            I => \N__60490\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__60490\,
            I => \N__60487\
        );

    \I__13055\ : Odrv4
    port map (
            O => \N__60487\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n311\
        );

    \I__13054\ : InMux
    port map (
            O => \N__60484\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18238\
        );

    \I__13053\ : CascadeMux
    port map (
            O => \N__60481\,
            I => \N__60478\
        );

    \I__13052\ : InMux
    port map (
            O => \N__60478\,
            I => \N__60475\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__60475\,
            I => \N__60472\
        );

    \I__13050\ : Odrv12
    port map (
            O => \N__60472\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n360\
        );

    \I__13049\ : InMux
    port map (
            O => \N__60469\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18239\
        );

    \I__13048\ : InMux
    port map (
            O => \N__60466\,
            I => \N__60463\
        );

    \I__13047\ : LocalMux
    port map (
            O => \N__60463\,
            I => \N__60460\
        );

    \I__13046\ : Span4Mux_v
    port map (
            O => \N__60460\,
            I => \N__60457\
        );

    \I__13045\ : Odrv4
    port map (
            O => \N__60457\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n409\
        );

    \I__13044\ : InMux
    port map (
            O => \N__60454\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18240\
        );

    \I__13043\ : InMux
    port map (
            O => \N__60451\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n16002\
        );

    \I__13042\ : CascadeMux
    port map (
            O => \N__60448\,
            I => \N__60444\
        );

    \I__13041\ : CascadeMux
    port map (
            O => \N__60447\,
            I => \N__60438\
        );

    \I__13040\ : InMux
    port map (
            O => \N__60444\,
            I => \N__60433\
        );

    \I__13039\ : InMux
    port map (
            O => \N__60443\,
            I => \N__60433\
        );

    \I__13038\ : InMux
    port map (
            O => \N__60442\,
            I => \N__60426\
        );

    \I__13037\ : InMux
    port map (
            O => \N__60441\,
            I => \N__60426\
        );

    \I__13036\ : InMux
    port map (
            O => \N__60438\,
            I => \N__60426\
        );

    \I__13035\ : LocalMux
    port map (
            O => \N__60433\,
            I => \N__60421\
        );

    \I__13034\ : LocalMux
    port map (
            O => \N__60426\,
            I => \N__60421\
        );

    \I__13033\ : Span4Mux_v
    port map (
            O => \N__60421\,
            I => \N__60418\
        );

    \I__13032\ : Odrv4
    port map (
            O => \N__60418\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_31\
        );

    \I__13031\ : InMux
    port map (
            O => \N__60415\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n16003\
        );

    \I__13030\ : InMux
    port map (
            O => \N__60412\,
            I => \N__60408\
        );

    \I__13029\ : InMux
    port map (
            O => \N__60411\,
            I => \N__60405\
        );

    \I__13028\ : LocalMux
    port map (
            O => \N__60408\,
            I => \N__60402\
        );

    \I__13027\ : LocalMux
    port map (
            O => \N__60405\,
            I => \N__60399\
        );

    \I__13026\ : Span4Mux_h
    port map (
            O => \N__60402\,
            I => \N__60395\
        );

    \I__13025\ : Span12Mux_h
    port map (
            O => \N__60399\,
            I => \N__60392\
        );

    \I__13024\ : InMux
    port map (
            O => \N__60398\,
            I => \N__60389\
        );

    \I__13023\ : Odrv4
    port map (
            O => \N__60395\,
            I => \Add_add_temp_14_adj_2406\
        );

    \I__13022\ : Odrv12
    port map (
            O => \N__60392\,
            I => \Add_add_temp_14_adj_2406\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__60389\,
            I => \Add_add_temp_14_adj_2406\
        );

    \I__13020\ : InMux
    port map (
            O => \N__60382\,
            I => \N__60376\
        );

    \I__13019\ : InMux
    port map (
            O => \N__60381\,
            I => \N__60376\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__60376\,
            I => \N__60372\
        );

    \I__13017\ : CascadeMux
    port map (
            O => \N__60375\,
            I => \N__60369\
        );

    \I__13016\ : Span4Mux_v
    port map (
            O => \N__60372\,
            I => \N__60366\
        );

    \I__13015\ : InMux
    port map (
            O => \N__60369\,
            I => \N__60363\
        );

    \I__13014\ : Odrv4
    port map (
            O => \N__60366\,
            I => \Add_add_temp_12_adj_2408\
        );

    \I__13013\ : LocalMux
    port map (
            O => \N__60363\,
            I => \Add_add_temp_12_adj_2408\
        );

    \I__13012\ : InMux
    port map (
            O => \N__60358\,
            I => \N__60355\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__60355\,
            I => \N__60351\
        );

    \I__13010\ : CascadeMux
    port map (
            O => \N__60354\,
            I => \N__60348\
        );

    \I__13009\ : Span4Mux_h
    port map (
            O => \N__60351\,
            I => \N__60345\
        );

    \I__13008\ : InMux
    port map (
            O => \N__60348\,
            I => \N__60342\
        );

    \I__13007\ : Span4Mux_h
    port map (
            O => \N__60345\,
            I => \N__60336\
        );

    \I__13006\ : LocalMux
    port map (
            O => \N__60342\,
            I => \N__60336\
        );

    \I__13005\ : InMux
    port map (
            O => \N__60341\,
            I => \N__60333\
        );

    \I__13004\ : Odrv4
    port map (
            O => \N__60336\,
            I => \Add_add_temp_13_adj_2407\
        );

    \I__13003\ : LocalMux
    port map (
            O => \N__60333\,
            I => \Add_add_temp_13_adj_2407\
        );

    \I__13002\ : InMux
    port map (
            O => \N__60328\,
            I => \N__60322\
        );

    \I__13001\ : InMux
    port map (
            O => \N__60327\,
            I => \N__60322\
        );

    \I__13000\ : LocalMux
    port map (
            O => \N__60322\,
            I => \N__60318\
        );

    \I__12999\ : InMux
    port map (
            O => \N__60321\,
            I => \N__60315\
        );

    \I__12998\ : Odrv4
    port map (
            O => \N__60318\,
            I => \Add_add_temp_16_adj_2404\
        );

    \I__12997\ : LocalMux
    port map (
            O => \N__60315\,
            I => \Add_add_temp_16_adj_2404\
        );

    \I__12996\ : InMux
    port map (
            O => \N__60310\,
            I => \N__60304\
        );

    \I__12995\ : InMux
    port map (
            O => \N__60309\,
            I => \N__60304\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__60304\,
            I => \N__60300\
        );

    \I__12993\ : InMux
    port map (
            O => \N__60303\,
            I => \N__60297\
        );

    \I__12992\ : Odrv4
    port map (
            O => \N__60300\,
            I => \Add_add_temp_17_adj_2403\
        );

    \I__12991\ : LocalMux
    port map (
            O => \N__60297\,
            I => \Add_add_temp_17_adj_2403\
        );

    \I__12990\ : CascadeMux
    port map (
            O => \N__60292\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15200_cascade_\
        );

    \I__12989\ : InMux
    port map (
            O => \N__60289\,
            I => \N__60286\
        );

    \I__12988\ : LocalMux
    port map (
            O => \N__60286\,
            I => \N__60282\
        );

    \I__12987\ : InMux
    port map (
            O => \N__60285\,
            I => \N__60279\
        );

    \I__12986\ : Span4Mux_v
    port map (
            O => \N__60282\,
            I => \N__60274\
        );

    \I__12985\ : LocalMux
    port map (
            O => \N__60279\,
            I => \N__60274\
        );

    \I__12984\ : Span4Mux_v
    port map (
            O => \N__60274\,
            I => \N__60271\
        );

    \I__12983\ : Sp12to4
    port map (
            O => \N__60271\,
            I => \N__60267\
        );

    \I__12982\ : InMux
    port map (
            O => \N__60270\,
            I => \N__60264\
        );

    \I__12981\ : Odrv12
    port map (
            O => \N__60267\,
            I => \Add_add_temp_15_adj_2405\
        );

    \I__12980\ : LocalMux
    port map (
            O => \N__60264\,
            I => \Add_add_temp_15_adj_2405\
        );

    \I__12979\ : InMux
    port map (
            O => \N__60259\,
            I => \N__60255\
        );

    \I__12978\ : InMux
    port map (
            O => \N__60258\,
            I => \N__60252\
        );

    \I__12977\ : LocalMux
    port map (
            O => \N__60255\,
            I => \N__60248\
        );

    \I__12976\ : LocalMux
    port map (
            O => \N__60252\,
            I => \N__60245\
        );

    \I__12975\ : InMux
    port map (
            O => \N__60251\,
            I => \N__60242\
        );

    \I__12974\ : Span4Mux_h
    port map (
            O => \N__60248\,
            I => \N__60239\
        );

    \I__12973\ : Span4Mux_h
    port map (
            O => \N__60245\,
            I => \N__60234\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__60242\,
            I => \N__60234\
        );

    \I__12971\ : Odrv4
    port map (
            O => \N__60239\,
            I => \Add_add_temp_20_adj_2400\
        );

    \I__12970\ : Odrv4
    port map (
            O => \N__60234\,
            I => \Add_add_temp_20_adj_2400\
        );

    \I__12969\ : InMux
    port map (
            O => \N__60229\,
            I => \N__60226\
        );

    \I__12968\ : LocalMux
    port map (
            O => \N__60226\,
            I => \N__60223\
        );

    \I__12967\ : Span4Mux_h
    port map (
            O => \N__60223\,
            I => \N__60219\
        );

    \I__12966\ : InMux
    port map (
            O => \N__60222\,
            I => \N__60216\
        );

    \I__12965\ : Span4Mux_v
    port map (
            O => \N__60219\,
            I => \N__60212\
        );

    \I__12964\ : LocalMux
    port map (
            O => \N__60216\,
            I => \N__60209\
        );

    \I__12963\ : InMux
    port map (
            O => \N__60215\,
            I => \N__60206\
        );

    \I__12962\ : Odrv4
    port map (
            O => \N__60212\,
            I => \Add_add_temp_19_adj_2401\
        );

    \I__12961\ : Odrv4
    port map (
            O => \N__60209\,
            I => \Add_add_temp_19_adj_2401\
        );

    \I__12960\ : LocalMux
    port map (
            O => \N__60206\,
            I => \Add_add_temp_19_adj_2401\
        );

    \I__12959\ : CascadeMux
    port map (
            O => \N__60199\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20680_cascade_\
        );

    \I__12958\ : InMux
    port map (
            O => \N__60196\,
            I => \N__60193\
        );

    \I__12957\ : LocalMux
    port map (
            O => \N__60193\,
            I => \N__60190\
        );

    \I__12956\ : Span4Mux_h
    port map (
            O => \N__60190\,
            I => \N__60186\
        );

    \I__12955\ : InMux
    port map (
            O => \N__60189\,
            I => \N__60183\
        );

    \I__12954\ : Span4Mux_v
    port map (
            O => \N__60186\,
            I => \N__60178\
        );

    \I__12953\ : LocalMux
    port map (
            O => \N__60183\,
            I => \N__60178\
        );

    \I__12952\ : Span4Mux_v
    port map (
            O => \N__60178\,
            I => \N__60175\
        );

    \I__12951\ : Span4Mux_h
    port map (
            O => \N__60175\,
            I => \N__60171\
        );

    \I__12950\ : InMux
    port map (
            O => \N__60174\,
            I => \N__60168\
        );

    \I__12949\ : Odrv4
    port map (
            O => \N__60171\,
            I => \Add_add_temp_18_adj_2402\
        );

    \I__12948\ : LocalMux
    port map (
            O => \N__60168\,
            I => \Add_add_temp_18_adj_2402\
        );

    \I__12947\ : InMux
    port map (
            O => \N__60163\,
            I => \N__60160\
        );

    \I__12946\ : LocalMux
    port map (
            O => \N__60160\,
            I => \N__60157\
        );

    \I__12945\ : Span4Mux_h
    port map (
            O => \N__60157\,
            I => \N__60154\
        );

    \I__12944\ : Odrv4
    port map (
            O => \N__60154\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19733\
        );

    \I__12943\ : InMux
    port map (
            O => \N__60151\,
            I => \N__60148\
        );

    \I__12942\ : LocalMux
    port map (
            O => \N__60148\,
            I => \N__60144\
        );

    \I__12941\ : CascadeMux
    port map (
            O => \N__60147\,
            I => \N__60141\
        );

    \I__12940\ : Span4Mux_h
    port map (
            O => \N__60144\,
            I => \N__60137\
        );

    \I__12939\ : InMux
    port map (
            O => \N__60141\,
            I => \N__60132\
        );

    \I__12938\ : InMux
    port map (
            O => \N__60140\,
            I => \N__60132\
        );

    \I__12937\ : Odrv4
    port map (
            O => \N__60137\,
            I => \Add_add_temp_5_adj_2415\
        );

    \I__12936\ : LocalMux
    port map (
            O => \N__60132\,
            I => \Add_add_temp_5_adj_2415\
        );

    \I__12935\ : InMux
    port map (
            O => \N__60127\,
            I => \N__60124\
        );

    \I__12934\ : LocalMux
    port map (
            O => \N__60124\,
            I => \N__60120\
        );

    \I__12933\ : InMux
    port map (
            O => \N__60123\,
            I => \N__60117\
        );

    \I__12932\ : Odrv4
    port map (
            O => \N__60120\,
            I => \Add_add_temp_4_adj_2416\
        );

    \I__12931\ : LocalMux
    port map (
            O => \N__60117\,
            I => \Add_add_temp_4_adj_2416\
        );

    \I__12930\ : InMux
    port map (
            O => \N__60112\,
            I => \N__60107\
        );

    \I__12929\ : InMux
    port map (
            O => \N__60111\,
            I => \N__60102\
        );

    \I__12928\ : InMux
    port map (
            O => \N__60110\,
            I => \N__60102\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__60107\,
            I => \Add_add_temp_8_adj_2412\
        );

    \I__12926\ : LocalMux
    port map (
            O => \N__60102\,
            I => \Add_add_temp_8_adj_2412\
        );

    \I__12925\ : InMux
    port map (
            O => \N__60097\,
            I => \N__60094\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__60094\,
            I => \N__60089\
        );

    \I__12923\ : InMux
    port map (
            O => \N__60093\,
            I => \N__60084\
        );

    \I__12922\ : InMux
    port map (
            O => \N__60092\,
            I => \N__60084\
        );

    \I__12921\ : Odrv12
    port map (
            O => \N__60089\,
            I => \Add_add_temp_7_adj_2413\
        );

    \I__12920\ : LocalMux
    port map (
            O => \N__60084\,
            I => \Add_add_temp_7_adj_2413\
        );

    \I__12919\ : CascadeMux
    port map (
            O => \N__60079\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20722_cascade_\
        );

    \I__12918\ : InMux
    port map (
            O => \N__60076\,
            I => \N__60073\
        );

    \I__12917\ : LocalMux
    port map (
            O => \N__60073\,
            I => \N__60070\
        );

    \I__12916\ : Span4Mux_v
    port map (
            O => \N__60070\,
            I => \N__60065\
        );

    \I__12915\ : InMux
    port map (
            O => \N__60069\,
            I => \N__60060\
        );

    \I__12914\ : InMux
    port map (
            O => \N__60068\,
            I => \N__60060\
        );

    \I__12913\ : Odrv4
    port map (
            O => \N__60065\,
            I => \Add_add_temp_6_adj_2414\
        );

    \I__12912\ : LocalMux
    port map (
            O => \N__60060\,
            I => \Add_add_temp_6_adj_2414\
        );

    \I__12911\ : InMux
    port map (
            O => \N__60055\,
            I => \N__60052\
        );

    \I__12910\ : LocalMux
    port map (
            O => \N__60052\,
            I => \N__60049\
        );

    \I__12909\ : Span4Mux_h
    port map (
            O => \N__60049\,
            I => \N__60046\
        );

    \I__12908\ : Odrv4
    port map (
            O => \N__60046\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_26\
        );

    \I__12907\ : InMux
    port map (
            O => \N__60043\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15994\
        );

    \I__12906\ : CascadeMux
    port map (
            O => \N__60040\,
            I => \N__60037\
        );

    \I__12905\ : InMux
    port map (
            O => \N__60037\,
            I => \N__60034\
        );

    \I__12904\ : LocalMux
    port map (
            O => \N__60034\,
            I => \N__60031\
        );

    \I__12903\ : Span4Mux_h
    port map (
            O => \N__60031\,
            I => \N__60028\
        );

    \I__12902\ : Odrv4
    port map (
            O => \N__60028\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_27\
        );

    \I__12901\ : InMux
    port map (
            O => \N__60025\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15995\
        );

    \I__12900\ : CascadeMux
    port map (
            O => \N__60022\,
            I => \N__60019\
        );

    \I__12899\ : InMux
    port map (
            O => \N__60019\,
            I => \N__60016\
        );

    \I__12898\ : LocalMux
    port map (
            O => \N__60016\,
            I => \N__60013\
        );

    \I__12897\ : Span4Mux_v
    port map (
            O => \N__60013\,
            I => \N__60010\
        );

    \I__12896\ : Odrv4
    port map (
            O => \N__60010\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_28\
        );

    \I__12895\ : InMux
    port map (
            O => \N__60007\,
            I => \N__59998\
        );

    \I__12894\ : InMux
    port map (
            O => \N__60006\,
            I => \N__59998\
        );

    \I__12893\ : InMux
    port map (
            O => \N__60005\,
            I => \N__59998\
        );

    \I__12892\ : LocalMux
    port map (
            O => \N__59998\,
            I => \N__59995\
        );

    \I__12891\ : Odrv12
    port map (
            O => \N__59995\,
            I => \Add_add_temp_28\
        );

    \I__12890\ : InMux
    port map (
            O => \N__59992\,
            I => \bfn_22_22_0_\
        );

    \I__12889\ : CascadeMux
    port map (
            O => \N__59989\,
            I => \N__59986\
        );

    \I__12888\ : InMux
    port map (
            O => \N__59986\,
            I => \N__59983\
        );

    \I__12887\ : LocalMux
    port map (
            O => \N__59983\,
            I => \N__59980\
        );

    \I__12886\ : Span4Mux_v
    port map (
            O => \N__59980\,
            I => \N__59977\
        );

    \I__12885\ : Odrv4
    port map (
            O => \N__59977\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_29\
        );

    \I__12884\ : InMux
    port map (
            O => \N__59974\,
            I => \N__59965\
        );

    \I__12883\ : InMux
    port map (
            O => \N__59973\,
            I => \N__59965\
        );

    \I__12882\ : InMux
    port map (
            O => \N__59972\,
            I => \N__59965\
        );

    \I__12881\ : LocalMux
    port map (
            O => \N__59965\,
            I => \N__59962\
        );

    \I__12880\ : Span4Mux_v
    port map (
            O => \N__59962\,
            I => \N__59959\
        );

    \I__12879\ : Odrv4
    port map (
            O => \N__59959\,
            I => \Add_add_temp_29\
        );

    \I__12878\ : InMux
    port map (
            O => \N__59956\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15997\
        );

    \I__12877\ : CascadeMux
    port map (
            O => \N__59953\,
            I => \N__59950\
        );

    \I__12876\ : InMux
    port map (
            O => \N__59950\,
            I => \N__59947\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__59947\,
            I => \N__59944\
        );

    \I__12874\ : Span4Mux_v
    port map (
            O => \N__59944\,
            I => \N__59941\
        );

    \I__12873\ : Span4Mux_h
    port map (
            O => \N__59941\,
            I => \N__59938\
        );

    \I__12872\ : Odrv4
    port map (
            O => \N__59938\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_30\
        );

    \I__12871\ : InMux
    port map (
            O => \N__59935\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15998\
        );

    \I__12870\ : InMux
    port map (
            O => \N__59932\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15999\
        );

    \I__12869\ : InMux
    port map (
            O => \N__59929\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n16000\
        );

    \I__12868\ : InMux
    port map (
            O => \N__59926\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n16001\
        );

    \I__12867\ : CascadeMux
    port map (
            O => \N__59923\,
            I => \N__59920\
        );

    \I__12866\ : InMux
    port map (
            O => \N__59920\,
            I => \N__59917\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__59917\,
            I => \N__59914\
        );

    \I__12864\ : Span4Mux_h
    port map (
            O => \N__59914\,
            I => \N__59911\
        );

    \I__12863\ : Odrv4
    port map (
            O => \N__59911\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_17\
        );

    \I__12862\ : InMux
    port map (
            O => \N__59908\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15985\
        );

    \I__12861\ : CascadeMux
    port map (
            O => \N__59905\,
            I => \N__59902\
        );

    \I__12860\ : InMux
    port map (
            O => \N__59902\,
            I => \N__59899\
        );

    \I__12859\ : LocalMux
    port map (
            O => \N__59899\,
            I => \N__59896\
        );

    \I__12858\ : Span4Mux_h
    port map (
            O => \N__59896\,
            I => \N__59893\
        );

    \I__12857\ : Odrv4
    port map (
            O => \N__59893\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_18\
        );

    \I__12856\ : InMux
    port map (
            O => \N__59890\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15986\
        );

    \I__12855\ : InMux
    port map (
            O => \N__59887\,
            I => \N__59884\
        );

    \I__12854\ : LocalMux
    port map (
            O => \N__59884\,
            I => \N__59881\
        );

    \I__12853\ : Span4Mux_h
    port map (
            O => \N__59881\,
            I => \N__59878\
        );

    \I__12852\ : Odrv4
    port map (
            O => \N__59878\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_19\
        );

    \I__12851\ : InMux
    port map (
            O => \N__59875\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15987\
        );

    \I__12850\ : CascadeMux
    port map (
            O => \N__59872\,
            I => \N__59869\
        );

    \I__12849\ : InMux
    port map (
            O => \N__59869\,
            I => \N__59866\
        );

    \I__12848\ : LocalMux
    port map (
            O => \N__59866\,
            I => \N__59863\
        );

    \I__12847\ : Span4Mux_v
    port map (
            O => \N__59863\,
            I => \N__59860\
        );

    \I__12846\ : Odrv4
    port map (
            O => \N__59860\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_20\
        );

    \I__12845\ : InMux
    port map (
            O => \N__59857\,
            I => \bfn_22_21_0_\
        );

    \I__12844\ : CascadeMux
    port map (
            O => \N__59854\,
            I => \N__59851\
        );

    \I__12843\ : InMux
    port map (
            O => \N__59851\,
            I => \N__59848\
        );

    \I__12842\ : LocalMux
    port map (
            O => \N__59848\,
            I => \N__59845\
        );

    \I__12841\ : Span4Mux_v
    port map (
            O => \N__59845\,
            I => \N__59842\
        );

    \I__12840\ : Odrv4
    port map (
            O => \N__59842\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_21\
        );

    \I__12839\ : InMux
    port map (
            O => \N__59839\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15989\
        );

    \I__12838\ : CascadeMux
    port map (
            O => \N__59836\,
            I => \N__59833\
        );

    \I__12837\ : InMux
    port map (
            O => \N__59833\,
            I => \N__59830\
        );

    \I__12836\ : LocalMux
    port map (
            O => \N__59830\,
            I => \N__59827\
        );

    \I__12835\ : Span4Mux_v
    port map (
            O => \N__59827\,
            I => \N__59824\
        );

    \I__12834\ : Odrv4
    port map (
            O => \N__59824\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_22\
        );

    \I__12833\ : InMux
    port map (
            O => \N__59821\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15990\
        );

    \I__12832\ : InMux
    port map (
            O => \N__59818\,
            I => \N__59815\
        );

    \I__12831\ : LocalMux
    port map (
            O => \N__59815\,
            I => \N__59812\
        );

    \I__12830\ : Span4Mux_v
    port map (
            O => \N__59812\,
            I => \N__59809\
        );

    \I__12829\ : Odrv4
    port map (
            O => \N__59809\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_23\
        );

    \I__12828\ : InMux
    port map (
            O => \N__59806\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15991\
        );

    \I__12827\ : InMux
    port map (
            O => \N__59803\,
            I => \N__59800\
        );

    \I__12826\ : LocalMux
    port map (
            O => \N__59800\,
            I => \N__59797\
        );

    \I__12825\ : Span4Mux_v
    port map (
            O => \N__59797\,
            I => \N__59794\
        );

    \I__12824\ : Odrv4
    port map (
            O => \N__59794\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_24\
        );

    \I__12823\ : InMux
    port map (
            O => \N__59791\,
            I => \N__59788\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__59788\,
            I => \N__59783\
        );

    \I__12821\ : InMux
    port map (
            O => \N__59787\,
            I => \N__59778\
        );

    \I__12820\ : InMux
    port map (
            O => \N__59786\,
            I => \N__59778\
        );

    \I__12819\ : Span4Mux_h
    port map (
            O => \N__59783\,
            I => \N__59773\
        );

    \I__12818\ : LocalMux
    port map (
            O => \N__59778\,
            I => \N__59773\
        );

    \I__12817\ : Odrv4
    port map (
            O => \N__59773\,
            I => \Add_add_temp_24\
        );

    \I__12816\ : InMux
    port map (
            O => \N__59770\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15992\
        );

    \I__12815\ : CascadeMux
    port map (
            O => \N__59767\,
            I => \N__59764\
        );

    \I__12814\ : InMux
    port map (
            O => \N__59764\,
            I => \N__59761\
        );

    \I__12813\ : LocalMux
    port map (
            O => \N__59761\,
            I => \N__59758\
        );

    \I__12812\ : Span4Mux_h
    port map (
            O => \N__59758\,
            I => \N__59755\
        );

    \I__12811\ : Odrv4
    port map (
            O => \N__59755\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_25\
        );

    \I__12810\ : InMux
    port map (
            O => \N__59752\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15993\
        );

    \I__12809\ : CascadeMux
    port map (
            O => \N__59749\,
            I => \N__59746\
        );

    \I__12808\ : InMux
    port map (
            O => \N__59746\,
            I => \N__59743\
        );

    \I__12807\ : LocalMux
    port map (
            O => \N__59743\,
            I => \N__59740\
        );

    \I__12806\ : Odrv4
    port map (
            O => \N__59740\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_9\
        );

    \I__12805\ : InMux
    port map (
            O => \N__59737\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15977\
        );

    \I__12804\ : InMux
    port map (
            O => \N__59734\,
            I => \N__59731\
        );

    \I__12803\ : LocalMux
    port map (
            O => \N__59731\,
            I => \N__59728\
        );

    \I__12802\ : Odrv12
    port map (
            O => \N__59728\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_6\
        );

    \I__12801\ : CascadeMux
    port map (
            O => \N__59725\,
            I => \N__59722\
        );

    \I__12800\ : InMux
    port map (
            O => \N__59722\,
            I => \N__59719\
        );

    \I__12799\ : LocalMux
    port map (
            O => \N__59719\,
            I => \N__59716\
        );

    \I__12798\ : Span4Mux_h
    port map (
            O => \N__59716\,
            I => \N__59713\
        );

    \I__12797\ : Odrv4
    port map (
            O => \N__59713\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_10\
        );

    \I__12796\ : InMux
    port map (
            O => \N__59710\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15978\
        );

    \I__12795\ : InMux
    port map (
            O => \N__59707\,
            I => \N__59704\
        );

    \I__12794\ : LocalMux
    port map (
            O => \N__59704\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_11\
        );

    \I__12793\ : InMux
    port map (
            O => \N__59701\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15979\
        );

    \I__12792\ : CascadeMux
    port map (
            O => \N__59698\,
            I => \N__59695\
        );

    \I__12791\ : InMux
    port map (
            O => \N__59695\,
            I => \N__59692\
        );

    \I__12790\ : LocalMux
    port map (
            O => \N__59692\,
            I => \N__59689\
        );

    \I__12789\ : Odrv4
    port map (
            O => \N__59689\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_12\
        );

    \I__12788\ : InMux
    port map (
            O => \N__59686\,
            I => \bfn_22_20_0_\
        );

    \I__12787\ : CascadeMux
    port map (
            O => \N__59683\,
            I => \N__59680\
        );

    \I__12786\ : InMux
    port map (
            O => \N__59680\,
            I => \N__59677\
        );

    \I__12785\ : LocalMux
    port map (
            O => \N__59677\,
            I => \N__59674\
        );

    \I__12784\ : Odrv4
    port map (
            O => \N__59674\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_13\
        );

    \I__12783\ : InMux
    port map (
            O => \N__59671\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15981\
        );

    \I__12782\ : CascadeMux
    port map (
            O => \N__59668\,
            I => \N__59665\
        );

    \I__12781\ : InMux
    port map (
            O => \N__59665\,
            I => \N__59662\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__59662\,
            I => \N__59659\
        );

    \I__12779\ : Odrv4
    port map (
            O => \N__59659\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_14\
        );

    \I__12778\ : InMux
    port map (
            O => \N__59656\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15982\
        );

    \I__12777\ : InMux
    port map (
            O => \N__59653\,
            I => \N__59650\
        );

    \I__12776\ : LocalMux
    port map (
            O => \N__59650\,
            I => \N__59647\
        );

    \I__12775\ : Odrv4
    port map (
            O => \N__59647\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_15\
        );

    \I__12774\ : InMux
    port map (
            O => \N__59644\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15983\
        );

    \I__12773\ : CascadeMux
    port map (
            O => \N__59641\,
            I => \N__59638\
        );

    \I__12772\ : InMux
    port map (
            O => \N__59638\,
            I => \N__59635\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__59635\,
            I => \N__59632\
        );

    \I__12770\ : Span4Mux_v
    port map (
            O => \N__59632\,
            I => \N__59629\
        );

    \I__12769\ : Span4Mux_h
    port map (
            O => \N__59629\,
            I => \N__59626\
        );

    \I__12768\ : Odrv4
    port map (
            O => \N__59626\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_16\
        );

    \I__12767\ : InMux
    port map (
            O => \N__59623\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15984\
        );

    \I__12766\ : CascadeMux
    port map (
            O => \N__59620\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20658_cascade_\
        );

    \I__12765\ : CascadeMux
    port map (
            O => \N__59617\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20648_cascade_\
        );

    \I__12764\ : InMux
    port map (
            O => \N__59614\,
            I => \N__59611\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__59611\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20634\
        );

    \I__12762\ : InMux
    port map (
            O => \N__59608\,
            I => \N__59605\
        );

    \I__12761\ : LocalMux
    port map (
            O => \N__59605\,
            I => \N__59602\
        );

    \I__12760\ : Odrv4
    port map (
            O => \N__59602\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_0\
        );

    \I__12759\ : CascadeMux
    port map (
            O => \N__59599\,
            I => \N__59596\
        );

    \I__12758\ : InMux
    port map (
            O => \N__59596\,
            I => \N__59593\
        );

    \I__12757\ : LocalMux
    port map (
            O => \N__59593\,
            I => \N__59590\
        );

    \I__12756\ : Odrv4
    port map (
            O => \N__59590\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_4\
        );

    \I__12755\ : InMux
    port map (
            O => \N__59587\,
            I => \N__59584\
        );

    \I__12754\ : LocalMux
    port map (
            O => \N__59584\,
            I => \N__59581\
        );

    \I__12753\ : Odrv4
    port map (
            O => \N__59581\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_1\
        );

    \I__12752\ : CascadeMux
    port map (
            O => \N__59578\,
            I => \N__59575\
        );

    \I__12751\ : InMux
    port map (
            O => \N__59575\,
            I => \N__59572\
        );

    \I__12750\ : LocalMux
    port map (
            O => \N__59572\,
            I => \N__59569\
        );

    \I__12749\ : Span4Mux_v
    port map (
            O => \N__59569\,
            I => \N__59566\
        );

    \I__12748\ : Odrv4
    port map (
            O => \N__59566\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_5\
        );

    \I__12747\ : InMux
    port map (
            O => \N__59563\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15973\
        );

    \I__12746\ : InMux
    port map (
            O => \N__59560\,
            I => \N__59557\
        );

    \I__12745\ : LocalMux
    port map (
            O => \N__59557\,
            I => \N__59554\
        );

    \I__12744\ : Odrv4
    port map (
            O => \N__59554\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_2\
        );

    \I__12743\ : CascadeMux
    port map (
            O => \N__59551\,
            I => \N__59548\
        );

    \I__12742\ : InMux
    port map (
            O => \N__59548\,
            I => \N__59545\
        );

    \I__12741\ : LocalMux
    port map (
            O => \N__59545\,
            I => \N__59542\
        );

    \I__12740\ : Odrv4
    port map (
            O => \N__59542\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_6\
        );

    \I__12739\ : InMux
    port map (
            O => \N__59539\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15974\
        );

    \I__12738\ : InMux
    port map (
            O => \N__59536\,
            I => \N__59533\
        );

    \I__12737\ : LocalMux
    port map (
            O => \N__59533\,
            I => \N__59530\
        );

    \I__12736\ : Odrv4
    port map (
            O => \N__59530\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_3\
        );

    \I__12735\ : CascadeMux
    port map (
            O => \N__59527\,
            I => \N__59524\
        );

    \I__12734\ : InMux
    port map (
            O => \N__59524\,
            I => \N__59521\
        );

    \I__12733\ : LocalMux
    port map (
            O => \N__59521\,
            I => \N__59518\
        );

    \I__12732\ : Span4Mux_v
    port map (
            O => \N__59518\,
            I => \N__59515\
        );

    \I__12731\ : Odrv4
    port map (
            O => \N__59515\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_7\
        );

    \I__12730\ : InMux
    port map (
            O => \N__59512\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15975\
        );

    \I__12729\ : CascadeMux
    port map (
            O => \N__59509\,
            I => \N__59506\
        );

    \I__12728\ : InMux
    port map (
            O => \N__59506\,
            I => \N__59503\
        );

    \I__12727\ : LocalMux
    port map (
            O => \N__59503\,
            I => \N__59500\
        );

    \I__12726\ : Span4Mux_v
    port map (
            O => \N__59500\,
            I => \N__59497\
        );

    \I__12725\ : Odrv4
    port map (
            O => \N__59497\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_8\
        );

    \I__12724\ : InMux
    port map (
            O => \N__59494\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15976\
        );

    \I__12723\ : CascadeMux
    port map (
            O => \N__59491\,
            I => \Saturate_out1_31__N_267_cascade_\
        );

    \I__12722\ : CascadeMux
    port map (
            O => \N__59488\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19842_cascade_\
        );

    \I__12721\ : CascadeMux
    port map (
            O => \N__59485\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20666_cascade_\
        );

    \I__12720\ : InMux
    port map (
            O => \N__59482\,
            I => \N__59476\
        );

    \I__12719\ : InMux
    port map (
            O => \N__59481\,
            I => \N__59476\
        );

    \I__12718\ : LocalMux
    port map (
            O => \N__59476\,
            I => \N__59473\
        );

    \I__12717\ : Span4Mux_h
    port map (
            O => \N__59473\,
            I => \N__59470\
        );

    \I__12716\ : Span4Mux_v
    port map (
            O => \N__59470\,
            I => \N__59467\
        );

    \I__12715\ : Span4Mux_v
    port map (
            O => \N__59467\,
            I => \N__59462\
        );

    \I__12714\ : InMux
    port map (
            O => \N__59466\,
            I => \N__59459\
        );

    \I__12713\ : InMux
    port map (
            O => \N__59465\,
            I => \N__59456\
        );

    \I__12712\ : Odrv4
    port map (
            O => \N__59462\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__59459\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15\
        );

    \I__12710\ : LocalMux
    port map (
            O => \N__59456\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15\
        );

    \I__12709\ : InMux
    port map (
            O => \N__59449\,
            I => \N__59446\
        );

    \I__12708\ : LocalMux
    port map (
            O => \N__59446\,
            I => \foc.qVoltage_6\
        );

    \I__12707\ : InMux
    port map (
            O => \N__59443\,
            I => \N__59437\
        );

    \I__12706\ : InMux
    port map (
            O => \N__59442\,
            I => \N__59434\
        );

    \I__12705\ : CascadeMux
    port map (
            O => \N__59441\,
            I => \N__59430\
        );

    \I__12704\ : CascadeMux
    port map (
            O => \N__59440\,
            I => \N__59420\
        );

    \I__12703\ : LocalMux
    port map (
            O => \N__59437\,
            I => \N__59412\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__59434\,
            I => \N__59409\
        );

    \I__12701\ : InMux
    port map (
            O => \N__59433\,
            I => \N__59402\
        );

    \I__12700\ : InMux
    port map (
            O => \N__59430\,
            I => \N__59402\
        );

    \I__12699\ : InMux
    port map (
            O => \N__59429\,
            I => \N__59402\
        );

    \I__12698\ : InMux
    port map (
            O => \N__59428\,
            I => \N__59391\
        );

    \I__12697\ : InMux
    port map (
            O => \N__59427\,
            I => \N__59391\
        );

    \I__12696\ : InMux
    port map (
            O => \N__59426\,
            I => \N__59391\
        );

    \I__12695\ : InMux
    port map (
            O => \N__59425\,
            I => \N__59391\
        );

    \I__12694\ : InMux
    port map (
            O => \N__59424\,
            I => \N__59391\
        );

    \I__12693\ : InMux
    port map (
            O => \N__59423\,
            I => \N__59388\
        );

    \I__12692\ : InMux
    port map (
            O => \N__59420\,
            I => \N__59381\
        );

    \I__12691\ : InMux
    port map (
            O => \N__59419\,
            I => \N__59381\
        );

    \I__12690\ : InMux
    port map (
            O => \N__59418\,
            I => \N__59381\
        );

    \I__12689\ : InMux
    port map (
            O => \N__59417\,
            I => \N__59374\
        );

    \I__12688\ : InMux
    port map (
            O => \N__59416\,
            I => \N__59374\
        );

    \I__12687\ : InMux
    port map (
            O => \N__59415\,
            I => \N__59374\
        );

    \I__12686\ : Odrv4
    port map (
            O => \N__59412\,
            I => \foc.Out_31__N_332\
        );

    \I__12685\ : Odrv4
    port map (
            O => \N__59409\,
            I => \foc.Out_31__N_332\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__59402\,
            I => \foc.Out_31__N_332\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__59391\,
            I => \foc.Out_31__N_332\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__59388\,
            I => \foc.Out_31__N_332\
        );

    \I__12681\ : LocalMux
    port map (
            O => \N__59381\,
            I => \foc.Out_31__N_332\
        );

    \I__12680\ : LocalMux
    port map (
            O => \N__59374\,
            I => \foc.Out_31__N_332\
        );

    \I__12679\ : InMux
    port map (
            O => \N__59359\,
            I => \N__59355\
        );

    \I__12678\ : InMux
    port map (
            O => \N__59358\,
            I => \N__59352\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__59355\,
            I => \N__59345\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__59352\,
            I => \N__59345\
        );

    \I__12675\ : InMux
    port map (
            O => \N__59351\,
            I => \N__59342\
        );

    \I__12674\ : InMux
    port map (
            O => \N__59350\,
            I => \N__59339\
        );

    \I__12673\ : Span12Mux_v
    port map (
            O => \N__59345\,
            I => \N__59336\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__59342\,
            I => \N__59331\
        );

    \I__12671\ : LocalMux
    port map (
            O => \N__59339\,
            I => \N__59331\
        );

    \I__12670\ : Odrv12
    port map (
            O => \N__59336\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21\
        );

    \I__12669\ : Odrv12
    port map (
            O => \N__59331\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21\
        );

    \I__12668\ : CascadeMux
    port map (
            O => \N__59326\,
            I => \N__59322\
        );

    \I__12667\ : InMux
    port map (
            O => \N__59325\,
            I => \N__59319\
        );

    \I__12666\ : InMux
    port map (
            O => \N__59322\,
            I => \N__59316\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__59319\,
            I => \N__59312\
        );

    \I__12664\ : LocalMux
    port map (
            O => \N__59316\,
            I => \N__59309\
        );

    \I__12663\ : CascadeMux
    port map (
            O => \N__59315\,
            I => \N__59301\
        );

    \I__12662\ : Span12Mux_s11_h
    port map (
            O => \N__59312\,
            I => \N__59287\
        );

    \I__12661\ : Sp12to4
    port map (
            O => \N__59309\,
            I => \N__59287\
        );

    \I__12660\ : InMux
    port map (
            O => \N__59308\,
            I => \N__59280\
        );

    \I__12659\ : InMux
    port map (
            O => \N__59307\,
            I => \N__59280\
        );

    \I__12658\ : InMux
    port map (
            O => \N__59306\,
            I => \N__59280\
        );

    \I__12657\ : InMux
    port map (
            O => \N__59305\,
            I => \N__59269\
        );

    \I__12656\ : InMux
    port map (
            O => \N__59304\,
            I => \N__59269\
        );

    \I__12655\ : InMux
    port map (
            O => \N__59301\,
            I => \N__59269\
        );

    \I__12654\ : InMux
    port map (
            O => \N__59300\,
            I => \N__59269\
        );

    \I__12653\ : InMux
    port map (
            O => \N__59299\,
            I => \N__59269\
        );

    \I__12652\ : InMux
    port map (
            O => \N__59298\,
            I => \N__59266\
        );

    \I__12651\ : InMux
    port map (
            O => \N__59297\,
            I => \N__59259\
        );

    \I__12650\ : InMux
    port map (
            O => \N__59296\,
            I => \N__59259\
        );

    \I__12649\ : InMux
    port map (
            O => \N__59295\,
            I => \N__59259\
        );

    \I__12648\ : InMux
    port map (
            O => \N__59294\,
            I => \N__59252\
        );

    \I__12647\ : InMux
    port map (
            O => \N__59293\,
            I => \N__59252\
        );

    \I__12646\ : InMux
    port map (
            O => \N__59292\,
            I => \N__59252\
        );

    \I__12645\ : Odrv12
    port map (
            O => \N__59287\,
            I => \foc.Out_31__N_333\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__59280\,
            I => \foc.Out_31__N_333\
        );

    \I__12643\ : LocalMux
    port map (
            O => \N__59269\,
            I => \foc.Out_31__N_333\
        );

    \I__12642\ : LocalMux
    port map (
            O => \N__59266\,
            I => \foc.Out_31__N_333\
        );

    \I__12641\ : LocalMux
    port map (
            O => \N__59259\,
            I => \foc.Out_31__N_333\
        );

    \I__12640\ : LocalMux
    port map (
            O => \N__59252\,
            I => \foc.Out_31__N_333\
        );

    \I__12639\ : InMux
    port map (
            O => \N__59239\,
            I => \N__59236\
        );

    \I__12638\ : LocalMux
    port map (
            O => \N__59236\,
            I => \foc.qVoltage_12\
        );

    \I__12637\ : CascadeMux
    port map (
            O => \N__59233\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15264_cascade_\
        );

    \I__12636\ : CascadeMux
    port map (
            O => \N__59230\,
            I => \foc.Out_31__N_333_adj_2310_cascade_\
        );

    \I__12635\ : InMux
    port map (
            O => \N__59227\,
            I => \N__59224\
        );

    \I__12634\ : LocalMux
    port map (
            O => \N__59224\,
            I => \foc.dVoltage_14\
        );

    \I__12633\ : CascadeMux
    port map (
            O => \N__59221\,
            I => \foc.dVoltage_3_cascade_\
        );

    \I__12632\ : InMux
    port map (
            O => \N__59218\,
            I => \N__59215\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__59215\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20572\
        );

    \I__12630\ : CascadeMux
    port map (
            O => \N__59212\,
            I => \foc.dVoltage_11_cascade_\
        );

    \I__12629\ : InMux
    port map (
            O => \N__59209\,
            I => \N__59206\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__59206\,
            I => \foc.dVoltage_9\
        );

    \I__12627\ : InMux
    port map (
            O => \N__59203\,
            I => \N__59200\
        );

    \I__12626\ : LocalMux
    port map (
            O => \N__59200\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20566\
        );

    \I__12625\ : InMux
    port map (
            O => \N__59197\,
            I => \N__59191\
        );

    \I__12624\ : InMux
    port map (
            O => \N__59196\,
            I => \N__59191\
        );

    \I__12623\ : LocalMux
    port map (
            O => \N__59191\,
            I => \N__59188\
        );

    \I__12622\ : Span4Mux_h
    port map (
            O => \N__59188\,
            I => \N__59185\
        );

    \I__12621\ : Span4Mux_v
    port map (
            O => \N__59185\,
            I => \N__59182\
        );

    \I__12620\ : Span4Mux_v
    port map (
            O => \N__59182\,
            I => \N__59177\
        );

    \I__12619\ : InMux
    port map (
            O => \N__59181\,
            I => \N__59174\
        );

    \I__12618\ : InMux
    port map (
            O => \N__59180\,
            I => \N__59171\
        );

    \I__12617\ : Odrv4
    port map (
            O => \N__59177\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__59174\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11\
        );

    \I__12615\ : LocalMux
    port map (
            O => \N__59171\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11\
        );

    \I__12614\ : CascadeMux
    port map (
            O => \N__59164\,
            I => \foc.qVoltage_2_cascade_\
        );

    \I__12613\ : InMux
    port map (
            O => \N__59161\,
            I => \N__59158\
        );

    \I__12612\ : LocalMux
    port map (
            O => \N__59158\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20594\
        );

    \I__12611\ : InMux
    port map (
            O => \N__59155\,
            I => \N__59152\
        );

    \I__12610\ : LocalMux
    port map (
            O => \N__59152\,
            I => \N__59147\
        );

    \I__12609\ : InMux
    port map (
            O => \N__59151\,
            I => \N__59144\
        );

    \I__12608\ : InMux
    port map (
            O => \N__59150\,
            I => \N__59141\
        );

    \I__12607\ : Span12Mux_h
    port map (
            O => \N__59147\,
            I => \N__59134\
        );

    \I__12606\ : LocalMux
    port map (
            O => \N__59144\,
            I => \N__59134\
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__59141\,
            I => \N__59134\
        );

    \I__12604\ : Odrv12
    port map (
            O => \N__59134\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_20\
        );

    \I__12603\ : CascadeMux
    port map (
            O => \N__59131\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_cascade_\
        );

    \I__12602\ : InMux
    port map (
            O => \N__59128\,
            I => \N__59125\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__59125\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20612\
        );

    \I__12600\ : InMux
    port map (
            O => \N__59122\,
            I => \N__59119\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__59119\,
            I => \N__59116\
        );

    \I__12598\ : Span4Mux_h
    port map (
            O => \N__59116\,
            I => \N__59113\
        );

    \I__12597\ : Span4Mux_v
    port map (
            O => \N__59113\,
            I => \N__59110\
        );

    \I__12596\ : Odrv4
    port map (
            O => \N__59110\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20618\
        );

    \I__12595\ : CascadeMux
    port map (
            O => \N__59107\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20550_cascade_\
        );

    \I__12594\ : InMux
    port map (
            O => \N__59104\,
            I => \N__59101\
        );

    \I__12593\ : LocalMux
    port map (
            O => \N__59101\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20556\
        );

    \I__12592\ : CascadeMux
    port map (
            O => \N__59098\,
            I => \foc.dVoltage_5_cascade_\
        );

    \I__12591\ : InMux
    port map (
            O => \N__59095\,
            I => \N__59092\
        );

    \I__12590\ : LocalMux
    port map (
            O => \N__59092\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20554\
        );

    \I__12589\ : CascadeMux
    port map (
            O => \N__59089\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15_cascade_\
        );

    \I__12588\ : InMux
    port map (
            O => \N__59086\,
            I => \N__59083\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__59083\,
            I => \foc.dVoltage_12\
        );

    \I__12586\ : InMux
    port map (
            O => \N__59080\,
            I => \N__59077\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__59077\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20560\
        );

    \I__12584\ : CascadeMux
    port map (
            O => \N__59074\,
            I => \foc.Out_31__N_332_adj_2312_cascade_\
        );

    \I__12583\ : InMux
    port map (
            O => \N__59071\,
            I => \N__59068\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__59068\,
            I => \foc.dVoltage_8\
        );

    \I__12581\ : InMux
    port map (
            O => \N__59065\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17542\
        );

    \I__12580\ : InMux
    port map (
            O => \N__59062\,
            I => \N__59059\
        );

    \I__12579\ : LocalMux
    port map (
            O => \N__59059\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n400\
        );

    \I__12578\ : InMux
    port map (
            O => \N__59056\,
            I => \bfn_22_12_0_\
        );

    \I__12577\ : CascadeMux
    port map (
            O => \N__59053\,
            I => \N__59050\
        );

    \I__12576\ : InMux
    port map (
            O => \N__59050\,
            I => \N__59047\
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__59047\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n449\
        );

    \I__12574\ : InMux
    port map (
            O => \N__59044\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17544\
        );

    \I__12573\ : InMux
    port map (
            O => \N__59041\,
            I => \N__59038\
        );

    \I__12572\ : LocalMux
    port map (
            O => \N__59038\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n498\
        );

    \I__12571\ : InMux
    port map (
            O => \N__59035\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17545\
        );

    \I__12570\ : CascadeMux
    port map (
            O => \N__59032\,
            I => \N__59029\
        );

    \I__12569\ : InMux
    port map (
            O => \N__59029\,
            I => \N__59026\
        );

    \I__12568\ : LocalMux
    port map (
            O => \N__59026\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n547\
        );

    \I__12567\ : InMux
    port map (
            O => \N__59023\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17546\
        );

    \I__12566\ : InMux
    port map (
            O => \N__59020\,
            I => \N__59017\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__59017\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n596\
        );

    \I__12564\ : InMux
    port map (
            O => \N__59014\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17547\
        );

    \I__12563\ : CascadeMux
    port map (
            O => \N__59011\,
            I => \N__59008\
        );

    \I__12562\ : InMux
    port map (
            O => \N__59008\,
            I => \N__59005\
        );

    \I__12561\ : LocalMux
    port map (
            O => \N__59005\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n645\
        );

    \I__12560\ : InMux
    port map (
            O => \N__59002\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17548\
        );

    \I__12559\ : InMux
    port map (
            O => \N__58999\,
            I => \N__58996\
        );

    \I__12558\ : LocalMux
    port map (
            O => \N__58996\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n694\
        );

    \I__12557\ : CascadeMux
    port map (
            O => \N__58993\,
            I => \N__58990\
        );

    \I__12556\ : InMux
    port map (
            O => \N__58990\,
            I => \N__58987\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__58987\,
            I => \N__58984\
        );

    \I__12554\ : Span4Mux_h
    port map (
            O => \N__58984\,
            I => \N__58980\
        );

    \I__12553\ : InMux
    port map (
            O => \N__58983\,
            I => \N__58977\
        );

    \I__12552\ : Span4Mux_v
    port map (
            O => \N__58980\,
            I => \N__58972\
        );

    \I__12551\ : LocalMux
    port map (
            O => \N__58977\,
            I => \N__58972\
        );

    \I__12550\ : Span4Mux_h
    port map (
            O => \N__58972\,
            I => \N__58969\
        );

    \I__12549\ : Odrv4
    port map (
            O => \N__58969\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n741\
        );

    \I__12548\ : InMux
    port map (
            O => \N__58966\,
            I => \N__58963\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__58963\,
            I => \N__58960\
        );

    \I__12546\ : Span12Mux_v
    port map (
            O => \N__58960\,
            I => \N__58957\
        );

    \I__12545\ : Odrv12
    port map (
            O => \N__58957\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n742_adj_411\
        );

    \I__12544\ : InMux
    port map (
            O => \N__58954\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17549\
        );

    \I__12543\ : InMux
    port map (
            O => \N__58951\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410\
        );

    \I__12542\ : InMux
    port map (
            O => \N__58948\,
            I => \N__58945\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__58945\,
            I => \N__58942\
        );

    \I__12540\ : Span4Mux_v
    port map (
            O => \N__58942\,
            I => \N__58939\
        );

    \I__12539\ : Odrv4
    port map (
            O => \N__58939\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_CO\
        );

    \I__12538\ : InMux
    port map (
            O => \N__58936\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590\
        );

    \I__12537\ : CascadeMux
    port map (
            O => \N__58933\,
            I => \N__58930\
        );

    \I__12536\ : InMux
    port map (
            O => \N__58930\,
            I => \N__58927\
        );

    \I__12535\ : LocalMux
    port map (
            O => \N__58927\,
            I => \N__58924\
        );

    \I__12534\ : Span4Mux_v
    port map (
            O => \N__58924\,
            I => \N__58921\
        );

    \I__12533\ : Span4Mux_v
    port map (
            O => \N__58921\,
            I => \N__58918\
        );

    \I__12532\ : Odrv4
    port map (
            O => \N__58918\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_CO\
        );

    \I__12531\ : CascadeMux
    port map (
            O => \N__58915\,
            I => \N__58912\
        );

    \I__12530\ : InMux
    port map (
            O => \N__58912\,
            I => \N__58896\
        );

    \I__12529\ : CascadeMux
    port map (
            O => \N__58911\,
            I => \N__58892\
        );

    \I__12528\ : CascadeMux
    port map (
            O => \N__58910\,
            I => \N__58888\
        );

    \I__12527\ : CascadeMux
    port map (
            O => \N__58909\,
            I => \N__58884\
        );

    \I__12526\ : CascadeMux
    port map (
            O => \N__58908\,
            I => \N__58881\
        );

    \I__12525\ : CascadeMux
    port map (
            O => \N__58907\,
            I => \N__58878\
        );

    \I__12524\ : CascadeMux
    port map (
            O => \N__58906\,
            I => \N__58875\
        );

    \I__12523\ : CascadeMux
    port map (
            O => \N__58905\,
            I => \N__58871\
        );

    \I__12522\ : CascadeMux
    port map (
            O => \N__58904\,
            I => \N__58867\
        );

    \I__12521\ : CascadeMux
    port map (
            O => \N__58903\,
            I => \N__58861\
        );

    \I__12520\ : CascadeMux
    port map (
            O => \N__58902\,
            I => \N__58857\
        );

    \I__12519\ : CascadeMux
    port map (
            O => \N__58901\,
            I => \N__58853\
        );

    \I__12518\ : CascadeMux
    port map (
            O => \N__58900\,
            I => \N__58849\
        );

    \I__12517\ : CascadeMux
    port map (
            O => \N__58899\,
            I => \N__58846\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__58896\,
            I => \N__58842\
        );

    \I__12515\ : InMux
    port map (
            O => \N__58895\,
            I => \N__58829\
        );

    \I__12514\ : InMux
    port map (
            O => \N__58892\,
            I => \N__58829\
        );

    \I__12513\ : InMux
    port map (
            O => \N__58891\,
            I => \N__58829\
        );

    \I__12512\ : InMux
    port map (
            O => \N__58888\,
            I => \N__58829\
        );

    \I__12511\ : InMux
    port map (
            O => \N__58887\,
            I => \N__58829\
        );

    \I__12510\ : InMux
    port map (
            O => \N__58884\,
            I => \N__58829\
        );

    \I__12509\ : InMux
    port map (
            O => \N__58881\,
            I => \N__58826\
        );

    \I__12508\ : InMux
    port map (
            O => \N__58878\,
            I => \N__58823\
        );

    \I__12507\ : InMux
    port map (
            O => \N__58875\,
            I => \N__58820\
        );

    \I__12506\ : CascadeMux
    port map (
            O => \N__58874\,
            I => \N__58817\
        );

    \I__12505\ : InMux
    port map (
            O => \N__58871\,
            I => \N__58814\
        );

    \I__12504\ : CascadeMux
    port map (
            O => \N__58870\,
            I => \N__58811\
        );

    \I__12503\ : InMux
    port map (
            O => \N__58867\,
            I => \N__58807\
        );

    \I__12502\ : InMux
    port map (
            O => \N__58866\,
            I => \N__58804\
        );

    \I__12501\ : InMux
    port map (
            O => \N__58865\,
            I => \N__58801\
        );

    \I__12500\ : InMux
    port map (
            O => \N__58864\,
            I => \N__58784\
        );

    \I__12499\ : InMux
    port map (
            O => \N__58861\,
            I => \N__58784\
        );

    \I__12498\ : InMux
    port map (
            O => \N__58860\,
            I => \N__58784\
        );

    \I__12497\ : InMux
    port map (
            O => \N__58857\,
            I => \N__58784\
        );

    \I__12496\ : InMux
    port map (
            O => \N__58856\,
            I => \N__58784\
        );

    \I__12495\ : InMux
    port map (
            O => \N__58853\,
            I => \N__58784\
        );

    \I__12494\ : InMux
    port map (
            O => \N__58852\,
            I => \N__58784\
        );

    \I__12493\ : InMux
    port map (
            O => \N__58849\,
            I => \N__58784\
        );

    \I__12492\ : InMux
    port map (
            O => \N__58846\,
            I => \N__58781\
        );

    \I__12491\ : CascadeMux
    port map (
            O => \N__58845\,
            I => \N__58777\
        );

    \I__12490\ : Span4Mux_v
    port map (
            O => \N__58842\,
            I => \N__58772\
        );

    \I__12489\ : LocalMux
    port map (
            O => \N__58829\,
            I => \N__58772\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__58826\,
            I => \N__58765\
        );

    \I__12487\ : LocalMux
    port map (
            O => \N__58823\,
            I => \N__58765\
        );

    \I__12486\ : LocalMux
    port map (
            O => \N__58820\,
            I => \N__58765\
        );

    \I__12485\ : InMux
    port map (
            O => \N__58817\,
            I => \N__58762\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__58814\,
            I => \N__58759\
        );

    \I__12483\ : InMux
    port map (
            O => \N__58811\,
            I => \N__58756\
        );

    \I__12482\ : CascadeMux
    port map (
            O => \N__58810\,
            I => \N__58752\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__58807\,
            I => \N__58747\
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__58804\,
            I => \N__58747\
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__58801\,
            I => \N__58740\
        );

    \I__12478\ : LocalMux
    port map (
            O => \N__58784\,
            I => \N__58740\
        );

    \I__12477\ : LocalMux
    port map (
            O => \N__58781\,
            I => \N__58740\
        );

    \I__12476\ : InMux
    port map (
            O => \N__58780\,
            I => \N__58737\
        );

    \I__12475\ : InMux
    port map (
            O => \N__58777\,
            I => \N__58734\
        );

    \I__12474\ : Span4Mux_v
    port map (
            O => \N__58772\,
            I => \N__58731\
        );

    \I__12473\ : Span4Mux_v
    port map (
            O => \N__58765\,
            I => \N__58722\
        );

    \I__12472\ : LocalMux
    port map (
            O => \N__58762\,
            I => \N__58722\
        );

    \I__12471\ : Span4Mux_h
    port map (
            O => \N__58759\,
            I => \N__58722\
        );

    \I__12470\ : LocalMux
    port map (
            O => \N__58756\,
            I => \N__58722\
        );

    \I__12469\ : InMux
    port map (
            O => \N__58755\,
            I => \N__58719\
        );

    \I__12468\ : InMux
    port map (
            O => \N__58752\,
            I => \N__58716\
        );

    \I__12467\ : Span4Mux_v
    port map (
            O => \N__58747\,
            I => \N__58707\
        );

    \I__12466\ : Span4Mux_h
    port map (
            O => \N__58740\,
            I => \N__58707\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__58737\,
            I => \N__58707\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__58734\,
            I => \N__58707\
        );

    \I__12463\ : Span4Mux_h
    port map (
            O => \N__58731\,
            I => \N__58698\
        );

    \I__12462\ : Span4Mux_v
    port map (
            O => \N__58722\,
            I => \N__58698\
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__58719\,
            I => \N__58698\
        );

    \I__12460\ : LocalMux
    port map (
            O => \N__58716\,
            I => \N__58698\
        );

    \I__12459\ : Span4Mux_v
    port map (
            O => \N__58707\,
            I => \N__58695\
        );

    \I__12458\ : Span4Mux_v
    port map (
            O => \N__58698\,
            I => \N__58692\
        );

    \I__12457\ : Odrv4
    port map (
            O => \N__58695\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n105\
        );

    \I__12456\ : Odrv4
    port map (
            O => \N__58692\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n105\
        );

    \I__12455\ : CascadeMux
    port map (
            O => \N__58687\,
            I => \N__58684\
        );

    \I__12454\ : InMux
    port map (
            O => \N__58684\,
            I => \N__58681\
        );

    \I__12453\ : LocalMux
    port map (
            O => \N__58681\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n57_adj_491\
        );

    \I__12452\ : InMux
    port map (
            O => \N__58678\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17536\
        );

    \I__12451\ : InMux
    port map (
            O => \N__58675\,
            I => \N__58672\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__58672\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n106_adj_509\
        );

    \I__12449\ : InMux
    port map (
            O => \N__58669\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17537\
        );

    \I__12448\ : CascadeMux
    port map (
            O => \N__58666\,
            I => \N__58663\
        );

    \I__12447\ : InMux
    port map (
            O => \N__58663\,
            I => \N__58660\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__58660\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n155\
        );

    \I__12445\ : InMux
    port map (
            O => \N__58657\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17538\
        );

    \I__12444\ : InMux
    port map (
            O => \N__58654\,
            I => \N__58651\
        );

    \I__12443\ : LocalMux
    port map (
            O => \N__58651\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n204\
        );

    \I__12442\ : InMux
    port map (
            O => \N__58648\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17539\
        );

    \I__12441\ : CascadeMux
    port map (
            O => \N__58645\,
            I => \N__58642\
        );

    \I__12440\ : InMux
    port map (
            O => \N__58642\,
            I => \N__58639\
        );

    \I__12439\ : LocalMux
    port map (
            O => \N__58639\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n253_adj_464\
        );

    \I__12438\ : InMux
    port map (
            O => \N__58636\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17540\
        );

    \I__12437\ : InMux
    port map (
            O => \N__58633\,
            I => \N__58630\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__58630\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n302\
        );

    \I__12435\ : InMux
    port map (
            O => \N__58627\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17541\
        );

    \I__12434\ : CascadeMux
    port map (
            O => \N__58624\,
            I => \N__58621\
        );

    \I__12433\ : InMux
    port map (
            O => \N__58621\,
            I => \N__58618\
        );

    \I__12432\ : LocalMux
    port map (
            O => \N__58618\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n351_adj_396\
        );

    \I__12431\ : CascadeMux
    port map (
            O => \N__58615\,
            I => \N__58612\
        );

    \I__12430\ : InMux
    port map (
            O => \N__58612\,
            I => \N__58609\
        );

    \I__12429\ : LocalMux
    port map (
            O => \N__58609\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n375_adj_587\
        );

    \I__12428\ : InMux
    port map (
            O => \N__58606\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18300\
        );

    \I__12427\ : CascadeMux
    port map (
            O => \N__58603\,
            I => \N__58600\
        );

    \I__12426\ : InMux
    port map (
            O => \N__58600\,
            I => \N__58597\
        );

    \I__12425\ : LocalMux
    port map (
            O => \N__58597\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n424_adj_586\
        );

    \I__12424\ : InMux
    port map (
            O => \N__58594\,
            I => \bfn_21_29_0_\
        );

    \I__12423\ : InMux
    port map (
            O => \N__58591\,
            I => \N__58588\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__58588\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n473_adj_585\
        );

    \I__12421\ : InMux
    port map (
            O => \N__58585\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18302\
        );

    \I__12420\ : InMux
    port map (
            O => \N__58582\,
            I => \N__58579\
        );

    \I__12419\ : LocalMux
    port map (
            O => \N__58579\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n522_adj_584\
        );

    \I__12418\ : InMux
    port map (
            O => \N__58576\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18303\
        );

    \I__12417\ : InMux
    port map (
            O => \N__58573\,
            I => \N__58570\
        );

    \I__12416\ : LocalMux
    port map (
            O => \N__58570\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n571\
        );

    \I__12415\ : InMux
    port map (
            O => \N__58567\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18304\
        );

    \I__12414\ : InMux
    port map (
            O => \N__58564\,
            I => \N__58561\
        );

    \I__12413\ : LocalMux
    port map (
            O => \N__58561\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n620\
        );

    \I__12412\ : InMux
    port map (
            O => \N__58558\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18305\
        );

    \I__12411\ : CascadeMux
    port map (
            O => \N__58555\,
            I => \N__58552\
        );

    \I__12410\ : InMux
    port map (
            O => \N__58552\,
            I => \N__58549\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__58549\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n669\
        );

    \I__12408\ : InMux
    port map (
            O => \N__58546\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18306\
        );

    \I__12407\ : CascadeMux
    port map (
            O => \N__58543\,
            I => \N__58540\
        );

    \I__12406\ : InMux
    port map (
            O => \N__58540\,
            I => \N__58537\
        );

    \I__12405\ : LocalMux
    port map (
            O => \N__58537\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n718\
        );

    \I__12404\ : InMux
    port map (
            O => \N__58534\,
            I => \N__58531\
        );

    \I__12403\ : LocalMux
    port map (
            O => \N__58531\,
            I => \N__58528\
        );

    \I__12402\ : Span12Mux_v
    port map (
            O => \N__58528\,
            I => \N__58525\
        );

    \I__12401\ : Odrv12
    port map (
            O => \N__58525\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n774_adj_589\
        );

    \I__12400\ : InMux
    port map (
            O => \N__58522\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18307\
        );

    \I__12399\ : CascadeMux
    port map (
            O => \N__58519\,
            I => \N__58516\
        );

    \I__12398\ : InMux
    port map (
            O => \N__58516\,
            I => \N__58513\
        );

    \I__12397\ : LocalMux
    port map (
            O => \N__58513\,
            I => \N__58509\
        );

    \I__12396\ : InMux
    port map (
            O => \N__58512\,
            I => \N__58506\
        );

    \I__12395\ : Sp12to4
    port map (
            O => \N__58509\,
            I => \N__58503\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__58506\,
            I => \N__58500\
        );

    \I__12393\ : Span12Mux_s11_v
    port map (
            O => \N__58503\,
            I => \N__58497\
        );

    \I__12392\ : Span12Mux_s11_v
    port map (
            O => \N__58500\,
            I => \N__58494\
        );

    \I__12391\ : Odrv12
    port map (
            O => \N__58497\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30\
        );

    \I__12390\ : Odrv12
    port map (
            O => \N__58494\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30\
        );

    \I__12389\ : InMux
    port map (
            O => \N__58489\,
            I => \N__58482\
        );

    \I__12388\ : InMux
    port map (
            O => \N__58488\,
            I => \N__58482\
        );

    \I__12387\ : InMux
    port map (
            O => \N__58487\,
            I => \N__58479\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__58482\,
            I => \N__58476\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__58479\,
            I => \N__58473\
        );

    \I__12384\ : Span4Mux_h
    port map (
            O => \N__58476\,
            I => \N__58470\
        );

    \I__12383\ : Span12Mux_h
    port map (
            O => \N__58473\,
            I => \N__58467\
        );

    \I__12382\ : Span4Mux_v
    port map (
            O => \N__58470\,
            I => \N__58464\
        );

    \I__12381\ : Odrv12
    port map (
            O => \N__58467\,
            I => \Add_add_temp_34_adj_2386\
        );

    \I__12380\ : Odrv4
    port map (
            O => \N__58464\,
            I => \Add_add_temp_34_adj_2386\
        );

    \I__12379\ : InMux
    port map (
            O => \N__58459\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15942\
        );

    \I__12378\ : InMux
    port map (
            O => \N__58456\,
            I => \N__58453\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__58453\,
            I => \N__58447\
        );

    \I__12376\ : CascadeMux
    port map (
            O => \N__58452\,
            I => \N__58443\
        );

    \I__12375\ : CascadeMux
    port map (
            O => \N__58451\,
            I => \N__58439\
        );

    \I__12374\ : CascadeMux
    port map (
            O => \N__58450\,
            I => \N__58435\
        );

    \I__12373\ : Span4Mux_v
    port map (
            O => \N__58447\,
            I => \N__58430\
        );

    \I__12372\ : InMux
    port map (
            O => \N__58446\,
            I => \N__58415\
        );

    \I__12371\ : InMux
    port map (
            O => \N__58443\,
            I => \N__58415\
        );

    \I__12370\ : InMux
    port map (
            O => \N__58442\,
            I => \N__58415\
        );

    \I__12369\ : InMux
    port map (
            O => \N__58439\,
            I => \N__58415\
        );

    \I__12368\ : InMux
    port map (
            O => \N__58438\,
            I => \N__58415\
        );

    \I__12367\ : InMux
    port map (
            O => \N__58435\,
            I => \N__58415\
        );

    \I__12366\ : InMux
    port map (
            O => \N__58434\,
            I => \N__58415\
        );

    \I__12365\ : InMux
    port map (
            O => \N__58433\,
            I => \N__58412\
        );

    \I__12364\ : Odrv4
    port map (
            O => \N__58430\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31\
        );

    \I__12363\ : LocalMux
    port map (
            O => \N__58415\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31\
        );

    \I__12362\ : LocalMux
    port map (
            O => \N__58412\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31\
        );

    \I__12361\ : CascadeMux
    port map (
            O => \N__58405\,
            I => \N__58400\
        );

    \I__12360\ : CascadeMux
    port map (
            O => \N__58404\,
            I => \N__58396\
        );

    \I__12359\ : CascadeMux
    port map (
            O => \N__58403\,
            I => \N__58392\
        );

    \I__12358\ : InMux
    port map (
            O => \N__58400\,
            I => \N__58381\
        );

    \I__12357\ : InMux
    port map (
            O => \N__58399\,
            I => \N__58381\
        );

    \I__12356\ : InMux
    port map (
            O => \N__58396\,
            I => \N__58381\
        );

    \I__12355\ : InMux
    port map (
            O => \N__58395\,
            I => \N__58381\
        );

    \I__12354\ : InMux
    port map (
            O => \N__58392\,
            I => \N__58381\
        );

    \I__12353\ : LocalMux
    port map (
            O => \N__58381\,
            I => \N__58378\
        );

    \I__12352\ : Span4Mux_v
    port map (
            O => \N__58378\,
            I => \N__58375\
        );

    \I__12351\ : Odrv4
    port map (
            O => \N__58375\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_31\
        );

    \I__12350\ : InMux
    port map (
            O => \N__58372\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15943\
        );

    \I__12349\ : InMux
    port map (
            O => \N__58369\,
            I => \N__58364\
        );

    \I__12348\ : InMux
    port map (
            O => \N__58368\,
            I => \N__58361\
        );

    \I__12347\ : InMux
    port map (
            O => \N__58367\,
            I => \N__58358\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__58364\,
            I => \N__58353\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__58361\,
            I => \N__58353\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__58358\,
            I => \N__58350\
        );

    \I__12343\ : Span4Mux_v
    port map (
            O => \N__58353\,
            I => \N__58347\
        );

    \I__12342\ : Span4Mux_v
    port map (
            O => \N__58350\,
            I => \N__58344\
        );

    \I__12341\ : Odrv4
    port map (
            O => \N__58347\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31\
        );

    \I__12340\ : Odrv4
    port map (
            O => \N__58344\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31\
        );

    \I__12339\ : InMux
    port map (
            O => \N__58339\,
            I => \N__58336\
        );

    \I__12338\ : LocalMux
    port map (
            O => \N__58336\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n81\
        );

    \I__12337\ : InMux
    port map (
            O => \N__58333\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18294\
        );

    \I__12336\ : InMux
    port map (
            O => \N__58330\,
            I => \N__58327\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__58327\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n130\
        );

    \I__12334\ : InMux
    port map (
            O => \N__58324\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18295\
        );

    \I__12333\ : InMux
    port map (
            O => \N__58321\,
            I => \N__58318\
        );

    \I__12332\ : LocalMux
    port map (
            O => \N__58318\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n179\
        );

    \I__12331\ : InMux
    port map (
            O => \N__58315\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18296\
        );

    \I__12330\ : CascadeMux
    port map (
            O => \N__58312\,
            I => \N__58309\
        );

    \I__12329\ : InMux
    port map (
            O => \N__58309\,
            I => \N__58306\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__58306\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n228\
        );

    \I__12327\ : InMux
    port map (
            O => \N__58303\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18297\
        );

    \I__12326\ : InMux
    port map (
            O => \N__58300\,
            I => \N__58297\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__58297\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n277\
        );

    \I__12324\ : InMux
    port map (
            O => \N__58294\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18298\
        );

    \I__12323\ : CascadeMux
    port map (
            O => \N__58291\,
            I => \N__58288\
        );

    \I__12322\ : InMux
    port map (
            O => \N__58288\,
            I => \N__58285\
        );

    \I__12321\ : LocalMux
    port map (
            O => \N__58285\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n326_adj_588\
        );

    \I__12320\ : InMux
    port map (
            O => \N__58282\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18299\
        );

    \I__12319\ : InMux
    port map (
            O => \N__58279\,
            I => \N__58275\
        );

    \I__12318\ : InMux
    port map (
            O => \N__58278\,
            I => \N__58272\
        );

    \I__12317\ : LocalMux
    port map (
            O => \N__58275\,
            I => \N__58269\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__58272\,
            I => \N__58266\
        );

    \I__12315\ : Span4Mux_v
    port map (
            O => \N__58269\,
            I => \N__58263\
        );

    \I__12314\ : Span4Mux_h
    port map (
            O => \N__58266\,
            I => \N__58260\
        );

    \I__12313\ : Odrv4
    port map (
            O => \N__58263\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23\
        );

    \I__12312\ : Odrv4
    port map (
            O => \N__58260\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23\
        );

    \I__12311\ : CascadeMux
    port map (
            O => \N__58255\,
            I => \N__58252\
        );

    \I__12310\ : InMux
    port map (
            O => \N__58252\,
            I => \N__58249\
        );

    \I__12309\ : LocalMux
    port map (
            O => \N__58249\,
            I => \N__58246\
        );

    \I__12308\ : Span4Mux_h
    port map (
            O => \N__58246\,
            I => \N__58243\
        );

    \I__12307\ : Odrv4
    port map (
            O => \N__58243\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_27\
        );

    \I__12306\ : InMux
    port map (
            O => \N__58240\,
            I => \N__58235\
        );

    \I__12305\ : InMux
    port map (
            O => \N__58239\,
            I => \N__58232\
        );

    \I__12304\ : InMux
    port map (
            O => \N__58238\,
            I => \N__58229\
        );

    \I__12303\ : LocalMux
    port map (
            O => \N__58235\,
            I => \N__58222\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__58232\,
            I => \N__58222\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__58229\,
            I => \N__58222\
        );

    \I__12300\ : Span4Mux_v
    port map (
            O => \N__58222\,
            I => \N__58219\
        );

    \I__12299\ : Odrv4
    port map (
            O => \N__58219\,
            I => \Add_add_temp_27_adj_2393\
        );

    \I__12298\ : InMux
    port map (
            O => \N__58216\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15935\
        );

    \I__12297\ : CascadeMux
    port map (
            O => \N__58213\,
            I => \N__58209\
        );

    \I__12296\ : InMux
    port map (
            O => \N__58212\,
            I => \N__58206\
        );

    \I__12295\ : InMux
    port map (
            O => \N__58209\,
            I => \N__58203\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__58206\,
            I => \N__58200\
        );

    \I__12293\ : LocalMux
    port map (
            O => \N__58203\,
            I => \N__58197\
        );

    \I__12292\ : Span4Mux_v
    port map (
            O => \N__58200\,
            I => \N__58194\
        );

    \I__12291\ : Span4Mux_v
    port map (
            O => \N__58197\,
            I => \N__58191\
        );

    \I__12290\ : Odrv4
    port map (
            O => \N__58194\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24\
        );

    \I__12289\ : Odrv4
    port map (
            O => \N__58191\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24\
        );

    \I__12288\ : CascadeMux
    port map (
            O => \N__58186\,
            I => \N__58183\
        );

    \I__12287\ : InMux
    port map (
            O => \N__58183\,
            I => \N__58180\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__58180\,
            I => \N__58177\
        );

    \I__12285\ : Span4Mux_v
    port map (
            O => \N__58177\,
            I => \N__58174\
        );

    \I__12284\ : Odrv4
    port map (
            O => \N__58174\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_28\
        );

    \I__12283\ : InMux
    port map (
            O => \N__58171\,
            I => \N__58164\
        );

    \I__12282\ : InMux
    port map (
            O => \N__58170\,
            I => \N__58164\
        );

    \I__12281\ : InMux
    port map (
            O => \N__58169\,
            I => \N__58161\
        );

    \I__12280\ : LocalMux
    port map (
            O => \N__58164\,
            I => \N__58156\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__58161\,
            I => \N__58156\
        );

    \I__12278\ : Span4Mux_v
    port map (
            O => \N__58156\,
            I => \N__58153\
        );

    \I__12277\ : Odrv4
    port map (
            O => \N__58153\,
            I => \Add_add_temp_28_adj_2392\
        );

    \I__12276\ : InMux
    port map (
            O => \N__58150\,
            I => \bfn_21_26_0_\
        );

    \I__12275\ : InMux
    port map (
            O => \N__58147\,
            I => \N__58144\
        );

    \I__12274\ : LocalMux
    port map (
            O => \N__58144\,
            I => \N__58141\
        );

    \I__12273\ : Span4Mux_h
    port map (
            O => \N__58141\,
            I => \N__58137\
        );

    \I__12272\ : InMux
    port map (
            O => \N__58140\,
            I => \N__58134\
        );

    \I__12271\ : Sp12to4
    port map (
            O => \N__58137\,
            I => \N__58129\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__58134\,
            I => \N__58129\
        );

    \I__12269\ : Odrv12
    port map (
            O => \N__58129\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_25\
        );

    \I__12268\ : CascadeMux
    port map (
            O => \N__58126\,
            I => \N__58123\
        );

    \I__12267\ : InMux
    port map (
            O => \N__58123\,
            I => \N__58120\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__58120\,
            I => \N__58117\
        );

    \I__12265\ : Span4Mux_v
    port map (
            O => \N__58117\,
            I => \N__58114\
        );

    \I__12264\ : Odrv4
    port map (
            O => \N__58114\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_29\
        );

    \I__12263\ : InMux
    port map (
            O => \N__58111\,
            I => \N__58106\
        );

    \I__12262\ : InMux
    port map (
            O => \N__58110\,
            I => \N__58101\
        );

    \I__12261\ : InMux
    port map (
            O => \N__58109\,
            I => \N__58101\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__58106\,
            I => \N__58098\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__58101\,
            I => \N__58095\
        );

    \I__12258\ : Sp12to4
    port map (
            O => \N__58098\,
            I => \N__58092\
        );

    \I__12257\ : Span4Mux_v
    port map (
            O => \N__58095\,
            I => \N__58089\
        );

    \I__12256\ : Odrv12
    port map (
            O => \N__58092\,
            I => \Add_add_temp_29_adj_2391\
        );

    \I__12255\ : Odrv4
    port map (
            O => \N__58089\,
            I => \Add_add_temp_29_adj_2391\
        );

    \I__12254\ : InMux
    port map (
            O => \N__58084\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15937\
        );

    \I__12253\ : InMux
    port map (
            O => \N__58081\,
            I => \N__58077\
        );

    \I__12252\ : InMux
    port map (
            O => \N__58080\,
            I => \N__58074\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__58077\,
            I => \N__58071\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__58074\,
            I => \N__58068\
        );

    \I__12249\ : Span12Mux_v
    port map (
            O => \N__58071\,
            I => \N__58065\
        );

    \I__12248\ : Span4Mux_v
    port map (
            O => \N__58068\,
            I => \N__58062\
        );

    \I__12247\ : Odrv12
    port map (
            O => \N__58065\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26\
        );

    \I__12246\ : Odrv4
    port map (
            O => \N__58062\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26\
        );

    \I__12245\ : CascadeMux
    port map (
            O => \N__58057\,
            I => \N__58054\
        );

    \I__12244\ : InMux
    port map (
            O => \N__58054\,
            I => \N__58051\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__58051\,
            I => \N__58048\
        );

    \I__12242\ : Span4Mux_v
    port map (
            O => \N__58048\,
            I => \N__58045\
        );

    \I__12241\ : Odrv4
    port map (
            O => \N__58045\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_30\
        );

    \I__12240\ : InMux
    port map (
            O => \N__58042\,
            I => \N__58035\
        );

    \I__12239\ : InMux
    port map (
            O => \N__58041\,
            I => \N__58035\
        );

    \I__12238\ : InMux
    port map (
            O => \N__58040\,
            I => \N__58032\
        );

    \I__12237\ : LocalMux
    port map (
            O => \N__58035\,
            I => \N__58029\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__58032\,
            I => \N__58026\
        );

    \I__12235\ : Span4Mux_v
    port map (
            O => \N__58029\,
            I => \N__58021\
        );

    \I__12234\ : Span4Mux_v
    port map (
            O => \N__58026\,
            I => \N__58021\
        );

    \I__12233\ : Odrv4
    port map (
            O => \N__58021\,
            I => \Add_add_temp_30_adj_2390\
        );

    \I__12232\ : InMux
    port map (
            O => \N__58018\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15938\
        );

    \I__12231\ : InMux
    port map (
            O => \N__58015\,
            I => \N__58012\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__58012\,
            I => \N__58008\
        );

    \I__12229\ : CascadeMux
    port map (
            O => \N__58011\,
            I => \N__58005\
        );

    \I__12228\ : Span4Mux_v
    port map (
            O => \N__58008\,
            I => \N__58002\
        );

    \I__12227\ : InMux
    port map (
            O => \N__58005\,
            I => \N__57999\
        );

    \I__12226\ : Span4Mux_h
    port map (
            O => \N__58002\,
            I => \N__57994\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__57999\,
            I => \N__57994\
        );

    \I__12224\ : Span4Mux_v
    port map (
            O => \N__57994\,
            I => \N__57991\
        );

    \I__12223\ : Odrv4
    port map (
            O => \N__57991\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_27\
        );

    \I__12222\ : InMux
    port map (
            O => \N__57988\,
            I => \N__57981\
        );

    \I__12221\ : InMux
    port map (
            O => \N__57987\,
            I => \N__57981\
        );

    \I__12220\ : InMux
    port map (
            O => \N__57986\,
            I => \N__57978\
        );

    \I__12219\ : LocalMux
    port map (
            O => \N__57981\,
            I => \N__57973\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__57978\,
            I => \N__57973\
        );

    \I__12217\ : Span4Mux_v
    port map (
            O => \N__57973\,
            I => \N__57970\
        );

    \I__12216\ : Odrv4
    port map (
            O => \N__57970\,
            I => \Add_add_temp_31_adj_2389\
        );

    \I__12215\ : InMux
    port map (
            O => \N__57967\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15939\
        );

    \I__12214\ : InMux
    port map (
            O => \N__57964\,
            I => \N__57960\
        );

    \I__12213\ : CascadeMux
    port map (
            O => \N__57963\,
            I => \N__57957\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__57960\,
            I => \N__57954\
        );

    \I__12211\ : InMux
    port map (
            O => \N__57957\,
            I => \N__57951\
        );

    \I__12210\ : Span4Mux_v
    port map (
            O => \N__57954\,
            I => \N__57948\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__57951\,
            I => \N__57945\
        );

    \I__12208\ : Odrv4
    port map (
            O => \N__57948\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28\
        );

    \I__12207\ : Odrv12
    port map (
            O => \N__57945\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28\
        );

    \I__12206\ : InMux
    port map (
            O => \N__57940\,
            I => \N__57935\
        );

    \I__12205\ : InMux
    port map (
            O => \N__57939\,
            I => \N__57932\
        );

    \I__12204\ : InMux
    port map (
            O => \N__57938\,
            I => \N__57929\
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__57935\,
            I => \N__57922\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__57932\,
            I => \N__57922\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__57929\,
            I => \N__57922\
        );

    \I__12200\ : Span4Mux_v
    port map (
            O => \N__57922\,
            I => \N__57919\
        );

    \I__12199\ : Odrv4
    port map (
            O => \N__57919\,
            I => \Add_add_temp_32_adj_2388\
        );

    \I__12198\ : InMux
    port map (
            O => \N__57916\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15940\
        );

    \I__12197\ : InMux
    port map (
            O => \N__57913\,
            I => \N__57910\
        );

    \I__12196\ : LocalMux
    port map (
            O => \N__57910\,
            I => \N__57906\
        );

    \I__12195\ : InMux
    port map (
            O => \N__57909\,
            I => \N__57903\
        );

    \I__12194\ : Span4Mux_v
    port map (
            O => \N__57906\,
            I => \N__57898\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__57903\,
            I => \N__57898\
        );

    \I__12192\ : Span4Mux_h
    port map (
            O => \N__57898\,
            I => \N__57895\
        );

    \I__12191\ : Span4Mux_v
    port map (
            O => \N__57895\,
            I => \N__57892\
        );

    \I__12190\ : Odrv4
    port map (
            O => \N__57892\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_29\
        );

    \I__12189\ : CascadeMux
    port map (
            O => \N__57889\,
            I => \N__57884\
        );

    \I__12188\ : InMux
    port map (
            O => \N__57888\,
            I => \N__57879\
        );

    \I__12187\ : InMux
    port map (
            O => \N__57887\,
            I => \N__57879\
        );

    \I__12186\ : InMux
    port map (
            O => \N__57884\,
            I => \N__57876\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__57879\,
            I => \N__57871\
        );

    \I__12184\ : LocalMux
    port map (
            O => \N__57876\,
            I => \N__57871\
        );

    \I__12183\ : Span12Mux_v
    port map (
            O => \N__57871\,
            I => \N__57868\
        );

    \I__12182\ : Odrv12
    port map (
            O => \N__57868\,
            I => \Add_add_temp_33_adj_2387\
        );

    \I__12181\ : InMux
    port map (
            O => \N__57865\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15941\
        );

    \I__12180\ : InMux
    port map (
            O => \N__57862\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15927\
        );

    \I__12179\ : InMux
    port map (
            O => \N__57859\,
            I => \N__57856\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__57856\,
            I => \N__57853\
        );

    \I__12177\ : Span4Mux_h
    port map (
            O => \N__57853\,
            I => \N__57849\
        );

    \I__12176\ : InMux
    port map (
            O => \N__57852\,
            I => \N__57846\
        );

    \I__12175\ : Odrv4
    port map (
            O => \N__57849\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16\
        );

    \I__12174\ : LocalMux
    port map (
            O => \N__57846\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16\
        );

    \I__12173\ : CascadeMux
    port map (
            O => \N__57841\,
            I => \N__57838\
        );

    \I__12172\ : InMux
    port map (
            O => \N__57838\,
            I => \N__57835\
        );

    \I__12171\ : LocalMux
    port map (
            O => \N__57835\,
            I => \N__57832\
        );

    \I__12170\ : Span4Mux_v
    port map (
            O => \N__57832\,
            I => \N__57829\
        );

    \I__12169\ : Span4Mux_h
    port map (
            O => \N__57829\,
            I => \N__57826\
        );

    \I__12168\ : Odrv4
    port map (
            O => \N__57826\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_20\
        );

    \I__12167\ : InMux
    port map (
            O => \N__57823\,
            I => \bfn_21_25_0_\
        );

    \I__12166\ : InMux
    port map (
            O => \N__57820\,
            I => \N__57817\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__57817\,
            I => \N__57814\
        );

    \I__12164\ : Span4Mux_h
    port map (
            O => \N__57814\,
            I => \N__57810\
        );

    \I__12163\ : InMux
    port map (
            O => \N__57813\,
            I => \N__57807\
        );

    \I__12162\ : Odrv4
    port map (
            O => \N__57810\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__57807\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17\
        );

    \I__12160\ : CascadeMux
    port map (
            O => \N__57802\,
            I => \N__57799\
        );

    \I__12159\ : InMux
    port map (
            O => \N__57799\,
            I => \N__57796\
        );

    \I__12158\ : LocalMux
    port map (
            O => \N__57796\,
            I => \N__57793\
        );

    \I__12157\ : Span4Mux_v
    port map (
            O => \N__57793\,
            I => \N__57790\
        );

    \I__12156\ : Odrv4
    port map (
            O => \N__57790\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_21\
        );

    \I__12155\ : InMux
    port map (
            O => \N__57787\,
            I => \N__57782\
        );

    \I__12154\ : InMux
    port map (
            O => \N__57786\,
            I => \N__57779\
        );

    \I__12153\ : InMux
    port map (
            O => \N__57785\,
            I => \N__57776\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__57782\,
            I => \N__57773\
        );

    \I__12151\ : LocalMux
    port map (
            O => \N__57779\,
            I => \N__57770\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__57776\,
            I => \N__57767\
        );

    \I__12149\ : Span4Mux_v
    port map (
            O => \N__57773\,
            I => \N__57762\
        );

    \I__12148\ : Span4Mux_h
    port map (
            O => \N__57770\,
            I => \N__57762\
        );

    \I__12147\ : Span4Mux_h
    port map (
            O => \N__57767\,
            I => \N__57759\
        );

    \I__12146\ : Odrv4
    port map (
            O => \N__57762\,
            I => \Add_add_temp_21_adj_2399\
        );

    \I__12145\ : Odrv4
    port map (
            O => \N__57759\,
            I => \Add_add_temp_21_adj_2399\
        );

    \I__12144\ : InMux
    port map (
            O => \N__57754\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15929\
        );

    \I__12143\ : InMux
    port map (
            O => \N__57751\,
            I => \N__57748\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__57748\,
            I => \N__57745\
        );

    \I__12141\ : Span4Mux_v
    port map (
            O => \N__57745\,
            I => \N__57741\
        );

    \I__12140\ : InMux
    port map (
            O => \N__57744\,
            I => \N__57738\
        );

    \I__12139\ : Odrv4
    port map (
            O => \N__57741\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__57738\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18\
        );

    \I__12137\ : CascadeMux
    port map (
            O => \N__57733\,
            I => \N__57730\
        );

    \I__12136\ : InMux
    port map (
            O => \N__57730\,
            I => \N__57727\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__57727\,
            I => \N__57724\
        );

    \I__12134\ : Span4Mux_v
    port map (
            O => \N__57724\,
            I => \N__57721\
        );

    \I__12133\ : Odrv4
    port map (
            O => \N__57721\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_22\
        );

    \I__12132\ : CascadeMux
    port map (
            O => \N__57718\,
            I => \N__57713\
        );

    \I__12131\ : InMux
    port map (
            O => \N__57717\,
            I => \N__57710\
        );

    \I__12130\ : InMux
    port map (
            O => \N__57716\,
            I => \N__57707\
        );

    \I__12129\ : InMux
    port map (
            O => \N__57713\,
            I => \N__57704\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__57710\,
            I => \N__57699\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__57707\,
            I => \N__57699\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__57704\,
            I => \N__57696\
        );

    \I__12125\ : Span4Mux_v
    port map (
            O => \N__57699\,
            I => \N__57693\
        );

    \I__12124\ : Odrv12
    port map (
            O => \N__57696\,
            I => \Add_add_temp_22_adj_2398\
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__57693\,
            I => \Add_add_temp_22_adj_2398\
        );

    \I__12122\ : InMux
    port map (
            O => \N__57688\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15930\
        );

    \I__12121\ : InMux
    port map (
            O => \N__57685\,
            I => \N__57681\
        );

    \I__12120\ : InMux
    port map (
            O => \N__57684\,
            I => \N__57678\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__57681\,
            I => \N__57675\
        );

    \I__12118\ : LocalMux
    port map (
            O => \N__57678\,
            I => \N__57672\
        );

    \I__12117\ : Span4Mux_h
    port map (
            O => \N__57675\,
            I => \N__57669\
        );

    \I__12116\ : Span4Mux_h
    port map (
            O => \N__57672\,
            I => \N__57666\
        );

    \I__12115\ : Sp12to4
    port map (
            O => \N__57669\,
            I => \N__57661\
        );

    \I__12114\ : Sp12to4
    port map (
            O => \N__57666\,
            I => \N__57661\
        );

    \I__12113\ : Odrv12
    port map (
            O => \N__57661\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_19\
        );

    \I__12112\ : CascadeMux
    port map (
            O => \N__57658\,
            I => \N__57655\
        );

    \I__12111\ : InMux
    port map (
            O => \N__57655\,
            I => \N__57652\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__57652\,
            I => \N__57649\
        );

    \I__12109\ : Span4Mux_v
    port map (
            O => \N__57649\,
            I => \N__57646\
        );

    \I__12108\ : Sp12to4
    port map (
            O => \N__57646\,
            I => \N__57643\
        );

    \I__12107\ : Odrv12
    port map (
            O => \N__57643\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_23\
        );

    \I__12106\ : InMux
    port map (
            O => \N__57640\,
            I => \N__57636\
        );

    \I__12105\ : InMux
    port map (
            O => \N__57639\,
            I => \N__57632\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__57636\,
            I => \N__57629\
        );

    \I__12103\ : InMux
    port map (
            O => \N__57635\,
            I => \N__57626\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__57632\,
            I => \N__57623\
        );

    \I__12101\ : Span4Mux_h
    port map (
            O => \N__57629\,
            I => \N__57620\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__57626\,
            I => \N__57615\
        );

    \I__12099\ : Span4Mux_h
    port map (
            O => \N__57623\,
            I => \N__57615\
        );

    \I__12098\ : Span4Mux_v
    port map (
            O => \N__57620\,
            I => \N__57612\
        );

    \I__12097\ : Span4Mux_v
    port map (
            O => \N__57615\,
            I => \N__57609\
        );

    \I__12096\ : Odrv4
    port map (
            O => \N__57612\,
            I => \Add_add_temp_23_adj_2397\
        );

    \I__12095\ : Odrv4
    port map (
            O => \N__57609\,
            I => \Add_add_temp_23_adj_2397\
        );

    \I__12094\ : InMux
    port map (
            O => \N__57604\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15931\
        );

    \I__12093\ : InMux
    port map (
            O => \N__57601\,
            I => \N__57597\
        );

    \I__12092\ : InMux
    port map (
            O => \N__57600\,
            I => \N__57594\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__57597\,
            I => \N__57591\
        );

    \I__12090\ : LocalMux
    port map (
            O => \N__57594\,
            I => \N__57588\
        );

    \I__12089\ : Span4Mux_v
    port map (
            O => \N__57591\,
            I => \N__57585\
        );

    \I__12088\ : Span4Mux_v
    port map (
            O => \N__57588\,
            I => \N__57582\
        );

    \I__12087\ : Odrv4
    port map (
            O => \N__57585\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20\
        );

    \I__12086\ : Odrv4
    port map (
            O => \N__57582\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20\
        );

    \I__12085\ : CascadeMux
    port map (
            O => \N__57577\,
            I => \N__57574\
        );

    \I__12084\ : InMux
    port map (
            O => \N__57574\,
            I => \N__57571\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__57571\,
            I => \N__57568\
        );

    \I__12082\ : Span4Mux_v
    port map (
            O => \N__57568\,
            I => \N__57565\
        );

    \I__12081\ : Odrv4
    port map (
            O => \N__57565\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_24\
        );

    \I__12080\ : InMux
    port map (
            O => \N__57562\,
            I => \N__57558\
        );

    \I__12079\ : InMux
    port map (
            O => \N__57561\,
            I => \N__57555\
        );

    \I__12078\ : LocalMux
    port map (
            O => \N__57558\,
            I => \N__57552\
        );

    \I__12077\ : LocalMux
    port map (
            O => \N__57555\,
            I => \N__57548\
        );

    \I__12076\ : Span4Mux_v
    port map (
            O => \N__57552\,
            I => \N__57545\
        );

    \I__12075\ : InMux
    port map (
            O => \N__57551\,
            I => \N__57542\
        );

    \I__12074\ : Sp12to4
    port map (
            O => \N__57548\,
            I => \N__57535\
        );

    \I__12073\ : Sp12to4
    port map (
            O => \N__57545\,
            I => \N__57535\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__57542\,
            I => \N__57535\
        );

    \I__12071\ : Odrv12
    port map (
            O => \N__57535\,
            I => \Add_add_temp_24_adj_2396\
        );

    \I__12070\ : InMux
    port map (
            O => \N__57532\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15932\
        );

    \I__12069\ : InMux
    port map (
            O => \N__57529\,
            I => \N__57526\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__57526\,
            I => \N__57522\
        );

    \I__12067\ : InMux
    port map (
            O => \N__57525\,
            I => \N__57519\
        );

    \I__12066\ : Span4Mux_h
    port map (
            O => \N__57522\,
            I => \N__57514\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__57519\,
            I => \N__57514\
        );

    \I__12064\ : Span4Mux_v
    port map (
            O => \N__57514\,
            I => \N__57511\
        );

    \I__12063\ : Odrv4
    port map (
            O => \N__57511\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_21\
        );

    \I__12062\ : CascadeMux
    port map (
            O => \N__57508\,
            I => \N__57505\
        );

    \I__12061\ : InMux
    port map (
            O => \N__57505\,
            I => \N__57502\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__57502\,
            I => \N__57499\
        );

    \I__12059\ : Span4Mux_h
    port map (
            O => \N__57499\,
            I => \N__57496\
        );

    \I__12058\ : Odrv4
    port map (
            O => \N__57496\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_25\
        );

    \I__12057\ : InMux
    port map (
            O => \N__57493\,
            I => \N__57488\
        );

    \I__12056\ : InMux
    port map (
            O => \N__57492\,
            I => \N__57485\
        );

    \I__12055\ : InMux
    port map (
            O => \N__57491\,
            I => \N__57482\
        );

    \I__12054\ : LocalMux
    port map (
            O => \N__57488\,
            I => \N__57479\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__57485\,
            I => \N__57474\
        );

    \I__12052\ : LocalMux
    port map (
            O => \N__57482\,
            I => \N__57474\
        );

    \I__12051\ : Span4Mux_h
    port map (
            O => \N__57479\,
            I => \N__57469\
        );

    \I__12050\ : Span4Mux_v
    port map (
            O => \N__57474\,
            I => \N__57469\
        );

    \I__12049\ : Odrv4
    port map (
            O => \N__57469\,
            I => \Add_add_temp_25_adj_2395\
        );

    \I__12048\ : InMux
    port map (
            O => \N__57466\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15933\
        );

    \I__12047\ : CascadeMux
    port map (
            O => \N__57463\,
            I => \N__57460\
        );

    \I__12046\ : InMux
    port map (
            O => \N__57460\,
            I => \N__57457\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__57457\,
            I => \N__57453\
        );

    \I__12044\ : InMux
    port map (
            O => \N__57456\,
            I => \N__57450\
        );

    \I__12043\ : Span4Mux_v
    port map (
            O => \N__57453\,
            I => \N__57447\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__57450\,
            I => \N__57444\
        );

    \I__12041\ : Odrv4
    port map (
            O => \N__57447\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22\
        );

    \I__12040\ : Odrv12
    port map (
            O => \N__57444\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22\
        );

    \I__12039\ : CascadeMux
    port map (
            O => \N__57439\,
            I => \N__57436\
        );

    \I__12038\ : InMux
    port map (
            O => \N__57436\,
            I => \N__57433\
        );

    \I__12037\ : LocalMux
    port map (
            O => \N__57433\,
            I => \N__57430\
        );

    \I__12036\ : Span12Mux_h
    port map (
            O => \N__57430\,
            I => \N__57427\
        );

    \I__12035\ : Odrv12
    port map (
            O => \N__57427\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_26\
        );

    \I__12034\ : CascadeMux
    port map (
            O => \N__57424\,
            I => \N__57421\
        );

    \I__12033\ : InMux
    port map (
            O => \N__57421\,
            I => \N__57416\
        );

    \I__12032\ : InMux
    port map (
            O => \N__57420\,
            I => \N__57411\
        );

    \I__12031\ : InMux
    port map (
            O => \N__57419\,
            I => \N__57411\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__57416\,
            I => \N__57408\
        );

    \I__12029\ : LocalMux
    port map (
            O => \N__57411\,
            I => \N__57405\
        );

    \I__12028\ : Span4Mux_h
    port map (
            O => \N__57408\,
            I => \N__57402\
        );

    \I__12027\ : Span4Mux_v
    port map (
            O => \N__57405\,
            I => \N__57399\
        );

    \I__12026\ : Span4Mux_v
    port map (
            O => \N__57402\,
            I => \N__57396\
        );

    \I__12025\ : Span4Mux_h
    port map (
            O => \N__57399\,
            I => \N__57393\
        );

    \I__12024\ : Odrv4
    port map (
            O => \N__57396\,
            I => \Add_add_temp_26_adj_2394\
        );

    \I__12023\ : Odrv4
    port map (
            O => \N__57393\,
            I => \Add_add_temp_26_adj_2394\
        );

    \I__12022\ : InMux
    port map (
            O => \N__57388\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15934\
        );

    \I__12021\ : InMux
    port map (
            O => \N__57385\,
            I => \N__57381\
        );

    \I__12020\ : InMux
    port map (
            O => \N__57384\,
            I => \N__57378\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__57381\,
            I => \N__57375\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__57378\,
            I => \N__57372\
        );

    \I__12017\ : Odrv4
    port map (
            O => \N__57375\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8\
        );

    \I__12016\ : Odrv12
    port map (
            O => \N__57372\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8\
        );

    \I__12015\ : CascadeMux
    port map (
            O => \N__57367\,
            I => \N__57364\
        );

    \I__12014\ : InMux
    port map (
            O => \N__57364\,
            I => \N__57361\
        );

    \I__12013\ : LocalMux
    port map (
            O => \N__57361\,
            I => \N__57358\
        );

    \I__12012\ : Span4Mux_v
    port map (
            O => \N__57358\,
            I => \N__57355\
        );

    \I__12011\ : Odrv4
    port map (
            O => \N__57355\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_12\
        );

    \I__12010\ : InMux
    port map (
            O => \N__57352\,
            I => \bfn_21_24_0_\
        );

    \I__12009\ : InMux
    port map (
            O => \N__57349\,
            I => \N__57346\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__57346\,
            I => \N__57343\
        );

    \I__12007\ : Odrv12
    port map (
            O => \N__57343\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_13\
        );

    \I__12006\ : CascadeMux
    port map (
            O => \N__57340\,
            I => \N__57337\
        );

    \I__12005\ : InMux
    port map (
            O => \N__57337\,
            I => \N__57334\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__57334\,
            I => \N__57330\
        );

    \I__12003\ : InMux
    port map (
            O => \N__57333\,
            I => \N__57327\
        );

    \I__12002\ : Span4Mux_v
    port map (
            O => \N__57330\,
            I => \N__57324\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__57327\,
            I => \N__57321\
        );

    \I__12000\ : Odrv4
    port map (
            O => \N__57324\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9\
        );

    \I__11999\ : Odrv4
    port map (
            O => \N__57321\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9\
        );

    \I__11998\ : InMux
    port map (
            O => \N__57316\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15921\
        );

    \I__11997\ : InMux
    port map (
            O => \N__57313\,
            I => \N__57310\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__57310\,
            I => \N__57307\
        );

    \I__11995\ : Odrv4
    port map (
            O => \N__57307\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_14\
        );

    \I__11994\ : CascadeMux
    port map (
            O => \N__57304\,
            I => \N__57301\
        );

    \I__11993\ : InMux
    port map (
            O => \N__57301\,
            I => \N__57298\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__57298\,
            I => \N__57294\
        );

    \I__11991\ : InMux
    port map (
            O => \N__57297\,
            I => \N__57291\
        );

    \I__11990\ : Span4Mux_v
    port map (
            O => \N__57294\,
            I => \N__57288\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__57291\,
            I => \N__57285\
        );

    \I__11988\ : Odrv4
    port map (
            O => \N__57288\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10\
        );

    \I__11987\ : Odrv4
    port map (
            O => \N__57285\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10\
        );

    \I__11986\ : InMux
    port map (
            O => \N__57280\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15922\
        );

    \I__11985\ : InMux
    port map (
            O => \N__57277\,
            I => \N__57273\
        );

    \I__11984\ : CascadeMux
    port map (
            O => \N__57276\,
            I => \N__57270\
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__57273\,
            I => \N__57267\
        );

    \I__11982\ : InMux
    port map (
            O => \N__57270\,
            I => \N__57264\
        );

    \I__11981\ : Span4Mux_v
    port map (
            O => \N__57267\,
            I => \N__57261\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__57264\,
            I => \N__57258\
        );

    \I__11979\ : Odrv4
    port map (
            O => \N__57261\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11\
        );

    \I__11978\ : Odrv4
    port map (
            O => \N__57258\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11\
        );

    \I__11977\ : CascadeMux
    port map (
            O => \N__57253\,
            I => \N__57250\
        );

    \I__11976\ : InMux
    port map (
            O => \N__57250\,
            I => \N__57247\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__57247\,
            I => \N__57244\
        );

    \I__11974\ : Span4Mux_h
    port map (
            O => \N__57244\,
            I => \N__57241\
        );

    \I__11973\ : Odrv4
    port map (
            O => \N__57241\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_15\
        );

    \I__11972\ : InMux
    port map (
            O => \N__57238\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15923\
        );

    \I__11971\ : InMux
    port map (
            O => \N__57235\,
            I => \N__57232\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__57232\,
            I => \N__57229\
        );

    \I__11969\ : Span4Mux_v
    port map (
            O => \N__57229\,
            I => \N__57226\
        );

    \I__11968\ : Odrv4
    port map (
            O => \N__57226\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_16\
        );

    \I__11967\ : CascadeMux
    port map (
            O => \N__57223\,
            I => \N__57220\
        );

    \I__11966\ : InMux
    port map (
            O => \N__57220\,
            I => \N__57216\
        );

    \I__11965\ : InMux
    port map (
            O => \N__57219\,
            I => \N__57213\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__57216\,
            I => \N__57210\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__57213\,
            I => \N__57207\
        );

    \I__11962\ : Odrv4
    port map (
            O => \N__57210\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12\
        );

    \I__11961\ : Odrv12
    port map (
            O => \N__57207\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12\
        );

    \I__11960\ : InMux
    port map (
            O => \N__57202\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15924\
        );

    \I__11959\ : InMux
    port map (
            O => \N__57199\,
            I => \N__57196\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__57196\,
            I => \N__57192\
        );

    \I__11957\ : InMux
    port map (
            O => \N__57195\,
            I => \N__57189\
        );

    \I__11956\ : Span12Mux_s10_v
    port map (
            O => \N__57192\,
            I => \N__57186\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__57189\,
            I => \N__57183\
        );

    \I__11954\ : Odrv12
    port map (
            O => \N__57186\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13\
        );

    \I__11953\ : Odrv12
    port map (
            O => \N__57183\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13\
        );

    \I__11952\ : CascadeMux
    port map (
            O => \N__57178\,
            I => \N__57175\
        );

    \I__11951\ : InMux
    port map (
            O => \N__57175\,
            I => \N__57172\
        );

    \I__11950\ : LocalMux
    port map (
            O => \N__57172\,
            I => \N__57169\
        );

    \I__11949\ : Span4Mux_h
    port map (
            O => \N__57169\,
            I => \N__57166\
        );

    \I__11948\ : Odrv4
    port map (
            O => \N__57166\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_17\
        );

    \I__11947\ : InMux
    port map (
            O => \N__57163\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15925\
        );

    \I__11946\ : InMux
    port map (
            O => \N__57160\,
            I => \N__57157\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__57157\,
            I => \N__57154\
        );

    \I__11944\ : Span4Mux_h
    port map (
            O => \N__57154\,
            I => \N__57150\
        );

    \I__11943\ : InMux
    port map (
            O => \N__57153\,
            I => \N__57147\
        );

    \I__11942\ : Span4Mux_v
    port map (
            O => \N__57150\,
            I => \N__57144\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__57147\,
            I => \N__57141\
        );

    \I__11940\ : Odrv4
    port map (
            O => \N__57144\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14\
        );

    \I__11939\ : Odrv4
    port map (
            O => \N__57141\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14\
        );

    \I__11938\ : CascadeMux
    port map (
            O => \N__57136\,
            I => \N__57133\
        );

    \I__11937\ : InMux
    port map (
            O => \N__57133\,
            I => \N__57130\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__57130\,
            I => \N__57127\
        );

    \I__11935\ : Span4Mux_h
    port map (
            O => \N__57127\,
            I => \N__57124\
        );

    \I__11934\ : Odrv4
    port map (
            O => \N__57124\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_18\
        );

    \I__11933\ : InMux
    port map (
            O => \N__57121\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15926\
        );

    \I__11932\ : InMux
    port map (
            O => \N__57118\,
            I => \N__57115\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__57115\,
            I => \N__57111\
        );

    \I__11930\ : InMux
    port map (
            O => \N__57114\,
            I => \N__57108\
        );

    \I__11929\ : Span4Mux_h
    port map (
            O => \N__57111\,
            I => \N__57103\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__57108\,
            I => \N__57103\
        );

    \I__11927\ : Span4Mux_v
    port map (
            O => \N__57103\,
            I => \N__57100\
        );

    \I__11926\ : Odrv4
    port map (
            O => \N__57100\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_15\
        );

    \I__11925\ : CascadeMux
    port map (
            O => \N__57097\,
            I => \N__57094\
        );

    \I__11924\ : InMux
    port map (
            O => \N__57094\,
            I => \N__57091\
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__57091\,
            I => \N__57088\
        );

    \I__11922\ : Span4Mux_h
    port map (
            O => \N__57088\,
            I => \N__57085\
        );

    \I__11921\ : Odrv4
    port map (
            O => \N__57085\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_19\
        );

    \I__11920\ : InMux
    port map (
            O => \N__57082\,
            I => \N__57079\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__57079\,
            I => \N__57076\
        );

    \I__11918\ : Odrv12
    port map (
            O => \N__57076\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_0\
        );

    \I__11917\ : CascadeMux
    port map (
            O => \N__57073\,
            I => \N__57070\
        );

    \I__11916\ : InMux
    port map (
            O => \N__57070\,
            I => \N__57067\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__57067\,
            I => \N__57064\
        );

    \I__11914\ : Odrv4
    port map (
            O => \N__57064\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_4\
        );

    \I__11913\ : InMux
    port map (
            O => \N__57061\,
            I => \N__57058\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__57058\,
            I => \N__57055\
        );

    \I__11911\ : Odrv12
    port map (
            O => \N__57055\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_5\
        );

    \I__11910\ : CascadeMux
    port map (
            O => \N__57052\,
            I => \N__57049\
        );

    \I__11909\ : InMux
    port map (
            O => \N__57049\,
            I => \N__57046\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__57046\,
            I => \N__57043\
        );

    \I__11907\ : Odrv12
    port map (
            O => \N__57043\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_1\
        );

    \I__11906\ : InMux
    port map (
            O => \N__57040\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15913\
        );

    \I__11905\ : InMux
    port map (
            O => \N__57037\,
            I => \N__57034\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__57034\,
            I => \N__57031\
        );

    \I__11903\ : Odrv4
    port map (
            O => \N__57031\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_2\
        );

    \I__11902\ : CascadeMux
    port map (
            O => \N__57028\,
            I => \N__57025\
        );

    \I__11901\ : InMux
    port map (
            O => \N__57025\,
            I => \N__57022\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__57022\,
            I => \N__57019\
        );

    \I__11899\ : Span4Mux_v
    port map (
            O => \N__57019\,
            I => \N__57016\
        );

    \I__11898\ : Odrv4
    port map (
            O => \N__57016\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_6\
        );

    \I__11897\ : InMux
    port map (
            O => \N__57013\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15914\
        );

    \I__11896\ : InMux
    port map (
            O => \N__57010\,
            I => \N__57007\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__57007\,
            I => \N__57004\
        );

    \I__11894\ : Odrv12
    port map (
            O => \N__57004\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_3\
        );

    \I__11893\ : CascadeMux
    port map (
            O => \N__57001\,
            I => \N__56998\
        );

    \I__11892\ : InMux
    port map (
            O => \N__56998\,
            I => \N__56995\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__56995\,
            I => \N__56992\
        );

    \I__11890\ : Odrv12
    port map (
            O => \N__56992\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_7\
        );

    \I__11889\ : InMux
    port map (
            O => \N__56989\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15915\
        );

    \I__11888\ : InMux
    port map (
            O => \N__56986\,
            I => \N__56983\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__56983\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_4\
        );

    \I__11886\ : CascadeMux
    port map (
            O => \N__56980\,
            I => \N__56977\
        );

    \I__11885\ : InMux
    port map (
            O => \N__56977\,
            I => \N__56974\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__56974\,
            I => \N__56971\
        );

    \I__11883\ : Odrv4
    port map (
            O => \N__56971\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_8\
        );

    \I__11882\ : InMux
    port map (
            O => \N__56968\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15916\
        );

    \I__11881\ : InMux
    port map (
            O => \N__56965\,
            I => \N__56962\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__56962\,
            I => \N__56959\
        );

    \I__11879\ : Odrv12
    port map (
            O => \N__56959\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_5\
        );

    \I__11878\ : CascadeMux
    port map (
            O => \N__56956\,
            I => \N__56953\
        );

    \I__11877\ : InMux
    port map (
            O => \N__56953\,
            I => \N__56950\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__56950\,
            I => \N__56947\
        );

    \I__11875\ : Odrv4
    port map (
            O => \N__56947\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_9\
        );

    \I__11874\ : InMux
    port map (
            O => \N__56944\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15917\
        );

    \I__11873\ : InMux
    port map (
            O => \N__56941\,
            I => \N__56938\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__56938\,
            I => \N__56935\
        );

    \I__11871\ : Odrv4
    port map (
            O => \N__56935\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_6\
        );

    \I__11870\ : CascadeMux
    port map (
            O => \N__56932\,
            I => \N__56929\
        );

    \I__11869\ : InMux
    port map (
            O => \N__56929\,
            I => \N__56926\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__56926\,
            I => \N__56923\
        );

    \I__11867\ : Odrv4
    port map (
            O => \N__56923\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_10\
        );

    \I__11866\ : InMux
    port map (
            O => \N__56920\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15918\
        );

    \I__11865\ : InMux
    port map (
            O => \N__56917\,
            I => \N__56914\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__56914\,
            I => \N__56910\
        );

    \I__11863\ : InMux
    port map (
            O => \N__56913\,
            I => \N__56907\
        );

    \I__11862\ : Span4Mux_v
    port map (
            O => \N__56910\,
            I => \N__56904\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__56907\,
            I => \N__56901\
        );

    \I__11860\ : Odrv4
    port map (
            O => \N__56904\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0\
        );

    \I__11859\ : Odrv4
    port map (
            O => \N__56901\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0\
        );

    \I__11858\ : CascadeMux
    port map (
            O => \N__56896\,
            I => \N__56893\
        );

    \I__11857\ : InMux
    port map (
            O => \N__56893\,
            I => \N__56890\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__56890\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_11\
        );

    \I__11855\ : InMux
    port map (
            O => \N__56887\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15919\
        );

    \I__11854\ : InMux
    port map (
            O => \N__56884\,
            I => \N__56881\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__56881\,
            I => \N__56878\
        );

    \I__11852\ : Span4Mux_h
    port map (
            O => \N__56878\,
            I => \N__56875\
        );

    \I__11851\ : Odrv4
    port map (
            O => \N__56875\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n400\
        );

    \I__11850\ : InMux
    port map (
            O => \N__56872\,
            I => \bfn_21_22_0_\
        );

    \I__11849\ : InMux
    port map (
            O => \N__56869\,
            I => \N__56866\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__56866\,
            I => \N__56863\
        );

    \I__11847\ : Span4Mux_h
    port map (
            O => \N__56863\,
            I => \N__56860\
        );

    \I__11846\ : Odrv4
    port map (
            O => \N__56860\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n449\
        );

    \I__11845\ : InMux
    port map (
            O => \N__56857\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18182\
        );

    \I__11844\ : InMux
    port map (
            O => \N__56854\,
            I => \N__56851\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__56851\,
            I => \N__56848\
        );

    \I__11842\ : Span12Mux_h
    port map (
            O => \N__56848\,
            I => \N__56845\
        );

    \I__11841\ : Odrv12
    port map (
            O => \N__56845\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n498\
        );

    \I__11840\ : InMux
    port map (
            O => \N__56842\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18183\
        );

    \I__11839\ : InMux
    port map (
            O => \N__56839\,
            I => \N__56836\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__56836\,
            I => \N__56833\
        );

    \I__11837\ : Span4Mux_h
    port map (
            O => \N__56833\,
            I => \N__56830\
        );

    \I__11836\ : Odrv4
    port map (
            O => \N__56830\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n547\
        );

    \I__11835\ : InMux
    port map (
            O => \N__56827\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18184\
        );

    \I__11834\ : InMux
    port map (
            O => \N__56824\,
            I => \N__56814\
        );

    \I__11833\ : InMux
    port map (
            O => \N__56823\,
            I => \N__56794\
        );

    \I__11832\ : InMux
    port map (
            O => \N__56822\,
            I => \N__56794\
        );

    \I__11831\ : InMux
    port map (
            O => \N__56821\,
            I => \N__56794\
        );

    \I__11830\ : InMux
    port map (
            O => \N__56820\,
            I => \N__56785\
        );

    \I__11829\ : InMux
    port map (
            O => \N__56819\,
            I => \N__56785\
        );

    \I__11828\ : InMux
    port map (
            O => \N__56818\,
            I => \N__56785\
        );

    \I__11827\ : InMux
    port map (
            O => \N__56817\,
            I => \N__56785\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__56814\,
            I => \N__56775\
        );

    \I__11825\ : InMux
    port map (
            O => \N__56813\,
            I => \N__56766\
        );

    \I__11824\ : InMux
    port map (
            O => \N__56812\,
            I => \N__56766\
        );

    \I__11823\ : InMux
    port map (
            O => \N__56811\,
            I => \N__56766\
        );

    \I__11822\ : InMux
    port map (
            O => \N__56810\,
            I => \N__56766\
        );

    \I__11821\ : InMux
    port map (
            O => \N__56809\,
            I => \N__56757\
        );

    \I__11820\ : InMux
    port map (
            O => \N__56808\,
            I => \N__56757\
        );

    \I__11819\ : InMux
    port map (
            O => \N__56807\,
            I => \N__56757\
        );

    \I__11818\ : InMux
    port map (
            O => \N__56806\,
            I => \N__56757\
        );

    \I__11817\ : InMux
    port map (
            O => \N__56805\,
            I => \N__56752\
        );

    \I__11816\ : InMux
    port map (
            O => \N__56804\,
            I => \N__56752\
        );

    \I__11815\ : InMux
    port map (
            O => \N__56803\,
            I => \N__56745\
        );

    \I__11814\ : InMux
    port map (
            O => \N__56802\,
            I => \N__56745\
        );

    \I__11813\ : InMux
    port map (
            O => \N__56801\,
            I => \N__56745\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__56794\,
            I => \N__56740\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__56785\,
            I => \N__56740\
        );

    \I__11810\ : InMux
    port map (
            O => \N__56784\,
            I => \N__56733\
        );

    \I__11809\ : InMux
    port map (
            O => \N__56783\,
            I => \N__56733\
        );

    \I__11808\ : InMux
    port map (
            O => \N__56782\,
            I => \N__56733\
        );

    \I__11807\ : InMux
    port map (
            O => \N__56781\,
            I => \N__56724\
        );

    \I__11806\ : InMux
    port map (
            O => \N__56780\,
            I => \N__56724\
        );

    \I__11805\ : InMux
    port map (
            O => \N__56779\,
            I => \N__56724\
        );

    \I__11804\ : InMux
    port map (
            O => \N__56778\,
            I => \N__56724\
        );

    \I__11803\ : Odrv4
    port map (
            O => \N__56775\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11802\ : LocalMux
    port map (
            O => \N__56766\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__56757\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__56752\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__56745\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11798\ : Odrv12
    port map (
            O => \N__56740\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__56733\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__56724\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11795\ : InMux
    port map (
            O => \N__56707\,
            I => \N__56704\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__56704\,
            I => \N__56701\
        );

    \I__11793\ : Span4Mux_h
    port map (
            O => \N__56701\,
            I => \N__56698\
        );

    \I__11792\ : Odrv4
    port map (
            O => \N__56698\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n596\
        );

    \I__11791\ : InMux
    port map (
            O => \N__56695\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18185\
        );

    \I__11790\ : CascadeMux
    port map (
            O => \N__56692\,
            I => \N__56689\
        );

    \I__11789\ : InMux
    port map (
            O => \N__56689\,
            I => \N__56686\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__56686\,
            I => \N__56683\
        );

    \I__11787\ : Span4Mux_v
    port map (
            O => \N__56683\,
            I => \N__56680\
        );

    \I__11786\ : Odrv4
    port map (
            O => \N__56680\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n645\
        );

    \I__11785\ : InMux
    port map (
            O => \N__56677\,
            I => \N__56671\
        );

    \I__11784\ : InMux
    port map (
            O => \N__56676\,
            I => \N__56671\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__56671\,
            I => \N__56668\
        );

    \I__11782\ : Span4Mux_v
    port map (
            O => \N__56668\,
            I => \N__56665\
        );

    \I__11781\ : Odrv4
    port map (
            O => \N__56665\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n691\
        );

    \I__11780\ : InMux
    port map (
            O => \N__56662\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18186\
        );

    \I__11779\ : InMux
    port map (
            O => \N__56659\,
            I => \N__56656\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__56656\,
            I => \N__56653\
        );

    \I__11777\ : Span4Mux_v
    port map (
            O => \N__56653\,
            I => \N__56650\
        );

    \I__11776\ : Odrv4
    port map (
            O => \N__56650\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n694\
        );

    \I__11775\ : CascadeMux
    port map (
            O => \N__56647\,
            I => \N__56644\
        );

    \I__11774\ : InMux
    port map (
            O => \N__56644\,
            I => \N__56641\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__56641\,
            I => \N__56638\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__56638\,
            I => \N__56635\
        );

    \I__11771\ : Odrv4
    port map (
            O => \N__56635\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n742\
        );

    \I__11770\ : InMux
    port map (
            O => \N__56632\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18187\
        );

    \I__11769\ : InMux
    port map (
            O => \N__56629\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743\
        );

    \I__11768\ : CascadeMux
    port map (
            O => \N__56626\,
            I => \N__56623\
        );

    \I__11767\ : InMux
    port map (
            O => \N__56623\,
            I => \N__56620\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__56620\,
            I => \N__56617\
        );

    \I__11765\ : Span4Mux_h
    port map (
            O => \N__56617\,
            I => \N__56614\
        );

    \I__11764\ : Odrv4
    port map (
            O => \N__56614\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_CO\
        );

    \I__11763\ : CascadeMux
    port map (
            O => \N__56611\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20640_cascade_\
        );

    \I__11762\ : InMux
    port map (
            O => \N__56608\,
            I => \N__56605\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__56605\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19308\
        );

    \I__11760\ : InMux
    port map (
            O => \N__56602\,
            I => \N__56599\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__56599\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n57\
        );

    \I__11758\ : InMux
    port map (
            O => \N__56596\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18174\
        );

    \I__11757\ : CascadeMux
    port map (
            O => \N__56593\,
            I => \N__56590\
        );

    \I__11756\ : InMux
    port map (
            O => \N__56590\,
            I => \N__56587\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__56587\,
            I => \N__56584\
        );

    \I__11754\ : Span4Mux_v
    port map (
            O => \N__56584\,
            I => \N__56581\
        );

    \I__11753\ : Span4Mux_v
    port map (
            O => \N__56581\,
            I => \N__56578\
        );

    \I__11752\ : Odrv4
    port map (
            O => \N__56578\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n106\
        );

    \I__11751\ : InMux
    port map (
            O => \N__56575\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18175\
        );

    \I__11750\ : InMux
    port map (
            O => \N__56572\,
            I => \N__56569\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__56569\,
            I => \N__56566\
        );

    \I__11748\ : Span4Mux_h
    port map (
            O => \N__56566\,
            I => \N__56563\
        );

    \I__11747\ : Odrv4
    port map (
            O => \N__56563\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n155\
        );

    \I__11746\ : InMux
    port map (
            O => \N__56560\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18176\
        );

    \I__11745\ : InMux
    port map (
            O => \N__56557\,
            I => \N__56554\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__56554\,
            I => \N__56551\
        );

    \I__11743\ : Span4Mux_v
    port map (
            O => \N__56551\,
            I => \N__56548\
        );

    \I__11742\ : Odrv4
    port map (
            O => \N__56548\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n204\
        );

    \I__11741\ : InMux
    port map (
            O => \N__56545\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18177\
        );

    \I__11740\ : InMux
    port map (
            O => \N__56542\,
            I => \N__56539\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__56539\,
            I => \N__56536\
        );

    \I__11738\ : Span4Mux_v
    port map (
            O => \N__56536\,
            I => \N__56533\
        );

    \I__11737\ : Odrv4
    port map (
            O => \N__56533\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n253\
        );

    \I__11736\ : InMux
    port map (
            O => \N__56530\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18178\
        );

    \I__11735\ : InMux
    port map (
            O => \N__56527\,
            I => \N__56524\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__56524\,
            I => \N__56521\
        );

    \I__11733\ : Span4Mux_v
    port map (
            O => \N__56521\,
            I => \N__56518\
        );

    \I__11732\ : Sp12to4
    port map (
            O => \N__56518\,
            I => \N__56515\
        );

    \I__11731\ : Odrv12
    port map (
            O => \N__56515\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n302\
        );

    \I__11730\ : InMux
    port map (
            O => \N__56512\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18179\
        );

    \I__11729\ : InMux
    port map (
            O => \N__56509\,
            I => \N__56506\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__56506\,
            I => \N__56503\
        );

    \I__11727\ : Span4Mux_h
    port map (
            O => \N__56503\,
            I => \N__56500\
        );

    \I__11726\ : Odrv4
    port map (
            O => \N__56500\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n351\
        );

    \I__11725\ : InMux
    port map (
            O => \N__56497\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18180\
        );

    \I__11724\ : InMux
    port map (
            O => \N__56494\,
            I => \N__56485\
        );

    \I__11723\ : InMux
    port map (
            O => \N__56493\,
            I => \N__56485\
        );

    \I__11722\ : InMux
    port map (
            O => \N__56492\,
            I => \N__56485\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__56485\,
            I => \N__56473\
        );

    \I__11720\ : InMux
    port map (
            O => \N__56484\,
            I => \N__56464\
        );

    \I__11719\ : InMux
    port map (
            O => \N__56483\,
            I => \N__56464\
        );

    \I__11718\ : InMux
    port map (
            O => \N__56482\,
            I => \N__56464\
        );

    \I__11717\ : InMux
    port map (
            O => \N__56481\,
            I => \N__56464\
        );

    \I__11716\ : CascadeMux
    port map (
            O => \N__56480\,
            I => \N__56451\
        );

    \I__11715\ : CascadeMux
    port map (
            O => \N__56479\,
            I => \N__56444\
        );

    \I__11714\ : InMux
    port map (
            O => \N__56478\,
            I => \N__56433\
        );

    \I__11713\ : InMux
    port map (
            O => \N__56477\,
            I => \N__56433\
        );

    \I__11712\ : InMux
    port map (
            O => \N__56476\,
            I => \N__56433\
        );

    \I__11711\ : Span4Mux_v
    port map (
            O => \N__56473\,
            I => \N__56428\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__56464\,
            I => \N__56428\
        );

    \I__11709\ : InMux
    port map (
            O => \N__56463\,
            I => \N__56425\
        );

    \I__11708\ : InMux
    port map (
            O => \N__56462\,
            I => \N__56412\
        );

    \I__11707\ : InMux
    port map (
            O => \N__56461\,
            I => \N__56412\
        );

    \I__11706\ : InMux
    port map (
            O => \N__56460\,
            I => \N__56412\
        );

    \I__11705\ : InMux
    port map (
            O => \N__56459\,
            I => \N__56412\
        );

    \I__11704\ : InMux
    port map (
            O => \N__56458\,
            I => \N__56412\
        );

    \I__11703\ : InMux
    port map (
            O => \N__56457\,
            I => \N__56412\
        );

    \I__11702\ : InMux
    port map (
            O => \N__56456\,
            I => \N__56399\
        );

    \I__11701\ : InMux
    port map (
            O => \N__56455\,
            I => \N__56399\
        );

    \I__11700\ : InMux
    port map (
            O => \N__56454\,
            I => \N__56399\
        );

    \I__11699\ : InMux
    port map (
            O => \N__56451\,
            I => \N__56399\
        );

    \I__11698\ : InMux
    port map (
            O => \N__56450\,
            I => \N__56399\
        );

    \I__11697\ : InMux
    port map (
            O => \N__56449\,
            I => \N__56399\
        );

    \I__11696\ : InMux
    port map (
            O => \N__56448\,
            I => \N__56390\
        );

    \I__11695\ : InMux
    port map (
            O => \N__56447\,
            I => \N__56390\
        );

    \I__11694\ : InMux
    port map (
            O => \N__56444\,
            I => \N__56390\
        );

    \I__11693\ : InMux
    port map (
            O => \N__56443\,
            I => \N__56390\
        );

    \I__11692\ : InMux
    port map (
            O => \N__56442\,
            I => \N__56383\
        );

    \I__11691\ : InMux
    port map (
            O => \N__56441\,
            I => \N__56383\
        );

    \I__11690\ : InMux
    port map (
            O => \N__56440\,
            I => \N__56383\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__56433\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11688\ : Odrv4
    port map (
            O => \N__56428\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__56425\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__56412\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__56399\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__56390\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__56383\,
            I => \Saturate_out1_31__N_266_adj_2417\
        );

    \I__11682\ : InMux
    port map (
            O => \N__56368\,
            I => \N__56353\
        );

    \I__11681\ : InMux
    port map (
            O => \N__56367\,
            I => \N__56353\
        );

    \I__11680\ : InMux
    port map (
            O => \N__56366\,
            I => \N__56353\
        );

    \I__11679\ : CascadeMux
    port map (
            O => \N__56365\,
            I => \N__56349\
        );

    \I__11678\ : CascadeMux
    port map (
            O => \N__56364\,
            I => \N__56346\
        );

    \I__11677\ : InMux
    port map (
            O => \N__56363\,
            I => \N__56335\
        );

    \I__11676\ : InMux
    port map (
            O => \N__56362\,
            I => \N__56335\
        );

    \I__11675\ : InMux
    port map (
            O => \N__56361\,
            I => \N__56335\
        );

    \I__11674\ : CascadeMux
    port map (
            O => \N__56360\,
            I => \N__56332\
        );

    \I__11673\ : LocalMux
    port map (
            O => \N__56353\,
            I => \N__56326\
        );

    \I__11672\ : InMux
    port map (
            O => \N__56352\,
            I => \N__56313\
        );

    \I__11671\ : InMux
    port map (
            O => \N__56349\,
            I => \N__56313\
        );

    \I__11670\ : InMux
    port map (
            O => \N__56346\,
            I => \N__56313\
        );

    \I__11669\ : InMux
    port map (
            O => \N__56345\,
            I => \N__56313\
        );

    \I__11668\ : InMux
    port map (
            O => \N__56344\,
            I => \N__56313\
        );

    \I__11667\ : InMux
    port map (
            O => \N__56343\,
            I => \N__56313\
        );

    \I__11666\ : InMux
    port map (
            O => \N__56342\,
            I => \N__56310\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__56335\,
            I => \N__56294\
        );

    \I__11664\ : InMux
    port map (
            O => \N__56332\,
            I => \N__56285\
        );

    \I__11663\ : InMux
    port map (
            O => \N__56331\,
            I => \N__56285\
        );

    \I__11662\ : InMux
    port map (
            O => \N__56330\,
            I => \N__56285\
        );

    \I__11661\ : InMux
    port map (
            O => \N__56329\,
            I => \N__56285\
        );

    \I__11660\ : Span4Mux_v
    port map (
            O => \N__56326\,
            I => \N__56278\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__56313\,
            I => \N__56278\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__56310\,
            I => \N__56278\
        );

    \I__11657\ : InMux
    port map (
            O => \N__56309\,
            I => \N__56269\
        );

    \I__11656\ : InMux
    port map (
            O => \N__56308\,
            I => \N__56269\
        );

    \I__11655\ : InMux
    port map (
            O => \N__56307\,
            I => \N__56269\
        );

    \I__11654\ : InMux
    port map (
            O => \N__56306\,
            I => \N__56269\
        );

    \I__11653\ : InMux
    port map (
            O => \N__56305\,
            I => \N__56260\
        );

    \I__11652\ : InMux
    port map (
            O => \N__56304\,
            I => \N__56260\
        );

    \I__11651\ : InMux
    port map (
            O => \N__56303\,
            I => \N__56260\
        );

    \I__11650\ : InMux
    port map (
            O => \N__56302\,
            I => \N__56260\
        );

    \I__11649\ : InMux
    port map (
            O => \N__56301\,
            I => \N__56251\
        );

    \I__11648\ : InMux
    port map (
            O => \N__56300\,
            I => \N__56251\
        );

    \I__11647\ : InMux
    port map (
            O => \N__56299\,
            I => \N__56251\
        );

    \I__11646\ : InMux
    port map (
            O => \N__56298\,
            I => \N__56251\
        );

    \I__11645\ : InMux
    port map (
            O => \N__56297\,
            I => \N__56248\
        );

    \I__11644\ : Odrv4
    port map (
            O => \N__56294\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__56285\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11642\ : Odrv4
    port map (
            O => \N__56278\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__56269\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__56260\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__56251\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__56248\,
            I => \Saturate_out1_31__N_267_adj_2418\
        );

    \I__11637\ : CascadeMux
    port map (
            O => \N__56233\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20660_cascade_\
        );

    \I__11636\ : CascadeMux
    port map (
            O => \N__56230\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20654_cascade_\
        );

    \I__11635\ : InMux
    port map (
            O => \N__56227\,
            I => \N__56224\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__56224\,
            I => \N__56221\
        );

    \I__11633\ : Span4Mux_v
    port map (
            O => \N__56221\,
            I => \N__56218\
        );

    \I__11632\ : Odrv4
    port map (
            O => \N__56218\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n449_adj_492\
        );

    \I__11631\ : CascadeMux
    port map (
            O => \N__56215\,
            I => \N__56211\
        );

    \I__11630\ : CascadeMux
    port map (
            O => \N__56214\,
            I => \N__56208\
        );

    \I__11629\ : InMux
    port map (
            O => \N__56211\,
            I => \N__56201\
        );

    \I__11628\ : InMux
    port map (
            O => \N__56208\,
            I => \N__56198\
        );

    \I__11627\ : CascadeMux
    port map (
            O => \N__56207\,
            I => \N__56194\
        );

    \I__11626\ : CascadeMux
    port map (
            O => \N__56206\,
            I => \N__56191\
        );

    \I__11625\ : CascadeMux
    port map (
            O => \N__56205\,
            I => \N__56186\
        );

    \I__11624\ : CascadeMux
    port map (
            O => \N__56204\,
            I => \N__56183\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__56201\,
            I => \N__56179\
        );

    \I__11622\ : LocalMux
    port map (
            O => \N__56198\,
            I => \N__56176\
        );

    \I__11621\ : CascadeMux
    port map (
            O => \N__56197\,
            I => \N__56173\
        );

    \I__11620\ : InMux
    port map (
            O => \N__56194\,
            I => \N__56170\
        );

    \I__11619\ : InMux
    port map (
            O => \N__56191\,
            I => \N__56167\
        );

    \I__11618\ : CascadeMux
    port map (
            O => \N__56190\,
            I => \N__56164\
        );

    \I__11617\ : CascadeMux
    port map (
            O => \N__56189\,
            I => \N__56161\
        );

    \I__11616\ : InMux
    port map (
            O => \N__56186\,
            I => \N__56157\
        );

    \I__11615\ : InMux
    port map (
            O => \N__56183\,
            I => \N__56154\
        );

    \I__11614\ : CascadeMux
    port map (
            O => \N__56182\,
            I => \N__56151\
        );

    \I__11613\ : Span4Mux_v
    port map (
            O => \N__56179\,
            I => \N__56142\
        );

    \I__11612\ : Span4Mux_h
    port map (
            O => \N__56176\,
            I => \N__56139\
        );

    \I__11611\ : InMux
    port map (
            O => \N__56173\,
            I => \N__56136\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__56170\,
            I => \N__56131\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__56167\,
            I => \N__56131\
        );

    \I__11608\ : InMux
    port map (
            O => \N__56164\,
            I => \N__56128\
        );

    \I__11607\ : InMux
    port map (
            O => \N__56161\,
            I => \N__56125\
        );

    \I__11606\ : CascadeMux
    port map (
            O => \N__56160\,
            I => \N__56122\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__56157\,
            I => \N__56116\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__56154\,
            I => \N__56116\
        );

    \I__11603\ : InMux
    port map (
            O => \N__56151\,
            I => \N__56113\
        );

    \I__11602\ : CascadeMux
    port map (
            O => \N__56150\,
            I => \N__56110\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__56149\,
            I => \N__56107\
        );

    \I__11600\ : CascadeMux
    port map (
            O => \N__56148\,
            I => \N__56103\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__56147\,
            I => \N__56099\
        );

    \I__11598\ : CascadeMux
    port map (
            O => \N__56146\,
            I => \N__56095\
        );

    \I__11597\ : CascadeMux
    port map (
            O => \N__56145\,
            I => \N__56091\
        );

    \I__11596\ : Span4Mux_v
    port map (
            O => \N__56142\,
            I => \N__56083\
        );

    \I__11595\ : Span4Mux_v
    port map (
            O => \N__56139\,
            I => \N__56083\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__56136\,
            I => \N__56083\
        );

    \I__11593\ : Span4Mux_v
    port map (
            O => \N__56131\,
            I => \N__56076\
        );

    \I__11592\ : LocalMux
    port map (
            O => \N__56128\,
            I => \N__56076\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__56125\,
            I => \N__56076\
        );

    \I__11590\ : InMux
    port map (
            O => \N__56122\,
            I => \N__56073\
        );

    \I__11589\ : InMux
    port map (
            O => \N__56121\,
            I => \N__56070\
        );

    \I__11588\ : Span4Mux_v
    port map (
            O => \N__56116\,
            I => \N__56065\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__56113\,
            I => \N__56065\
        );

    \I__11586\ : InMux
    port map (
            O => \N__56110\,
            I => \N__56062\
        );

    \I__11585\ : InMux
    port map (
            O => \N__56107\,
            I => \N__56059\
        );

    \I__11584\ : InMux
    port map (
            O => \N__56106\,
            I => \N__56042\
        );

    \I__11583\ : InMux
    port map (
            O => \N__56103\,
            I => \N__56042\
        );

    \I__11582\ : InMux
    port map (
            O => \N__56102\,
            I => \N__56042\
        );

    \I__11581\ : InMux
    port map (
            O => \N__56099\,
            I => \N__56042\
        );

    \I__11580\ : InMux
    port map (
            O => \N__56098\,
            I => \N__56042\
        );

    \I__11579\ : InMux
    port map (
            O => \N__56095\,
            I => \N__56042\
        );

    \I__11578\ : InMux
    port map (
            O => \N__56094\,
            I => \N__56042\
        );

    \I__11577\ : InMux
    port map (
            O => \N__56091\,
            I => \N__56042\
        );

    \I__11576\ : CascadeMux
    port map (
            O => \N__56090\,
            I => \N__56039\
        );

    \I__11575\ : Span4Mux_h
    port map (
            O => \N__56083\,
            I => \N__56035\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__56076\,
            I => \N__56030\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__56073\,
            I => \N__56030\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__56070\,
            I => \N__56027\
        );

    \I__11571\ : Span4Mux_v
    port map (
            O => \N__56065\,
            I => \N__56020\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__56062\,
            I => \N__56020\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__56059\,
            I => \N__56020\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__56042\,
            I => \N__56017\
        );

    \I__11567\ : InMux
    port map (
            O => \N__56039\,
            I => \N__56014\
        );

    \I__11566\ : CascadeMux
    port map (
            O => \N__56038\,
            I => \N__56010\
        );

    \I__11565\ : Span4Mux_v
    port map (
            O => \N__56035\,
            I => \N__56007\
        );

    \I__11564\ : Span4Mux_v
    port map (
            O => \N__56030\,
            I => \N__56004\
        );

    \I__11563\ : Span4Mux_h
    port map (
            O => \N__56027\,
            I => \N__55995\
        );

    \I__11562\ : Span4Mux_v
    port map (
            O => \N__56020\,
            I => \N__55995\
        );

    \I__11561\ : Span4Mux_v
    port map (
            O => \N__56017\,
            I => \N__55995\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__56014\,
            I => \N__55995\
        );

    \I__11559\ : InMux
    port map (
            O => \N__56013\,
            I => \N__55990\
        );

    \I__11558\ : InMux
    port map (
            O => \N__56010\,
            I => \N__55990\
        );

    \I__11557\ : Odrv4
    port map (
            O => \N__56007\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n129\
        );

    \I__11556\ : Odrv4
    port map (
            O => \N__56004\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n129\
        );

    \I__11555\ : Odrv4
    port map (
            O => \N__55995\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n129\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__55990\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n129\
        );

    \I__11553\ : InMux
    port map (
            O => \N__55981\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17744\
        );

    \I__11552\ : InMux
    port map (
            O => \N__55978\,
            I => \N__55975\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__55975\,
            I => \N__55972\
        );

    \I__11550\ : Span4Mux_v
    port map (
            O => \N__55972\,
            I => \N__55969\
        );

    \I__11549\ : Odrv4
    port map (
            O => \N__55969\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n498_adj_469\
        );

    \I__11548\ : CascadeMux
    port map (
            O => \N__55966\,
            I => \N__55961\
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__55965\,
            I => \N__55957\
        );

    \I__11546\ : CascadeMux
    port map (
            O => \N__55964\,
            I => \N__55953\
        );

    \I__11545\ : InMux
    port map (
            O => \N__55961\,
            I => \N__55950\
        );

    \I__11544\ : InMux
    port map (
            O => \N__55960\,
            I => \N__55947\
        );

    \I__11543\ : InMux
    port map (
            O => \N__55957\,
            I => \N__55941\
        );

    \I__11542\ : CascadeMux
    port map (
            O => \N__55956\,
            I => \N__55936\
        );

    \I__11541\ : InMux
    port map (
            O => \N__55953\,
            I => \N__55933\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__55950\,
            I => \N__55928\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__55947\,
            I => \N__55928\
        );

    \I__11538\ : CascadeMux
    port map (
            O => \N__55946\,
            I => \N__55925\
        );

    \I__11537\ : CascadeMux
    port map (
            O => \N__55945\,
            I => \N__55922\
        );

    \I__11536\ : CascadeMux
    port map (
            O => \N__55944\,
            I => \N__55919\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__55941\,
            I => \N__55912\
        );

    \I__11534\ : CascadeMux
    port map (
            O => \N__55940\,
            I => \N__55909\
        );

    \I__11533\ : CascadeMux
    port map (
            O => \N__55939\,
            I => \N__55906\
        );

    \I__11532\ : InMux
    port map (
            O => \N__55936\,
            I => \N__55903\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__55933\,
            I => \N__55900\
        );

    \I__11530\ : Span4Mux_v
    port map (
            O => \N__55928\,
            I => \N__55897\
        );

    \I__11529\ : InMux
    port map (
            O => \N__55925\,
            I => \N__55894\
        );

    \I__11528\ : InMux
    port map (
            O => \N__55922\,
            I => \N__55891\
        );

    \I__11527\ : InMux
    port map (
            O => \N__55919\,
            I => \N__55888\
        );

    \I__11526\ : CascadeMux
    port map (
            O => \N__55918\,
            I => \N__55885\
        );

    \I__11525\ : CascadeMux
    port map (
            O => \N__55917\,
            I => \N__55882\
        );

    \I__11524\ : CascadeMux
    port map (
            O => \N__55916\,
            I => \N__55879\
        );

    \I__11523\ : CascadeMux
    port map (
            O => \N__55915\,
            I => \N__55876\
        );

    \I__11522\ : Span4Mux_v
    port map (
            O => \N__55912\,
            I => \N__55869\
        );

    \I__11521\ : InMux
    port map (
            O => \N__55909\,
            I => \N__55866\
        );

    \I__11520\ : InMux
    port map (
            O => \N__55906\,
            I => \N__55863\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__55903\,
            I => \N__55860\
        );

    \I__11518\ : Span4Mux_h
    port map (
            O => \N__55900\,
            I => \N__55849\
        );

    \I__11517\ : Span4Mux_h
    port map (
            O => \N__55897\,
            I => \N__55849\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__55894\,
            I => \N__55849\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__55891\,
            I => \N__55849\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__55888\,
            I => \N__55849\
        );

    \I__11513\ : InMux
    port map (
            O => \N__55885\,
            I => \N__55846\
        );

    \I__11512\ : InMux
    port map (
            O => \N__55882\,
            I => \N__55843\
        );

    \I__11511\ : InMux
    port map (
            O => \N__55879\,
            I => \N__55840\
        );

    \I__11510\ : InMux
    port map (
            O => \N__55876\,
            I => \N__55836\
        );

    \I__11509\ : CascadeMux
    port map (
            O => \N__55875\,
            I => \N__55832\
        );

    \I__11508\ : CascadeMux
    port map (
            O => \N__55874\,
            I => \N__55828\
        );

    \I__11507\ : CascadeMux
    port map (
            O => \N__55873\,
            I => \N__55824\
        );

    \I__11506\ : CascadeMux
    port map (
            O => \N__55872\,
            I => \N__55820\
        );

    \I__11505\ : Sp12to4
    port map (
            O => \N__55869\,
            I => \N__55813\
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__55866\,
            I => \N__55813\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__55863\,
            I => \N__55813\
        );

    \I__11502\ : Span4Mux_h
    port map (
            O => \N__55860\,
            I => \N__55806\
        );

    \I__11501\ : Span4Mux_v
    port map (
            O => \N__55849\,
            I => \N__55806\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__55846\,
            I => \N__55806\
        );

    \I__11499\ : LocalMux
    port map (
            O => \N__55843\,
            I => \N__55803\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__55840\,
            I => \N__55800\
        );

    \I__11497\ : InMux
    port map (
            O => \N__55839\,
            I => \N__55797\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__55836\,
            I => \N__55794\
        );

    \I__11495\ : InMux
    port map (
            O => \N__55835\,
            I => \N__55777\
        );

    \I__11494\ : InMux
    port map (
            O => \N__55832\,
            I => \N__55777\
        );

    \I__11493\ : InMux
    port map (
            O => \N__55831\,
            I => \N__55777\
        );

    \I__11492\ : InMux
    port map (
            O => \N__55828\,
            I => \N__55777\
        );

    \I__11491\ : InMux
    port map (
            O => \N__55827\,
            I => \N__55777\
        );

    \I__11490\ : InMux
    port map (
            O => \N__55824\,
            I => \N__55777\
        );

    \I__11489\ : InMux
    port map (
            O => \N__55823\,
            I => \N__55777\
        );

    \I__11488\ : InMux
    port map (
            O => \N__55820\,
            I => \N__55777\
        );

    \I__11487\ : Span12Mux_h
    port map (
            O => \N__55813\,
            I => \N__55774\
        );

    \I__11486\ : Span4Mux_v
    port map (
            O => \N__55806\,
            I => \N__55769\
        );

    \I__11485\ : Span4Mux_h
    port map (
            O => \N__55803\,
            I => \N__55769\
        );

    \I__11484\ : Span4Mux_v
    port map (
            O => \N__55800\,
            I => \N__55760\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__55797\,
            I => \N__55760\
        );

    \I__11482\ : Span4Mux_v
    port map (
            O => \N__55794\,
            I => \N__55760\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__55777\,
            I => \N__55760\
        );

    \I__11480\ : Odrv12
    port map (
            O => \N__55774\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n132\
        );

    \I__11479\ : Odrv4
    port map (
            O => \N__55769\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n132\
        );

    \I__11478\ : Odrv4
    port map (
            O => \N__55760\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n132\
        );

    \I__11477\ : InMux
    port map (
            O => \N__55753\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17745\
        );

    \I__11476\ : InMux
    port map (
            O => \N__55750\,
            I => \N__55747\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__55747\,
            I => \N__55744\
        );

    \I__11474\ : Span4Mux_v
    port map (
            O => \N__55744\,
            I => \N__55741\
        );

    \I__11473\ : Odrv4
    port map (
            O => \N__55741\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n547_adj_454\
        );

    \I__11472\ : CascadeMux
    port map (
            O => \N__55738\,
            I => \N__55733\
        );

    \I__11471\ : CascadeMux
    port map (
            O => \N__55737\,
            I => \N__55730\
        );

    \I__11470\ : CascadeMux
    port map (
            O => \N__55736\,
            I => \N__55726\
        );

    \I__11469\ : InMux
    port map (
            O => \N__55733\,
            I => \N__55719\
        );

    \I__11468\ : InMux
    port map (
            O => \N__55730\,
            I => \N__55714\
        );

    \I__11467\ : CascadeMux
    port map (
            O => \N__55729\,
            I => \N__55711\
        );

    \I__11466\ : InMux
    port map (
            O => \N__55726\,
            I => \N__55708\
        );

    \I__11465\ : CascadeMux
    port map (
            O => \N__55725\,
            I => \N__55705\
        );

    \I__11464\ : CascadeMux
    port map (
            O => \N__55724\,
            I => \N__55702\
        );

    \I__11463\ : CascadeMux
    port map (
            O => \N__55723\,
            I => \N__55699\
        );

    \I__11462\ : CascadeMux
    port map (
            O => \N__55722\,
            I => \N__55694\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__55719\,
            I => \N__55691\
        );

    \I__11460\ : CascadeMux
    port map (
            O => \N__55718\,
            I => \N__55688\
        );

    \I__11459\ : CascadeMux
    port map (
            O => \N__55717\,
            I => \N__55685\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__55714\,
            I => \N__55682\
        );

    \I__11457\ : InMux
    port map (
            O => \N__55711\,
            I => \N__55679\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__55708\,
            I => \N__55676\
        );

    \I__11455\ : InMux
    port map (
            O => \N__55705\,
            I => \N__55673\
        );

    \I__11454\ : InMux
    port map (
            O => \N__55702\,
            I => \N__55670\
        );

    \I__11453\ : InMux
    port map (
            O => \N__55699\,
            I => \N__55667\
        );

    \I__11452\ : CascadeMux
    port map (
            O => \N__55698\,
            I => \N__55664\
        );

    \I__11451\ : CascadeMux
    port map (
            O => \N__55697\,
            I => \N__55660\
        );

    \I__11450\ : InMux
    port map (
            O => \N__55694\,
            I => \N__55656\
        );

    \I__11449\ : Span4Mux_v
    port map (
            O => \N__55691\,
            I => \N__55653\
        );

    \I__11448\ : InMux
    port map (
            O => \N__55688\,
            I => \N__55650\
        );

    \I__11447\ : InMux
    port map (
            O => \N__55685\,
            I => \N__55647\
        );

    \I__11446\ : Span4Mux_v
    port map (
            O => \N__55682\,
            I => \N__55642\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__55679\,
            I => \N__55642\
        );

    \I__11444\ : Span4Mux_v
    port map (
            O => \N__55676\,
            I => \N__55633\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__55673\,
            I => \N__55633\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__55670\,
            I => \N__55633\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__55667\,
            I => \N__55633\
        );

    \I__11440\ : InMux
    port map (
            O => \N__55664\,
            I => \N__55630\
        );

    \I__11439\ : InMux
    port map (
            O => \N__55663\,
            I => \N__55627\
        );

    \I__11438\ : InMux
    port map (
            O => \N__55660\,
            I => \N__55624\
        );

    \I__11437\ : CascadeMux
    port map (
            O => \N__55659\,
            I => \N__55621\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__55656\,
            I => \N__55612\
        );

    \I__11435\ : Span4Mux_v
    port map (
            O => \N__55653\,
            I => \N__55605\
        );

    \I__11434\ : LocalMux
    port map (
            O => \N__55650\,
            I => \N__55605\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__55647\,
            I => \N__55605\
        );

    \I__11432\ : Span4Mux_h
    port map (
            O => \N__55642\,
            I => \N__55598\
        );

    \I__11431\ : Span4Mux_v
    port map (
            O => \N__55633\,
            I => \N__55598\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__55630\,
            I => \N__55598\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__55627\,
            I => \N__55595\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__55624\,
            I => \N__55592\
        );

    \I__11427\ : InMux
    port map (
            O => \N__55621\,
            I => \N__55589\
        );

    \I__11426\ : CascadeMux
    port map (
            O => \N__55620\,
            I => \N__55586\
        );

    \I__11425\ : CascadeMux
    port map (
            O => \N__55619\,
            I => \N__55583\
        );

    \I__11424\ : CascadeMux
    port map (
            O => \N__55618\,
            I => \N__55579\
        );

    \I__11423\ : CascadeMux
    port map (
            O => \N__55617\,
            I => \N__55576\
        );

    \I__11422\ : CascadeMux
    port map (
            O => \N__55616\,
            I => \N__55573\
        );

    \I__11421\ : CascadeMux
    port map (
            O => \N__55615\,
            I => \N__55570\
        );

    \I__11420\ : Span12Mux_h
    port map (
            O => \N__55612\,
            I => \N__55567\
        );

    \I__11419\ : Span4Mux_h
    port map (
            O => \N__55605\,
            I => \N__55564\
        );

    \I__11418\ : Span4Mux_v
    port map (
            O => \N__55598\,
            I => \N__55557\
        );

    \I__11417\ : Span4Mux_v
    port map (
            O => \N__55595\,
            I => \N__55557\
        );

    \I__11416\ : Span4Mux_h
    port map (
            O => \N__55592\,
            I => \N__55557\
        );

    \I__11415\ : LocalMux
    port map (
            O => \N__55589\,
            I => \N__55554\
        );

    \I__11414\ : InMux
    port map (
            O => \N__55586\,
            I => \N__55549\
        );

    \I__11413\ : InMux
    port map (
            O => \N__55583\,
            I => \N__55549\
        );

    \I__11412\ : InMux
    port map (
            O => \N__55582\,
            I => \N__55540\
        );

    \I__11411\ : InMux
    port map (
            O => \N__55579\,
            I => \N__55540\
        );

    \I__11410\ : InMux
    port map (
            O => \N__55576\,
            I => \N__55540\
        );

    \I__11409\ : InMux
    port map (
            O => \N__55573\,
            I => \N__55540\
        );

    \I__11408\ : InMux
    port map (
            O => \N__55570\,
            I => \N__55537\
        );

    \I__11407\ : Odrv12
    port map (
            O => \N__55567\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11406\ : Odrv4
    port map (
            O => \N__55564\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11405\ : Odrv4
    port map (
            O => \N__55557\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11404\ : Odrv4
    port map (
            O => \N__55554\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__55549\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__55540\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__55537\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\
        );

    \I__11400\ : InMux
    port map (
            O => \N__55522\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17746\
        );

    \I__11399\ : CascadeMux
    port map (
            O => \N__55519\,
            I => \N__55516\
        );

    \I__11398\ : InMux
    port map (
            O => \N__55516\,
            I => \N__55513\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__55513\,
            I => \N__55506\
        );

    \I__11396\ : InMux
    port map (
            O => \N__55512\,
            I => \N__55497\
        );

    \I__11395\ : InMux
    port map (
            O => \N__55511\,
            I => \N__55497\
        );

    \I__11394\ : InMux
    port map (
            O => \N__55510\,
            I => \N__55497\
        );

    \I__11393\ : InMux
    port map (
            O => \N__55509\,
            I => \N__55497\
        );

    \I__11392\ : Span4Mux_v
    port map (
            O => \N__55506\,
            I => \N__55481\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__55497\,
            I => \N__55481\
        );

    \I__11390\ : InMux
    port map (
            O => \N__55496\,
            I => \N__55472\
        );

    \I__11389\ : InMux
    port map (
            O => \N__55495\,
            I => \N__55472\
        );

    \I__11388\ : InMux
    port map (
            O => \N__55494\,
            I => \N__55472\
        );

    \I__11387\ : InMux
    port map (
            O => \N__55493\,
            I => \N__55472\
        );

    \I__11386\ : InMux
    port map (
            O => \N__55492\,
            I => \N__55465\
        );

    \I__11385\ : InMux
    port map (
            O => \N__55491\,
            I => \N__55465\
        );

    \I__11384\ : InMux
    port map (
            O => \N__55490\,
            I => \N__55465\
        );

    \I__11383\ : InMux
    port map (
            O => \N__55489\,
            I => \N__55456\
        );

    \I__11382\ : InMux
    port map (
            O => \N__55488\,
            I => \N__55456\
        );

    \I__11381\ : InMux
    port map (
            O => \N__55487\,
            I => \N__55456\
        );

    \I__11380\ : InMux
    port map (
            O => \N__55486\,
            I => \N__55456\
        );

    \I__11379\ : Span4Mux_h
    port map (
            O => \N__55481\,
            I => \N__55435\
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__55472\,
            I => \N__55435\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__55465\,
            I => \N__55435\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__55456\,
            I => \N__55435\
        );

    \I__11375\ : InMux
    port map (
            O => \N__55455\,
            I => \N__55430\
        );

    \I__11374\ : InMux
    port map (
            O => \N__55454\,
            I => \N__55430\
        );

    \I__11373\ : InMux
    port map (
            O => \N__55453\,
            I => \N__55423\
        );

    \I__11372\ : InMux
    port map (
            O => \N__55452\,
            I => \N__55423\
        );

    \I__11371\ : InMux
    port map (
            O => \N__55451\,
            I => \N__55423\
        );

    \I__11370\ : InMux
    port map (
            O => \N__55450\,
            I => \N__55416\
        );

    \I__11369\ : InMux
    port map (
            O => \N__55449\,
            I => \N__55416\
        );

    \I__11368\ : InMux
    port map (
            O => \N__55448\,
            I => \N__55416\
        );

    \I__11367\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55407\
        );

    \I__11366\ : InMux
    port map (
            O => \N__55446\,
            I => \N__55407\
        );

    \I__11365\ : InMux
    port map (
            O => \N__55445\,
            I => \N__55407\
        );

    \I__11364\ : InMux
    port map (
            O => \N__55444\,
            I => \N__55407\
        );

    \I__11363\ : Span4Mux_v
    port map (
            O => \N__55435\,
            I => \N__55404\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__55430\,
            I => \N__55395\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__55423\,
            I => \N__55395\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__55416\,
            I => \N__55395\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__55407\,
            I => \N__55395\
        );

    \I__11358\ : Odrv4
    port map (
            O => \N__55404\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11357\ : Odrv12
    port map (
            O => \N__55395\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201\
        );

    \I__11356\ : InMux
    port map (
            O => \N__55390\,
            I => \N__55387\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__55387\,
            I => \N__55384\
        );

    \I__11354\ : Span4Mux_v
    port map (
            O => \N__55384\,
            I => \N__55381\
        );

    \I__11353\ : Odrv4
    port map (
            O => \N__55381\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n596_adj_434\
        );

    \I__11352\ : CascadeMux
    port map (
            O => \N__55378\,
            I => \N__55374\
        );

    \I__11351\ : CascadeMux
    port map (
            O => \N__55377\,
            I => \N__55371\
        );

    \I__11350\ : InMux
    port map (
            O => \N__55374\,
            I => \N__55367\
        );

    \I__11349\ : InMux
    port map (
            O => \N__55371\,
            I => \N__55360\
        );

    \I__11348\ : InMux
    port map (
            O => \N__55370\,
            I => \N__55357\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__55367\,
            I => \N__55353\
        );

    \I__11346\ : CascadeMux
    port map (
            O => \N__55366\,
            I => \N__55350\
        );

    \I__11345\ : CascadeMux
    port map (
            O => \N__55365\,
            I => \N__55345\
        );

    \I__11344\ : CascadeMux
    port map (
            O => \N__55364\,
            I => \N__55342\
        );

    \I__11343\ : CascadeMux
    port map (
            O => \N__55363\,
            I => \N__55338\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__55360\,
            I => \N__55334\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__55357\,
            I => \N__55331\
        );

    \I__11340\ : CascadeMux
    port map (
            O => \N__55356\,
            I => \N__55328\
        );

    \I__11339\ : Span4Mux_v
    port map (
            O => \N__55353\,
            I => \N__55325\
        );

    \I__11338\ : InMux
    port map (
            O => \N__55350\,
            I => \N__55322\
        );

    \I__11337\ : CascadeMux
    port map (
            O => \N__55349\,
            I => \N__55319\
        );

    \I__11336\ : CascadeMux
    port map (
            O => \N__55348\,
            I => \N__55316\
        );

    \I__11335\ : InMux
    port map (
            O => \N__55345\,
            I => \N__55313\
        );

    \I__11334\ : InMux
    port map (
            O => \N__55342\,
            I => \N__55310\
        );

    \I__11333\ : CascadeMux
    port map (
            O => \N__55341\,
            I => \N__55307\
        );

    \I__11332\ : InMux
    port map (
            O => \N__55338\,
            I => \N__55303\
        );

    \I__11331\ : CascadeMux
    port map (
            O => \N__55337\,
            I => \N__55300\
        );

    \I__11330\ : Span4Mux_v
    port map (
            O => \N__55334\,
            I => \N__55297\
        );

    \I__11329\ : Span4Mux_h
    port map (
            O => \N__55331\,
            I => \N__55294\
        );

    \I__11328\ : InMux
    port map (
            O => \N__55328\,
            I => \N__55291\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__55325\,
            I => \N__55286\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__55322\,
            I => \N__55286\
        );

    \I__11325\ : InMux
    port map (
            O => \N__55319\,
            I => \N__55283\
        );

    \I__11324\ : InMux
    port map (
            O => \N__55316\,
            I => \N__55280\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__55313\,
            I => \N__55275\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__55310\,
            I => \N__55275\
        );

    \I__11321\ : InMux
    port map (
            O => \N__55307\,
            I => \N__55272\
        );

    \I__11320\ : CascadeMux
    port map (
            O => \N__55306\,
            I => \N__55269\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__55303\,
            I => \N__55263\
        );

    \I__11318\ : InMux
    port map (
            O => \N__55300\,
            I => \N__55260\
        );

    \I__11317\ : Span4Mux_v
    port map (
            O => \N__55297\,
            I => \N__55253\
        );

    \I__11316\ : Span4Mux_v
    port map (
            O => \N__55294\,
            I => \N__55253\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__55291\,
            I => \N__55253\
        );

    \I__11314\ : Span4Mux_h
    port map (
            O => \N__55286\,
            I => \N__55242\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__55283\,
            I => \N__55242\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__55280\,
            I => \N__55242\
        );

    \I__11311\ : Span4Mux_h
    port map (
            O => \N__55275\,
            I => \N__55242\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__55272\,
            I => \N__55242\
        );

    \I__11309\ : InMux
    port map (
            O => \N__55269\,
            I => \N__55239\
        );

    \I__11308\ : InMux
    port map (
            O => \N__55268\,
            I => \N__55234\
        );

    \I__11307\ : InMux
    port map (
            O => \N__55267\,
            I => \N__55234\
        );

    \I__11306\ : CascadeMux
    port map (
            O => \N__55266\,
            I => \N__55230\
        );

    \I__11305\ : Span12Mux_h
    port map (
            O => \N__55263\,
            I => \N__55224\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__55260\,
            I => \N__55224\
        );

    \I__11303\ : Span4Mux_h
    port map (
            O => \N__55253\,
            I => \N__55221\
        );

    \I__11302\ : Span4Mux_v
    port map (
            O => \N__55242\,
            I => \N__55216\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__55239\,
            I => \N__55216\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__55234\,
            I => \N__55213\
        );

    \I__11299\ : InMux
    port map (
            O => \N__55233\,
            I => \N__55210\
        );

    \I__11298\ : InMux
    port map (
            O => \N__55230\,
            I => \N__55207\
        );

    \I__11297\ : InMux
    port map (
            O => \N__55229\,
            I => \N__55204\
        );

    \I__11296\ : Odrv12
    port map (
            O => \N__55224\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11295\ : Odrv4
    port map (
            O => \N__55221\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11294\ : Odrv4
    port map (
            O => \N__55216\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11293\ : Odrv4
    port map (
            O => \N__55213\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__55210\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__55207\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__55204\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\
        );

    \I__11289\ : InMux
    port map (
            O => \N__55189\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17747\
        );

    \I__11288\ : InMux
    port map (
            O => \N__55186\,
            I => \N__55183\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__55183\,
            I => \N__55176\
        );

    \I__11286\ : InMux
    port map (
            O => \N__55182\,
            I => \N__55173\
        );

    \I__11285\ : InMux
    port map (
            O => \N__55181\,
            I => \N__55170\
        );

    \I__11284\ : CascadeMux
    port map (
            O => \N__55180\,
            I => \N__55167\
        );

    \I__11283\ : InMux
    port map (
            O => \N__55179\,
            I => \N__55163\
        );

    \I__11282\ : Span4Mux_h
    port map (
            O => \N__55176\,
            I => \N__55156\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__55173\,
            I => \N__55156\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__55170\,
            I => \N__55156\
        );

    \I__11279\ : InMux
    port map (
            O => \N__55167\,
            I => \N__55152\
        );

    \I__11278\ : CascadeMux
    port map (
            O => \N__55166\,
            I => \N__55147\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__55163\,
            I => \N__55144\
        );

    \I__11276\ : Span4Mux_v
    port map (
            O => \N__55156\,
            I => \N__55141\
        );

    \I__11275\ : InMux
    port map (
            O => \N__55155\,
            I => \N__55138\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__55152\,
            I => \N__55135\
        );

    \I__11273\ : InMux
    port map (
            O => \N__55151\,
            I => \N__55132\
        );

    \I__11272\ : InMux
    port map (
            O => \N__55150\,
            I => \N__55129\
        );

    \I__11271\ : InMux
    port map (
            O => \N__55147\,
            I => \N__55126\
        );

    \I__11270\ : Span4Mux_v
    port map (
            O => \N__55144\,
            I => \N__55115\
        );

    \I__11269\ : Span4Mux_h
    port map (
            O => \N__55141\,
            I => \N__55115\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__55138\,
            I => \N__55115\
        );

    \I__11267\ : Span4Mux_h
    port map (
            O => \N__55135\,
            I => \N__55106\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__55132\,
            I => \N__55106\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__55129\,
            I => \N__55106\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__55126\,
            I => \N__55106\
        );

    \I__11263\ : InMux
    port map (
            O => \N__55125\,
            I => \N__55103\
        );

    \I__11262\ : InMux
    port map (
            O => \N__55124\,
            I => \N__55100\
        );

    \I__11261\ : InMux
    port map (
            O => \N__55123\,
            I => \N__55097\
        );

    \I__11260\ : InMux
    port map (
            O => \N__55122\,
            I => \N__55094\
        );

    \I__11259\ : Span4Mux_v
    port map (
            O => \N__55115\,
            I => \N__55090\
        );

    \I__11258\ : Span4Mux_v
    port map (
            O => \N__55106\,
            I => \N__55084\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__55103\,
            I => \N__55084\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__55100\,
            I => \N__55077\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__55097\,
            I => \N__55077\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__55094\,
            I => \N__55077\
        );

    \I__11253\ : InMux
    port map (
            O => \N__55093\,
            I => \N__55074\
        );

    \I__11252\ : Span4Mux_h
    port map (
            O => \N__55090\,
            I => \N__55070\
        );

    \I__11251\ : InMux
    port map (
            O => \N__55089\,
            I => \N__55067\
        );

    \I__11250\ : Span4Mux_v
    port map (
            O => \N__55084\,
            I => \N__55060\
        );

    \I__11249\ : Span4Mux_v
    port map (
            O => \N__55077\,
            I => \N__55060\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__55074\,
            I => \N__55060\
        );

    \I__11247\ : InMux
    port map (
            O => \N__55073\,
            I => \N__55057\
        );

    \I__11246\ : Odrv4
    port map (
            O => \N__55070\,
            I => n141
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__55067\,
            I => n141
        );

    \I__11244\ : Odrv4
    port map (
            O => \N__55060\,
            I => n141
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__55057\,
            I => n141
        );

    \I__11242\ : CascadeMux
    port map (
            O => \N__55048\,
            I => \N__55045\
        );

    \I__11241\ : InMux
    port map (
            O => \N__55045\,
            I => \N__55042\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__55042\,
            I => \N__55039\
        );

    \I__11239\ : Span4Mux_h
    port map (
            O => \N__55039\,
            I => \N__55036\
        );

    \I__11238\ : Odrv4
    port map (
            O => \N__55036\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n645_adj_429\
        );

    \I__11237\ : InMux
    port map (
            O => \N__55033\,
            I => \N__55027\
        );

    \I__11236\ : InMux
    port map (
            O => \N__55032\,
            I => \N__55027\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__55027\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n691\
        );

    \I__11234\ : InMux
    port map (
            O => \N__55024\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17748\
        );

    \I__11233\ : InMux
    port map (
            O => \N__55021\,
            I => \N__55018\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__55018\,
            I => \N__55015\
        );

    \I__11231\ : Span12Mux_v
    port map (
            O => \N__55015\,
            I => \N__55012\
        );

    \I__11230\ : Odrv12
    port map (
            O => \N__55012\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n694_adj_427\
        );

    \I__11229\ : CascadeMux
    port map (
            O => \N__55009\,
            I => \N__55006\
        );

    \I__11228\ : InMux
    port map (
            O => \N__55006\,
            I => \N__55002\
        );

    \I__11227\ : CascadeMux
    port map (
            O => \N__55005\,
            I => \N__54998\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__55002\,
            I => \N__54993\
        );

    \I__11225\ : InMux
    port map (
            O => \N__55001\,
            I => \N__54990\
        );

    \I__11224\ : InMux
    port map (
            O => \N__54998\,
            I => \N__54984\
        );

    \I__11223\ : InMux
    port map (
            O => \N__54997\,
            I => \N__54981\
        );

    \I__11222\ : InMux
    port map (
            O => \N__54996\,
            I => \N__54978\
        );

    \I__11221\ : Span4Mux_v
    port map (
            O => \N__54993\,
            I => \N__54973\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__54990\,
            I => \N__54973\
        );

    \I__11219\ : InMux
    port map (
            O => \N__54989\,
            I => \N__54970\
        );

    \I__11218\ : InMux
    port map (
            O => \N__54988\,
            I => \N__54966\
        );

    \I__11217\ : InMux
    port map (
            O => \N__54987\,
            I => \N__54963\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__54984\,
            I => \N__54960\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__54981\,
            I => \N__54955\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__54978\,
            I => \N__54952\
        );

    \I__11213\ : Span4Mux_v
    port map (
            O => \N__54973\,
            I => \N__54947\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__54970\,
            I => \N__54947\
        );

    \I__11211\ : InMux
    port map (
            O => \N__54969\,
            I => \N__54942\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__54966\,
            I => \N__54935\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__54963\,
            I => \N__54935\
        );

    \I__11208\ : Span4Mux_v
    port map (
            O => \N__54960\,
            I => \N__54932\
        );

    \I__11207\ : InMux
    port map (
            O => \N__54959\,
            I => \N__54929\
        );

    \I__11206\ : InMux
    port map (
            O => \N__54958\,
            I => \N__54926\
        );

    \I__11205\ : Span4Mux_h
    port map (
            O => \N__54955\,
            I => \N__54923\
        );

    \I__11204\ : Span4Mux_h
    port map (
            O => \N__54952\,
            I => \N__54918\
        );

    \I__11203\ : Span4Mux_h
    port map (
            O => \N__54947\,
            I => \N__54918\
        );

    \I__11202\ : InMux
    port map (
            O => \N__54946\,
            I => \N__54915\
        );

    \I__11201\ : CascadeMux
    port map (
            O => \N__54945\,
            I => \N__54911\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__54942\,
            I => \N__54908\
        );

    \I__11199\ : InMux
    port map (
            O => \N__54941\,
            I => \N__54905\
        );

    \I__11198\ : InMux
    port map (
            O => \N__54940\,
            I => \N__54902\
        );

    \I__11197\ : Span4Mux_v
    port map (
            O => \N__54935\,
            I => \N__54895\
        );

    \I__11196\ : Span4Mux_h
    port map (
            O => \N__54932\,
            I => \N__54895\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__54929\,
            I => \N__54895\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__54926\,
            I => \N__54886\
        );

    \I__11193\ : Sp12to4
    port map (
            O => \N__54923\,
            I => \N__54886\
        );

    \I__11192\ : Sp12to4
    port map (
            O => \N__54918\,
            I => \N__54886\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__54915\,
            I => \N__54886\
        );

    \I__11190\ : InMux
    port map (
            O => \N__54914\,
            I => \N__54883\
        );

    \I__11189\ : InMux
    port map (
            O => \N__54911\,
            I => \N__54880\
        );

    \I__11188\ : Span4Mux_v
    port map (
            O => \N__54908\,
            I => \N__54873\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__54905\,
            I => \N__54873\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__54902\,
            I => \N__54873\
        );

    \I__11185\ : Odrv4
    port map (
            O => \N__54895\,
            I => n146
        );

    \I__11184\ : Odrv12
    port map (
            O => \N__54886\,
            I => n146
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__54883\,
            I => n146
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__54880\,
            I => n146
        );

    \I__11181\ : Odrv4
    port map (
            O => \N__54873\,
            I => n146
        );

    \I__11180\ : CascadeMux
    port map (
            O => \N__54862\,
            I => \N__54859\
        );

    \I__11179\ : InMux
    port map (
            O => \N__54859\,
            I => \N__54856\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__54856\,
            I => \N__54853\
        );

    \I__11177\ : Span4Mux_v
    port map (
            O => \N__54853\,
            I => \N__54850\
        );

    \I__11176\ : Odrv4
    port map (
            O => \N__54850\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n742\
        );

    \I__11175\ : InMux
    port map (
            O => \N__54847\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17749\
        );

    \I__11174\ : InMux
    port map (
            O => \N__54844\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n743\
        );

    \I__11173\ : CascadeMux
    port map (
            O => \N__54841\,
            I => \N__54838\
        );

    \I__11172\ : InMux
    port map (
            O => \N__54838\,
            I => \N__54835\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__54835\,
            I => \N__54832\
        );

    \I__11170\ : Span4Mux_h
    port map (
            O => \N__54832\,
            I => \N__54829\
        );

    \I__11169\ : Odrv4
    port map (
            O => \N__54829\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_CO\
        );

    \I__11168\ : InMux
    port map (
            O => \N__54826\,
            I => \N__54823\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__54823\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n57\
        );

    \I__11166\ : InMux
    port map (
            O => \N__54820\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17736\
        );

    \I__11165\ : InMux
    port map (
            O => \N__54817\,
            I => \N__54814\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__54814\,
            I => \N__54810\
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__54813\,
            I => \N__54807\
        );

    \I__11162\ : Span4Mux_v
    port map (
            O => \N__54810\,
            I => \N__54793\
        );

    \I__11161\ : InMux
    port map (
            O => \N__54807\,
            I => \N__54790\
        );

    \I__11160\ : CascadeMux
    port map (
            O => \N__54806\,
            I => \N__54787\
        );

    \I__11159\ : CascadeMux
    port map (
            O => \N__54805\,
            I => \N__54784\
        );

    \I__11158\ : CascadeMux
    port map (
            O => \N__54804\,
            I => \N__54781\
        );

    \I__11157\ : CascadeMux
    port map (
            O => \N__54803\,
            I => \N__54778\
        );

    \I__11156\ : CascadeMux
    port map (
            O => \N__54802\,
            I => \N__54775\
        );

    \I__11155\ : InMux
    port map (
            O => \N__54801\,
            I => \N__54765\
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__54800\,
            I => \N__54762\
        );

    \I__11153\ : CascadeMux
    port map (
            O => \N__54799\,
            I => \N__54758\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__54798\,
            I => \N__54754\
        );

    \I__11151\ : CascadeMux
    port map (
            O => \N__54797\,
            I => \N__54751\
        );

    \I__11150\ : CascadeMux
    port map (
            O => \N__54796\,
            I => \N__54747\
        );

    \I__11149\ : Span4Mux_h
    port map (
            O => \N__54793\,
            I => \N__54742\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__54790\,
            I => \N__54742\
        );

    \I__11147\ : InMux
    port map (
            O => \N__54787\,
            I => \N__54739\
        );

    \I__11146\ : InMux
    port map (
            O => \N__54784\,
            I => \N__54736\
        );

    \I__11145\ : InMux
    port map (
            O => \N__54781\,
            I => \N__54733\
        );

    \I__11144\ : InMux
    port map (
            O => \N__54778\,
            I => \N__54730\
        );

    \I__11143\ : InMux
    port map (
            O => \N__54775\,
            I => \N__54727\
        );

    \I__11142\ : CascadeMux
    port map (
            O => \N__54774\,
            I => \N__54724\
        );

    \I__11141\ : CascadeMux
    port map (
            O => \N__54773\,
            I => \N__54721\
        );

    \I__11140\ : CascadeMux
    port map (
            O => \N__54772\,
            I => \N__54718\
        );

    \I__11139\ : CascadeMux
    port map (
            O => \N__54771\,
            I => \N__54715\
        );

    \I__11138\ : CascadeMux
    port map (
            O => \N__54770\,
            I => \N__54710\
        );

    \I__11137\ : CascadeMux
    port map (
            O => \N__54769\,
            I => \N__54706\
        );

    \I__11136\ : CascadeMux
    port map (
            O => \N__54768\,
            I => \N__54702\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__54765\,
            I => \N__54699\
        );

    \I__11134\ : InMux
    port map (
            O => \N__54762\,
            I => \N__54696\
        );

    \I__11133\ : InMux
    port map (
            O => \N__54761\,
            I => \N__54681\
        );

    \I__11132\ : InMux
    port map (
            O => \N__54758\,
            I => \N__54681\
        );

    \I__11131\ : InMux
    port map (
            O => \N__54757\,
            I => \N__54681\
        );

    \I__11130\ : InMux
    port map (
            O => \N__54754\,
            I => \N__54681\
        );

    \I__11129\ : InMux
    port map (
            O => \N__54751\,
            I => \N__54681\
        );

    \I__11128\ : InMux
    port map (
            O => \N__54750\,
            I => \N__54681\
        );

    \I__11127\ : InMux
    port map (
            O => \N__54747\,
            I => \N__54681\
        );

    \I__11126\ : Span4Mux_v
    port map (
            O => \N__54742\,
            I => \N__54675\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__54739\,
            I => \N__54675\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__54736\,
            I => \N__54672\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__54733\,
            I => \N__54665\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__54730\,
            I => \N__54665\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__54727\,
            I => \N__54665\
        );

    \I__11120\ : InMux
    port map (
            O => \N__54724\,
            I => \N__54662\
        );

    \I__11119\ : InMux
    port map (
            O => \N__54721\,
            I => \N__54659\
        );

    \I__11118\ : InMux
    port map (
            O => \N__54718\,
            I => \N__54656\
        );

    \I__11117\ : InMux
    port map (
            O => \N__54715\,
            I => \N__54653\
        );

    \I__11116\ : CascadeMux
    port map (
            O => \N__54714\,
            I => \N__54650\
        );

    \I__11115\ : InMux
    port map (
            O => \N__54713\,
            I => \N__54637\
        );

    \I__11114\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54637\
        );

    \I__11113\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54637\
        );

    \I__11112\ : InMux
    port map (
            O => \N__54706\,
            I => \N__54637\
        );

    \I__11111\ : InMux
    port map (
            O => \N__54705\,
            I => \N__54637\
        );

    \I__11110\ : InMux
    port map (
            O => \N__54702\,
            I => \N__54637\
        );

    \I__11109\ : Span4Mux_v
    port map (
            O => \N__54699\,
            I => \N__54632\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__54696\,
            I => \N__54632\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__54681\,
            I => \N__54629\
        );

    \I__11106\ : CascadeMux
    port map (
            O => \N__54680\,
            I => \N__54626\
        );

    \I__11105\ : Span4Mux_v
    port map (
            O => \N__54675\,
            I => \N__54620\
        );

    \I__11104\ : Span4Mux_h
    port map (
            O => \N__54672\,
            I => \N__54620\
        );

    \I__11103\ : Span4Mux_v
    port map (
            O => \N__54665\,
            I => \N__54609\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__54662\,
            I => \N__54609\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__54659\,
            I => \N__54609\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__54656\,
            I => \N__54609\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__54653\,
            I => \N__54609\
        );

    \I__11098\ : InMux
    port map (
            O => \N__54650\,
            I => \N__54606\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__54637\,
            I => \N__54599\
        );

    \I__11096\ : Span4Mux_v
    port map (
            O => \N__54632\,
            I => \N__54599\
        );

    \I__11095\ : Span4Mux_v
    port map (
            O => \N__54629\,
            I => \N__54599\
        );

    \I__11094\ : InMux
    port map (
            O => \N__54626\,
            I => \N__54596\
        );

    \I__11093\ : CascadeMux
    port map (
            O => \N__54625\,
            I => \N__54593\
        );

    \I__11092\ : Span4Mux_v
    port map (
            O => \N__54620\,
            I => \N__54590\
        );

    \I__11091\ : Span4Mux_v
    port map (
            O => \N__54609\,
            I => \N__54585\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__54606\,
            I => \N__54585\
        );

    \I__11089\ : Span4Mux_h
    port map (
            O => \N__54599\,
            I => \N__54580\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__54596\,
            I => \N__54580\
        );

    \I__11087\ : InMux
    port map (
            O => \N__54593\,
            I => \N__54577\
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__54590\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n108\
        );

    \I__11085\ : Odrv4
    port map (
            O => \N__54585\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n108\
        );

    \I__11084\ : Odrv4
    port map (
            O => \N__54580\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n108\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__54577\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n108\
        );

    \I__11082\ : CascadeMux
    port map (
            O => \N__54568\,
            I => \N__54565\
        );

    \I__11081\ : InMux
    port map (
            O => \N__54565\,
            I => \N__54562\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__54562\,
            I => \N__54559\
        );

    \I__11079\ : Span4Mux_v
    port map (
            O => \N__54559\,
            I => \N__54556\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__54556\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n106\
        );

    \I__11077\ : InMux
    port map (
            O => \N__54553\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17737\
        );

    \I__11076\ : InMux
    port map (
            O => \N__54550\,
            I => \N__54547\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__54547\,
            I => \N__54544\
        );

    \I__11074\ : Span4Mux_v
    port map (
            O => \N__54544\,
            I => \N__54541\
        );

    \I__11073\ : Odrv4
    port map (
            O => \N__54541\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n155_adj_369\
        );

    \I__11072\ : CascadeMux
    port map (
            O => \N__54538\,
            I => \N__54535\
        );

    \I__11071\ : InMux
    port map (
            O => \N__54535\,
            I => \N__54531\
        );

    \I__11070\ : CascadeMux
    port map (
            O => \N__54534\,
            I => \N__54527\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__54531\,
            I => \N__54522\
        );

    \I__11068\ : CascadeMux
    port map (
            O => \N__54530\,
            I => \N__54518\
        );

    \I__11067\ : InMux
    port map (
            O => \N__54527\,
            I => \N__54513\
        );

    \I__11066\ : CascadeMux
    port map (
            O => \N__54526\,
            I => \N__54505\
        );

    \I__11065\ : CascadeMux
    port map (
            O => \N__54525\,
            I => \N__54502\
        );

    \I__11064\ : Span4Mux_v
    port map (
            O => \N__54522\,
            I => \N__54494\
        );

    \I__11063\ : InMux
    port map (
            O => \N__54521\,
            I => \N__54491\
        );

    \I__11062\ : InMux
    port map (
            O => \N__54518\,
            I => \N__54488\
        );

    \I__11061\ : CascadeMux
    port map (
            O => \N__54517\,
            I => \N__54485\
        );

    \I__11060\ : CascadeMux
    port map (
            O => \N__54516\,
            I => \N__54482\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__54513\,
            I => \N__54477\
        );

    \I__11058\ : CascadeMux
    port map (
            O => \N__54512\,
            I => \N__54474\
        );

    \I__11057\ : CascadeMux
    port map (
            O => \N__54511\,
            I => \N__54470\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__54510\,
            I => \N__54466\
        );

    \I__11055\ : CascadeMux
    port map (
            O => \N__54509\,
            I => \N__54463\
        );

    \I__11054\ : InMux
    port map (
            O => \N__54508\,
            I => \N__54460\
        );

    \I__11053\ : InMux
    port map (
            O => \N__54505\,
            I => \N__54457\
        );

    \I__11052\ : InMux
    port map (
            O => \N__54502\,
            I => \N__54454\
        );

    \I__11051\ : CascadeMux
    port map (
            O => \N__54501\,
            I => \N__54451\
        );

    \I__11050\ : CascadeMux
    port map (
            O => \N__54500\,
            I => \N__54446\
        );

    \I__11049\ : CascadeMux
    port map (
            O => \N__54499\,
            I => \N__54442\
        );

    \I__11048\ : CascadeMux
    port map (
            O => \N__54498\,
            I => \N__54438\
        );

    \I__11047\ : CascadeMux
    port map (
            O => \N__54497\,
            I => \N__54434\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__54494\,
            I => \N__54426\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__54491\,
            I => \N__54426\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__54488\,
            I => \N__54426\
        );

    \I__11043\ : InMux
    port map (
            O => \N__54485\,
            I => \N__54423\
        );

    \I__11042\ : InMux
    port map (
            O => \N__54482\,
            I => \N__54420\
        );

    \I__11041\ : CascadeMux
    port map (
            O => \N__54481\,
            I => \N__54417\
        );

    \I__11040\ : CascadeMux
    port map (
            O => \N__54480\,
            I => \N__54414\
        );

    \I__11039\ : Span4Mux_v
    port map (
            O => \N__54477\,
            I => \N__54411\
        );

    \I__11038\ : InMux
    port map (
            O => \N__54474\,
            I => \N__54400\
        );

    \I__11037\ : InMux
    port map (
            O => \N__54473\,
            I => \N__54400\
        );

    \I__11036\ : InMux
    port map (
            O => \N__54470\,
            I => \N__54400\
        );

    \I__11035\ : InMux
    port map (
            O => \N__54469\,
            I => \N__54400\
        );

    \I__11034\ : InMux
    port map (
            O => \N__54466\,
            I => \N__54400\
        );

    \I__11033\ : InMux
    port map (
            O => \N__54463\,
            I => \N__54397\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__54460\,
            I => \N__54390\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__54457\,
            I => \N__54390\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__54454\,
            I => \N__54390\
        );

    \I__11029\ : InMux
    port map (
            O => \N__54451\,
            I => \N__54387\
        );

    \I__11028\ : InMux
    port map (
            O => \N__54450\,
            I => \N__54383\
        );

    \I__11027\ : InMux
    port map (
            O => \N__54449\,
            I => \N__54374\
        );

    \I__11026\ : InMux
    port map (
            O => \N__54446\,
            I => \N__54374\
        );

    \I__11025\ : InMux
    port map (
            O => \N__54445\,
            I => \N__54374\
        );

    \I__11024\ : InMux
    port map (
            O => \N__54442\,
            I => \N__54374\
        );

    \I__11023\ : InMux
    port map (
            O => \N__54441\,
            I => \N__54365\
        );

    \I__11022\ : InMux
    port map (
            O => \N__54438\,
            I => \N__54365\
        );

    \I__11021\ : InMux
    port map (
            O => \N__54437\,
            I => \N__54365\
        );

    \I__11020\ : InMux
    port map (
            O => \N__54434\,
            I => \N__54365\
        );

    \I__11019\ : InMux
    port map (
            O => \N__54433\,
            I => \N__54362\
        );

    \I__11018\ : Span4Mux_v
    port map (
            O => \N__54426\,
            I => \N__54355\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__54423\,
            I => \N__54355\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__54420\,
            I => \N__54355\
        );

    \I__11015\ : InMux
    port map (
            O => \N__54417\,
            I => \N__54352\
        );

    \I__11014\ : InMux
    port map (
            O => \N__54414\,
            I => \N__54349\
        );

    \I__11013\ : Span4Mux_v
    port map (
            O => \N__54411\,
            I => \N__54344\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__54400\,
            I => \N__54344\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__54397\,
            I => \N__54341\
        );

    \I__11010\ : Span4Mux_v
    port map (
            O => \N__54390\,
            I => \N__54336\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__54387\,
            I => \N__54336\
        );

    \I__11008\ : CascadeMux
    port map (
            O => \N__54386\,
            I => \N__54333\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__54383\,
            I => \N__54324\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__54374\,
            I => \N__54324\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__54365\,
            I => \N__54324\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__54362\,
            I => \N__54324\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__54355\,
            I => \N__54317\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__54352\,
            I => \N__54317\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__54349\,
            I => \N__54317\
        );

    \I__11000\ : Span4Mux_v
    port map (
            O => \N__54344\,
            I => \N__54312\
        );

    \I__10999\ : Span4Mux_v
    port map (
            O => \N__54341\,
            I => \N__54312\
        );

    \I__10998\ : Span4Mux_v
    port map (
            O => \N__54336\,
            I => \N__54309\
        );

    \I__10997\ : InMux
    port map (
            O => \N__54333\,
            I => \N__54306\
        );

    \I__10996\ : Span12Mux_h
    port map (
            O => \N__54324\,
            I => \N__54303\
        );

    \I__10995\ : Span4Mux_v
    port map (
            O => \N__54317\,
            I => \N__54300\
        );

    \I__10994\ : Sp12to4
    port map (
            O => \N__54312\,
            I => \N__54293\
        );

    \I__10993\ : Sp12to4
    port map (
            O => \N__54309\,
            I => \N__54293\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__54306\,
            I => \N__54293\
        );

    \I__10991\ : Odrv12
    port map (
            O => \N__54303\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n111\
        );

    \I__10990\ : Odrv4
    port map (
            O => \N__54300\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n111\
        );

    \I__10989\ : Odrv12
    port map (
            O => \N__54293\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n111\
        );

    \I__10988\ : InMux
    port map (
            O => \N__54286\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17738\
        );

    \I__10987\ : InMux
    port map (
            O => \N__54283\,
            I => \N__54280\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__54280\,
            I => \N__54277\
        );

    \I__10985\ : Span4Mux_h
    port map (
            O => \N__54277\,
            I => \N__54274\
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__54274\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n204_adj_361\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__54271\,
            I => \N__54268\
        );

    \I__10982\ : InMux
    port map (
            O => \N__54268\,
            I => \N__54265\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__54265\,
            I => \N__54261\
        );

    \I__10980\ : CascadeMux
    port map (
            O => \N__54264\,
            I => \N__54258\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__54261\,
            I => \N__54245\
        );

    \I__10978\ : InMux
    port map (
            O => \N__54258\,
            I => \N__54242\
        );

    \I__10977\ : CascadeMux
    port map (
            O => \N__54257\,
            I => \N__54239\
        );

    \I__10976\ : CascadeMux
    port map (
            O => \N__54256\,
            I => \N__54236\
        );

    \I__10975\ : CascadeMux
    port map (
            O => \N__54255\,
            I => \N__54233\
        );

    \I__10974\ : CascadeMux
    port map (
            O => \N__54254\,
            I => \N__54229\
        );

    \I__10973\ : CascadeMux
    port map (
            O => \N__54253\,
            I => \N__54225\
        );

    \I__10972\ : CascadeMux
    port map (
            O => \N__54252\,
            I => \N__54221\
        );

    \I__10971\ : CascadeMux
    port map (
            O => \N__54251\,
            I => \N__54217\
        );

    \I__10970\ : CascadeMux
    port map (
            O => \N__54250\,
            I => \N__54214\
        );

    \I__10969\ : CascadeMux
    port map (
            O => \N__54249\,
            I => \N__54211\
        );

    \I__10968\ : CascadeMux
    port map (
            O => \N__54248\,
            I => \N__54208\
        );

    \I__10967\ : Span4Mux_v
    port map (
            O => \N__54245\,
            I => \N__54202\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__54242\,
            I => \N__54202\
        );

    \I__10965\ : InMux
    port map (
            O => \N__54239\,
            I => \N__54199\
        );

    \I__10964\ : InMux
    port map (
            O => \N__54236\,
            I => \N__54196\
        );

    \I__10963\ : InMux
    port map (
            O => \N__54233\,
            I => \N__54190\
        );

    \I__10962\ : InMux
    port map (
            O => \N__54232\,
            I => \N__54177\
        );

    \I__10961\ : InMux
    port map (
            O => \N__54229\,
            I => \N__54177\
        );

    \I__10960\ : InMux
    port map (
            O => \N__54228\,
            I => \N__54177\
        );

    \I__10959\ : InMux
    port map (
            O => \N__54225\,
            I => \N__54177\
        );

    \I__10958\ : InMux
    port map (
            O => \N__54224\,
            I => \N__54177\
        );

    \I__10957\ : InMux
    port map (
            O => \N__54221\,
            I => \N__54177\
        );

    \I__10956\ : CascadeMux
    port map (
            O => \N__54220\,
            I => \N__54172\
        );

    \I__10955\ : InMux
    port map (
            O => \N__54217\,
            I => \N__54169\
        );

    \I__10954\ : InMux
    port map (
            O => \N__54214\,
            I => \N__54166\
        );

    \I__10953\ : InMux
    port map (
            O => \N__54211\,
            I => \N__54163\
        );

    \I__10952\ : InMux
    port map (
            O => \N__54208\,
            I => \N__54160\
        );

    \I__10951\ : CascadeMux
    port map (
            O => \N__54207\,
            I => \N__54157\
        );

    \I__10950\ : Span4Mux_h
    port map (
            O => \N__54202\,
            I => \N__54153\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__54199\,
            I => \N__54148\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__54196\,
            I => \N__54148\
        );

    \I__10947\ : CascadeMux
    port map (
            O => \N__54195\,
            I => \N__54145\
        );

    \I__10946\ : CascadeMux
    port map (
            O => \N__54194\,
            I => \N__54142\
        );

    \I__10945\ : CascadeMux
    port map (
            O => \N__54193\,
            I => \N__54139\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__54190\,
            I => \N__54132\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__54177\,
            I => \N__54129\
        );

    \I__10942\ : InMux
    port map (
            O => \N__54176\,
            I => \N__54126\
        );

    \I__10941\ : InMux
    port map (
            O => \N__54175\,
            I => \N__54123\
        );

    \I__10940\ : InMux
    port map (
            O => \N__54172\,
            I => \N__54120\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__54169\,
            I => \N__54111\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__54166\,
            I => \N__54111\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__54163\,
            I => \N__54111\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__54160\,
            I => \N__54111\
        );

    \I__10935\ : InMux
    port map (
            O => \N__54157\,
            I => \N__54108\
        );

    \I__10934\ : CascadeMux
    port map (
            O => \N__54156\,
            I => \N__54105\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__54153\,
            I => \N__54100\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__54148\,
            I => \N__54100\
        );

    \I__10931\ : InMux
    port map (
            O => \N__54145\,
            I => \N__54091\
        );

    \I__10930\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54091\
        );

    \I__10929\ : InMux
    port map (
            O => \N__54139\,
            I => \N__54091\
        );

    \I__10928\ : InMux
    port map (
            O => \N__54138\,
            I => \N__54091\
        );

    \I__10927\ : CascadeMux
    port map (
            O => \N__54137\,
            I => \N__54088\
        );

    \I__10926\ : CascadeMux
    port map (
            O => \N__54136\,
            I => \N__54085\
        );

    \I__10925\ : CascadeMux
    port map (
            O => \N__54135\,
            I => \N__54081\
        );

    \I__10924\ : Span4Mux_h
    port map (
            O => \N__54132\,
            I => \N__54077\
        );

    \I__10923\ : Span4Mux_v
    port map (
            O => \N__54129\,
            I => \N__54070\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__54126\,
            I => \N__54070\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__54123\,
            I => \N__54070\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__54120\,
            I => \N__54063\
        );

    \I__10919\ : Span4Mux_v
    port map (
            O => \N__54111\,
            I => \N__54063\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__54108\,
            I => \N__54063\
        );

    \I__10917\ : InMux
    port map (
            O => \N__54105\,
            I => \N__54060\
        );

    \I__10916\ : Span4Mux_v
    port map (
            O => \N__54100\,
            I => \N__54055\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__54091\,
            I => \N__54055\
        );

    \I__10914\ : InMux
    port map (
            O => \N__54088\,
            I => \N__54046\
        );

    \I__10913\ : InMux
    port map (
            O => \N__54085\,
            I => \N__54046\
        );

    \I__10912\ : InMux
    port map (
            O => \N__54084\,
            I => \N__54046\
        );

    \I__10911\ : InMux
    port map (
            O => \N__54081\,
            I => \N__54046\
        );

    \I__10910\ : CascadeMux
    port map (
            O => \N__54080\,
            I => \N__54043\
        );

    \I__10909\ : Span4Mux_v
    port map (
            O => \N__54077\,
            I => \N__54038\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__54070\,
            I => \N__54038\
        );

    \I__10907\ : Span4Mux_v
    port map (
            O => \N__54063\,
            I => \N__54033\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__54060\,
            I => \N__54033\
        );

    \I__10905\ : Sp12to4
    port map (
            O => \N__54055\,
            I => \N__54028\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__54046\,
            I => \N__54028\
        );

    \I__10903\ : InMux
    port map (
            O => \N__54043\,
            I => \N__54025\
        );

    \I__10902\ : Odrv4
    port map (
            O => \N__54038\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n114\
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__54033\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n114\
        );

    \I__10900\ : Odrv12
    port map (
            O => \N__54028\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n114\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__54025\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n114\
        );

    \I__10898\ : InMux
    port map (
            O => \N__54016\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17739\
        );

    \I__10897\ : InMux
    port map (
            O => \N__54013\,
            I => \N__54010\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__54010\,
            I => \N__54007\
        );

    \I__10895\ : Span4Mux_h
    port map (
            O => \N__54007\,
            I => \N__54004\
        );

    \I__10894\ : Odrv4
    port map (
            O => \N__54004\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n253\
        );

    \I__10893\ : CascadeMux
    port map (
            O => \N__54001\,
            I => \N__53996\
        );

    \I__10892\ : CascadeMux
    port map (
            O => \N__54000\,
            I => \N__53993\
        );

    \I__10891\ : CascadeMux
    port map (
            O => \N__53999\,
            I => \N__53987\
        );

    \I__10890\ : InMux
    port map (
            O => \N__53996\,
            I => \N__53983\
        );

    \I__10889\ : InMux
    port map (
            O => \N__53993\,
            I => \N__53980\
        );

    \I__10888\ : CascadeMux
    port map (
            O => \N__53992\,
            I => \N__53977\
        );

    \I__10887\ : CascadeMux
    port map (
            O => \N__53991\,
            I => \N__53974\
        );

    \I__10886\ : CascadeMux
    port map (
            O => \N__53990\,
            I => \N__53971\
        );

    \I__10885\ : InMux
    port map (
            O => \N__53987\,
            I => \N__53966\
        );

    \I__10884\ : CascadeMux
    port map (
            O => \N__53986\,
            I => \N__53963\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__53983\,
            I => \N__53958\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__53980\,
            I => \N__53958\
        );

    \I__10881\ : InMux
    port map (
            O => \N__53977\,
            I => \N__53955\
        );

    \I__10880\ : InMux
    port map (
            O => \N__53974\,
            I => \N__53952\
        );

    \I__10879\ : InMux
    port map (
            O => \N__53971\,
            I => \N__53949\
        );

    \I__10878\ : CascadeMux
    port map (
            O => \N__53970\,
            I => \N__53946\
        );

    \I__10877\ : CascadeMux
    port map (
            O => \N__53969\,
            I => \N__53943\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__53966\,
            I => \N__53934\
        );

    \I__10875\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53931\
        );

    \I__10874\ : Span4Mux_v
    port map (
            O => \N__53958\,
            I => \N__53922\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__53955\,
            I => \N__53922\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__53952\,
            I => \N__53922\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__53949\,
            I => \N__53922\
        );

    \I__10870\ : InMux
    port map (
            O => \N__53946\,
            I => \N__53919\
        );

    \I__10869\ : InMux
    port map (
            O => \N__53943\,
            I => \N__53916\
        );

    \I__10868\ : CascadeMux
    port map (
            O => \N__53942\,
            I => \N__53912\
        );

    \I__10867\ : CascadeMux
    port map (
            O => \N__53941\,
            I => \N__53908\
        );

    \I__10866\ : CascadeMux
    port map (
            O => \N__53940\,
            I => \N__53904\
        );

    \I__10865\ : CascadeMux
    port map (
            O => \N__53939\,
            I => \N__53900\
        );

    \I__10864\ : CascadeMux
    port map (
            O => \N__53938\,
            I => \N__53897\
        );

    \I__10863\ : CascadeMux
    port map (
            O => \N__53937\,
            I => \N__53894\
        );

    \I__10862\ : Span4Mux_v
    port map (
            O => \N__53934\,
            I => \N__53889\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__53931\,
            I => \N__53889\
        );

    \I__10860\ : Span4Mux_v
    port map (
            O => \N__53922\,
            I => \N__53876\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__53919\,
            I => \N__53876\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__53916\,
            I => \N__53873\
        );

    \I__10857\ : InMux
    port map (
            O => \N__53915\,
            I => \N__53870\
        );

    \I__10856\ : InMux
    port map (
            O => \N__53912\,
            I => \N__53867\
        );

    \I__10855\ : InMux
    port map (
            O => \N__53911\,
            I => \N__53854\
        );

    \I__10854\ : InMux
    port map (
            O => \N__53908\,
            I => \N__53854\
        );

    \I__10853\ : InMux
    port map (
            O => \N__53907\,
            I => \N__53854\
        );

    \I__10852\ : InMux
    port map (
            O => \N__53904\,
            I => \N__53854\
        );

    \I__10851\ : InMux
    port map (
            O => \N__53903\,
            I => \N__53854\
        );

    \I__10850\ : InMux
    port map (
            O => \N__53900\,
            I => \N__53854\
        );

    \I__10849\ : InMux
    port map (
            O => \N__53897\,
            I => \N__53851\
        );

    \I__10848\ : InMux
    port map (
            O => \N__53894\,
            I => \N__53848\
        );

    \I__10847\ : Span4Mux_h
    port map (
            O => \N__53889\,
            I => \N__53845\
        );

    \I__10846\ : InMux
    port map (
            O => \N__53888\,
            I => \N__53842\
        );

    \I__10845\ : CascadeMux
    port map (
            O => \N__53887\,
            I => \N__53839\
        );

    \I__10844\ : CascadeMux
    port map (
            O => \N__53886\,
            I => \N__53836\
        );

    \I__10843\ : CascadeMux
    port map (
            O => \N__53885\,
            I => \N__53833\
        );

    \I__10842\ : CascadeMux
    port map (
            O => \N__53884\,
            I => \N__53829\
        );

    \I__10841\ : CascadeMux
    port map (
            O => \N__53883\,
            I => \N__53826\
        );

    \I__10840\ : CascadeMux
    port map (
            O => \N__53882\,
            I => \N__53823\
        );

    \I__10839\ : CascadeMux
    port map (
            O => \N__53881\,
            I => \N__53820\
        );

    \I__10838\ : Span4Mux_v
    port map (
            O => \N__53876\,
            I => \N__53816\
        );

    \I__10837\ : Span4Mux_v
    port map (
            O => \N__53873\,
            I => \N__53805\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__53870\,
            I => \N__53805\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__53867\,
            I => \N__53805\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__53854\,
            I => \N__53805\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__53851\,
            I => \N__53805\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__53848\,
            I => \N__53802\
        );

    \I__10831\ : Span4Mux_v
    port map (
            O => \N__53845\,
            I => \N__53799\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__53842\,
            I => \N__53796\
        );

    \I__10829\ : InMux
    port map (
            O => \N__53839\,
            I => \N__53785\
        );

    \I__10828\ : InMux
    port map (
            O => \N__53836\,
            I => \N__53785\
        );

    \I__10827\ : InMux
    port map (
            O => \N__53833\,
            I => \N__53785\
        );

    \I__10826\ : InMux
    port map (
            O => \N__53832\,
            I => \N__53785\
        );

    \I__10825\ : InMux
    port map (
            O => \N__53829\,
            I => \N__53785\
        );

    \I__10824\ : InMux
    port map (
            O => \N__53826\,
            I => \N__53778\
        );

    \I__10823\ : InMux
    port map (
            O => \N__53823\,
            I => \N__53778\
        );

    \I__10822\ : InMux
    port map (
            O => \N__53820\,
            I => \N__53778\
        );

    \I__10821\ : CascadeMux
    port map (
            O => \N__53819\,
            I => \N__53775\
        );

    \I__10820\ : Span4Mux_h
    port map (
            O => \N__53816\,
            I => \N__53772\
        );

    \I__10819\ : Span4Mux_v
    port map (
            O => \N__53805\,
            I => \N__53769\
        );

    \I__10818\ : Span4Mux_h
    port map (
            O => \N__53802\,
            I => \N__53766\
        );

    \I__10817\ : Span4Mux_v
    port map (
            O => \N__53799\,
            I => \N__53757\
        );

    \I__10816\ : Span4Mux_h
    port map (
            O => \N__53796\,
            I => \N__53757\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__53785\,
            I => \N__53757\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__53778\,
            I => \N__53757\
        );

    \I__10813\ : InMux
    port map (
            O => \N__53775\,
            I => \N__53754\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__53772\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n117\
        );

    \I__10811\ : Odrv4
    port map (
            O => \N__53769\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n117\
        );

    \I__10810\ : Odrv4
    port map (
            O => \N__53766\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n117\
        );

    \I__10809\ : Odrv4
    port map (
            O => \N__53757\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n117\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__53754\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n117\
        );

    \I__10807\ : InMux
    port map (
            O => \N__53743\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17740\
        );

    \I__10806\ : InMux
    port map (
            O => \N__53740\,
            I => \N__53737\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__53737\,
            I => \N__53734\
        );

    \I__10804\ : Span4Mux_h
    port map (
            O => \N__53734\,
            I => \N__53731\
        );

    \I__10803\ : Odrv4
    port map (
            O => \N__53731\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n302_adj_364\
        );

    \I__10802\ : CascadeMux
    port map (
            O => \N__53728\,
            I => \N__53725\
        );

    \I__10801\ : InMux
    port map (
            O => \N__53725\,
            I => \N__53719\
        );

    \I__10800\ : CascadeMux
    port map (
            O => \N__53724\,
            I => \N__53716\
        );

    \I__10799\ : CascadeMux
    port map (
            O => \N__53723\,
            I => \N__53712\
        );

    \I__10798\ : CascadeMux
    port map (
            O => \N__53722\,
            I => \N__53708\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__53719\,
            I => \N__53702\
        );

    \I__10796\ : InMux
    port map (
            O => \N__53716\,
            I => \N__53699\
        );

    \I__10795\ : CascadeMux
    port map (
            O => \N__53715\,
            I => \N__53696\
        );

    \I__10794\ : InMux
    port map (
            O => \N__53712\,
            I => \N__53690\
        );

    \I__10793\ : CascadeMux
    port map (
            O => \N__53711\,
            I => \N__53687\
        );

    \I__10792\ : InMux
    port map (
            O => \N__53708\,
            I => \N__53684\
        );

    \I__10791\ : CascadeMux
    port map (
            O => \N__53707\,
            I => \N__53681\
        );

    \I__10790\ : CascadeMux
    port map (
            O => \N__53706\,
            I => \N__53677\
        );

    \I__10789\ : InMux
    port map (
            O => \N__53705\,
            I => \N__53674\
        );

    \I__10788\ : Span4Mux_v
    port map (
            O => \N__53702\,
            I => \N__53669\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__53699\,
            I => \N__53669\
        );

    \I__10786\ : InMux
    port map (
            O => \N__53696\,
            I => \N__53666\
        );

    \I__10785\ : CascadeMux
    port map (
            O => \N__53695\,
            I => \N__53662\
        );

    \I__10784\ : CascadeMux
    port map (
            O => \N__53694\,
            I => \N__53658\
        );

    \I__10783\ : CascadeMux
    port map (
            O => \N__53693\,
            I => \N__53654\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__53690\,
            I => \N__53651\
        );

    \I__10781\ : InMux
    port map (
            O => \N__53687\,
            I => \N__53647\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__53684\,
            I => \N__53644\
        );

    \I__10779\ : InMux
    port map (
            O => \N__53681\,
            I => \N__53641\
        );

    \I__10778\ : InMux
    port map (
            O => \N__53680\,
            I => \N__53638\
        );

    \I__10777\ : InMux
    port map (
            O => \N__53677\,
            I => \N__53633\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__53674\,
            I => \N__53630\
        );

    \I__10775\ : Span4Mux_h
    port map (
            O => \N__53669\,
            I => \N__53625\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__53666\,
            I => \N__53625\
        );

    \I__10773\ : InMux
    port map (
            O => \N__53665\,
            I => \N__53612\
        );

    \I__10772\ : InMux
    port map (
            O => \N__53662\,
            I => \N__53612\
        );

    \I__10771\ : InMux
    port map (
            O => \N__53661\,
            I => \N__53612\
        );

    \I__10770\ : InMux
    port map (
            O => \N__53658\,
            I => \N__53612\
        );

    \I__10769\ : InMux
    port map (
            O => \N__53657\,
            I => \N__53612\
        );

    \I__10768\ : InMux
    port map (
            O => \N__53654\,
            I => \N__53612\
        );

    \I__10767\ : Span4Mux_v
    port map (
            O => \N__53651\,
            I => \N__53604\
        );

    \I__10766\ : InMux
    port map (
            O => \N__53650\,
            I => \N__53601\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__53647\,
            I => \N__53592\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__53644\,
            I => \N__53592\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__53641\,
            I => \N__53592\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__53638\,
            I => \N__53592\
        );

    \I__10761\ : InMux
    port map (
            O => \N__53637\,
            I => \N__53589\
        );

    \I__10760\ : CascadeMux
    port map (
            O => \N__53636\,
            I => \N__53586\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__53633\,
            I => \N__53582\
        );

    \I__10758\ : Span4Mux_v
    port map (
            O => \N__53630\,
            I => \N__53575\
        );

    \I__10757\ : Span4Mux_h
    port map (
            O => \N__53625\,
            I => \N__53575\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__53612\,
            I => \N__53575\
        );

    \I__10755\ : InMux
    port map (
            O => \N__53611\,
            I => \N__53572\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__53610\,
            I => \N__53569\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__53609\,
            I => \N__53564\
        );

    \I__10752\ : CascadeMux
    port map (
            O => \N__53608\,
            I => \N__53560\
        );

    \I__10751\ : CascadeMux
    port map (
            O => \N__53607\,
            I => \N__53556\
        );

    \I__10750\ : Span4Mux_h
    port map (
            O => \N__53604\,
            I => \N__53547\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__53601\,
            I => \N__53547\
        );

    \I__10748\ : Span4Mux_v
    port map (
            O => \N__53592\,
            I => \N__53547\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__53589\,
            I => \N__53547\
        );

    \I__10746\ : InMux
    port map (
            O => \N__53586\,
            I => \N__53544\
        );

    \I__10745\ : CascadeMux
    port map (
            O => \N__53585\,
            I => \N__53541\
        );

    \I__10744\ : Span4Mux_v
    port map (
            O => \N__53582\,
            I => \N__53534\
        );

    \I__10743\ : Span4Mux_v
    port map (
            O => \N__53575\,
            I => \N__53534\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__53572\,
            I => \N__53534\
        );

    \I__10741\ : InMux
    port map (
            O => \N__53569\,
            I => \N__53529\
        );

    \I__10740\ : InMux
    port map (
            O => \N__53568\,
            I => \N__53529\
        );

    \I__10739\ : InMux
    port map (
            O => \N__53567\,
            I => \N__53516\
        );

    \I__10738\ : InMux
    port map (
            O => \N__53564\,
            I => \N__53516\
        );

    \I__10737\ : InMux
    port map (
            O => \N__53563\,
            I => \N__53516\
        );

    \I__10736\ : InMux
    port map (
            O => \N__53560\,
            I => \N__53516\
        );

    \I__10735\ : InMux
    port map (
            O => \N__53559\,
            I => \N__53516\
        );

    \I__10734\ : InMux
    port map (
            O => \N__53556\,
            I => \N__53516\
        );

    \I__10733\ : Span4Mux_v
    port map (
            O => \N__53547\,
            I => \N__53511\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__53544\,
            I => \N__53511\
        );

    \I__10731\ : InMux
    port map (
            O => \N__53541\,
            I => \N__53508\
        );

    \I__10730\ : Sp12to4
    port map (
            O => \N__53534\,
            I => \N__53501\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__53529\,
            I => \N__53501\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__53516\,
            I => \N__53501\
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__53511\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n120\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__53508\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n120\
        );

    \I__10725\ : Odrv12
    port map (
            O => \N__53501\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n120\
        );

    \I__10724\ : InMux
    port map (
            O => \N__53494\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17741\
        );

    \I__10723\ : InMux
    port map (
            O => \N__53491\,
            I => \N__53488\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__53488\,
            I => \N__53485\
        );

    \I__10721\ : Span4Mux_v
    port map (
            O => \N__53485\,
            I => \N__53482\
        );

    \I__10720\ : Odrv4
    port map (
            O => \N__53482\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n351\
        );

    \I__10719\ : InMux
    port map (
            O => \N__53479\,
            I => \N__53475\
        );

    \I__10718\ : CascadeMux
    port map (
            O => \N__53478\,
            I => \N__53471\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__53475\,
            I => \N__53461\
        );

    \I__10716\ : InMux
    port map (
            O => \N__53474\,
            I => \N__53458\
        );

    \I__10715\ : InMux
    port map (
            O => \N__53471\,
            I => \N__53455\
        );

    \I__10714\ : CascadeMux
    port map (
            O => \N__53470\,
            I => \N__53452\
        );

    \I__10713\ : CascadeMux
    port map (
            O => \N__53469\,
            I => \N__53449\
        );

    \I__10712\ : CascadeMux
    port map (
            O => \N__53468\,
            I => \N__53446\
        );

    \I__10711\ : CascadeMux
    port map (
            O => \N__53467\,
            I => \N__53442\
        );

    \I__10710\ : CascadeMux
    port map (
            O => \N__53466\,
            I => \N__53439\
        );

    \I__10709\ : CascadeMux
    port map (
            O => \N__53465\,
            I => \N__53435\
        );

    \I__10708\ : CascadeMux
    port map (
            O => \N__53464\,
            I => \N__53431\
        );

    \I__10707\ : Span4Mux_v
    port map (
            O => \N__53461\,
            I => \N__53423\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__53458\,
            I => \N__53420\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__53455\,
            I => \N__53417\
        );

    \I__10704\ : InMux
    port map (
            O => \N__53452\,
            I => \N__53414\
        );

    \I__10703\ : InMux
    port map (
            O => \N__53449\,
            I => \N__53411\
        );

    \I__10702\ : InMux
    port map (
            O => \N__53446\,
            I => \N__53405\
        );

    \I__10701\ : InMux
    port map (
            O => \N__53445\,
            I => \N__53390\
        );

    \I__10700\ : InMux
    port map (
            O => \N__53442\,
            I => \N__53390\
        );

    \I__10699\ : InMux
    port map (
            O => \N__53439\,
            I => \N__53390\
        );

    \I__10698\ : InMux
    port map (
            O => \N__53438\,
            I => \N__53390\
        );

    \I__10697\ : InMux
    port map (
            O => \N__53435\,
            I => \N__53390\
        );

    \I__10696\ : InMux
    port map (
            O => \N__53434\,
            I => \N__53390\
        );

    \I__10695\ : InMux
    port map (
            O => \N__53431\,
            I => \N__53390\
        );

    \I__10694\ : CascadeMux
    port map (
            O => \N__53430\,
            I => \N__53387\
        );

    \I__10693\ : CascadeMux
    port map (
            O => \N__53429\,
            I => \N__53383\
        );

    \I__10692\ : CascadeMux
    port map (
            O => \N__53428\,
            I => \N__53379\
        );

    \I__10691\ : CascadeMux
    port map (
            O => \N__53427\,
            I => \N__53374\
        );

    \I__10690\ : InMux
    port map (
            O => \N__53426\,
            I => \N__53370\
        );

    \I__10689\ : Span4Mux_v
    port map (
            O => \N__53423\,
            I => \N__53364\
        );

    \I__10688\ : Span4Mux_v
    port map (
            O => \N__53420\,
            I => \N__53364\
        );

    \I__10687\ : Span4Mux_h
    port map (
            O => \N__53417\,
            I => \N__53359\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__53414\,
            I => \N__53359\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__53411\,
            I => \N__53356\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__53410\,
            I => \N__53353\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__53409\,
            I => \N__53350\
        );

    \I__10682\ : CascadeMux
    port map (
            O => \N__53408\,
            I => \N__53347\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__53405\,
            I => \N__53342\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__53390\,
            I => \N__53342\
        );

    \I__10679\ : InMux
    port map (
            O => \N__53387\,
            I => \N__53329\
        );

    \I__10678\ : InMux
    port map (
            O => \N__53386\,
            I => \N__53329\
        );

    \I__10677\ : InMux
    port map (
            O => \N__53383\,
            I => \N__53329\
        );

    \I__10676\ : InMux
    port map (
            O => \N__53382\,
            I => \N__53329\
        );

    \I__10675\ : InMux
    port map (
            O => \N__53379\,
            I => \N__53329\
        );

    \I__10674\ : InMux
    port map (
            O => \N__53378\,
            I => \N__53329\
        );

    \I__10673\ : InMux
    port map (
            O => \N__53377\,
            I => \N__53326\
        );

    \I__10672\ : InMux
    port map (
            O => \N__53374\,
            I => \N__53323\
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__53373\,
            I => \N__53320\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__53370\,
            I => \N__53317\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__53369\,
            I => \N__53313\
        );

    \I__10668\ : Span4Mux_h
    port map (
            O => \N__53364\,
            I => \N__53306\
        );

    \I__10667\ : Span4Mux_v
    port map (
            O => \N__53359\,
            I => \N__53306\
        );

    \I__10666\ : Span4Mux_v
    port map (
            O => \N__53356\,
            I => \N__53306\
        );

    \I__10665\ : InMux
    port map (
            O => \N__53353\,
            I => \N__53303\
        );

    \I__10664\ : InMux
    port map (
            O => \N__53350\,
            I => \N__53300\
        );

    \I__10663\ : InMux
    port map (
            O => \N__53347\,
            I => \N__53297\
        );

    \I__10662\ : Span4Mux_v
    port map (
            O => \N__53342\,
            I => \N__53288\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__53329\,
            I => \N__53288\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__53326\,
            I => \N__53288\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__53323\,
            I => \N__53288\
        );

    \I__10658\ : InMux
    port map (
            O => \N__53320\,
            I => \N__53285\
        );

    \I__10657\ : Span4Mux_v
    port map (
            O => \N__53317\,
            I => \N__53281\
        );

    \I__10656\ : InMux
    port map (
            O => \N__53316\,
            I => \N__53278\
        );

    \I__10655\ : InMux
    port map (
            O => \N__53313\,
            I => \N__53275\
        );

    \I__10654\ : Span4Mux_h
    port map (
            O => \N__53306\,
            I => \N__53262\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__53303\,
            I => \N__53262\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__53300\,
            I => \N__53262\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__53297\,
            I => \N__53262\
        );

    \I__10650\ : Span4Mux_v
    port map (
            O => \N__53288\,
            I => \N__53262\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__53285\,
            I => \N__53262\
        );

    \I__10648\ : CascadeMux
    port map (
            O => \N__53284\,
            I => \N__53259\
        );

    \I__10647\ : Span4Mux_h
    port map (
            O => \N__53281\,
            I => \N__53254\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__53278\,
            I => \N__53254\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__53275\,
            I => \N__53251\
        );

    \I__10644\ : Span4Mux_v
    port map (
            O => \N__53262\,
            I => \N__53248\
        );

    \I__10643\ : InMux
    port map (
            O => \N__53259\,
            I => \N__53245\
        );

    \I__10642\ : Span4Mux_v
    port map (
            O => \N__53254\,
            I => \N__53242\
        );

    \I__10641\ : Span4Mux_v
    port map (
            O => \N__53251\,
            I => \N__53239\
        );

    \I__10640\ : Sp12to4
    port map (
            O => \N__53248\,
            I => \N__53234\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__53245\,
            I => \N__53234\
        );

    \I__10638\ : Odrv4
    port map (
            O => \N__53242\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n123\
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__53239\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n123\
        );

    \I__10636\ : Odrv12
    port map (
            O => \N__53234\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n123\
        );

    \I__10635\ : InMux
    port map (
            O => \N__53227\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17742\
        );

    \I__10634\ : InMux
    port map (
            O => \N__53224\,
            I => \N__53221\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__53221\,
            I => \N__53218\
        );

    \I__10632\ : Odrv12
    port map (
            O => \N__53218\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n400_adj_511\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__53215\,
            I => \N__53212\
        );

    \I__10630\ : InMux
    port map (
            O => \N__53212\,
            I => \N__53207\
        );

    \I__10629\ : CascadeMux
    port map (
            O => \N__53211\,
            I => \N__53203\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__53210\,
            I => \N__53191\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__53207\,
            I => \N__53186\
        );

    \I__10626\ : InMux
    port map (
            O => \N__53206\,
            I => \N__53183\
        );

    \I__10625\ : InMux
    port map (
            O => \N__53203\,
            I => \N__53180\
        );

    \I__10624\ : CascadeMux
    port map (
            O => \N__53202\,
            I => \N__53177\
        );

    \I__10623\ : CascadeMux
    port map (
            O => \N__53201\,
            I => \N__53174\
        );

    \I__10622\ : CascadeMux
    port map (
            O => \N__53200\,
            I => \N__53171\
        );

    \I__10621\ : CascadeMux
    port map (
            O => \N__53199\,
            I => \N__53166\
        );

    \I__10620\ : CascadeMux
    port map (
            O => \N__53198\,
            I => \N__53162\
        );

    \I__10619\ : CascadeMux
    port map (
            O => \N__53197\,
            I => \N__53158\
        );

    \I__10618\ : CascadeMux
    port map (
            O => \N__53196\,
            I => \N__53155\
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__53195\,
            I => \N__53151\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__53194\,
            I => \N__53148\
        );

    \I__10615\ : InMux
    port map (
            O => \N__53191\,
            I => \N__53144\
        );

    \I__10614\ : CascadeMux
    port map (
            O => \N__53190\,
            I => \N__53141\
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__53189\,
            I => \N__53137\
        );

    \I__10612\ : Span4Mux_h
    port map (
            O => \N__53186\,
            I => \N__53131\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__53183\,
            I => \N__53131\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__53180\,
            I => \N__53127\
        );

    \I__10609\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53124\
        );

    \I__10608\ : InMux
    port map (
            O => \N__53174\,
            I => \N__53121\
        );

    \I__10607\ : InMux
    port map (
            O => \N__53171\,
            I => \N__53116\
        );

    \I__10606\ : InMux
    port map (
            O => \N__53170\,
            I => \N__53116\
        );

    \I__10605\ : InMux
    port map (
            O => \N__53169\,
            I => \N__53103\
        );

    \I__10604\ : InMux
    port map (
            O => \N__53166\,
            I => \N__53103\
        );

    \I__10603\ : InMux
    port map (
            O => \N__53165\,
            I => \N__53103\
        );

    \I__10602\ : InMux
    port map (
            O => \N__53162\,
            I => \N__53103\
        );

    \I__10601\ : InMux
    port map (
            O => \N__53161\,
            I => \N__53103\
        );

    \I__10600\ : InMux
    port map (
            O => \N__53158\,
            I => \N__53103\
        );

    \I__10599\ : InMux
    port map (
            O => \N__53155\,
            I => \N__53100\
        );

    \I__10598\ : InMux
    port map (
            O => \N__53154\,
            I => \N__53093\
        );

    \I__10597\ : InMux
    port map (
            O => \N__53151\,
            I => \N__53093\
        );

    \I__10596\ : InMux
    port map (
            O => \N__53148\,
            I => \N__53093\
        );

    \I__10595\ : InMux
    port map (
            O => \N__53147\,
            I => \N__53090\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__53144\,
            I => \N__53085\
        );

    \I__10593\ : InMux
    port map (
            O => \N__53141\,
            I => \N__53082\
        );

    \I__10592\ : CascadeMux
    port map (
            O => \N__53140\,
            I => \N__53079\
        );

    \I__10591\ : InMux
    port map (
            O => \N__53137\,
            I => \N__53076\
        );

    \I__10590\ : CascadeMux
    port map (
            O => \N__53136\,
            I => \N__53072\
        );

    \I__10589\ : Span4Mux_v
    port map (
            O => \N__53131\,
            I => \N__53069\
        );

    \I__10588\ : InMux
    port map (
            O => \N__53130\,
            I => \N__53066\
        );

    \I__10587\ : Span4Mux_h
    port map (
            O => \N__53127\,
            I => \N__53059\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__53124\,
            I => \N__53059\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__53121\,
            I => \N__53059\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__53116\,
            I => \N__53048\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__53103\,
            I => \N__53048\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__53100\,
            I => \N__53048\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__53093\,
            I => \N__53048\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__53090\,
            I => \N__53048\
        );

    \I__10579\ : InMux
    port map (
            O => \N__53089\,
            I => \N__53045\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__53088\,
            I => \N__53042\
        );

    \I__10577\ : Span4Mux_v
    port map (
            O => \N__53085\,
            I => \N__53037\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__53082\,
            I => \N__53037\
        );

    \I__10575\ : InMux
    port map (
            O => \N__53079\,
            I => \N__53034\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__53076\,
            I => \N__53031\
        );

    \I__10573\ : CascadeMux
    port map (
            O => \N__53075\,
            I => \N__53028\
        );

    \I__10572\ : InMux
    port map (
            O => \N__53072\,
            I => \N__53025\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__53069\,
            I => \N__53020\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__53066\,
            I => \N__53020\
        );

    \I__10569\ : Span4Mux_v
    port map (
            O => \N__53059\,
            I => \N__53013\
        );

    \I__10568\ : Span4Mux_v
    port map (
            O => \N__53048\,
            I => \N__53013\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__53045\,
            I => \N__53013\
        );

    \I__10566\ : InMux
    port map (
            O => \N__53042\,
            I => \N__53010\
        );

    \I__10565\ : Span4Mux_h
    port map (
            O => \N__53037\,
            I => \N__53005\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__53034\,
            I => \N__53005\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__53031\,
            I => \N__53002\
        );

    \I__10562\ : InMux
    port map (
            O => \N__53028\,
            I => \N__52999\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__53025\,
            I => \N__52996\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__53020\,
            I => \N__52989\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__53013\,
            I => \N__52989\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__53010\,
            I => \N__52989\
        );

    \I__10557\ : Span4Mux_v
    port map (
            O => \N__53005\,
            I => \N__52986\
        );

    \I__10556\ : Span4Mux_v
    port map (
            O => \N__53002\,
            I => \N__52981\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__52999\,
            I => \N__52981\
        );

    \I__10554\ : Span12Mux_h
    port map (
            O => \N__52996\,
            I => \N__52978\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__52989\,
            I => \N__52975\
        );

    \I__10552\ : Span4Mux_v
    port map (
            O => \N__52986\,
            I => \N__52970\
        );

    \I__10551\ : Span4Mux_h
    port map (
            O => \N__52981\,
            I => \N__52970\
        );

    \I__10550\ : Odrv12
    port map (
            O => \N__52978\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n126\
        );

    \I__10549\ : Odrv4
    port map (
            O => \N__52975\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n126\
        );

    \I__10548\ : Odrv4
    port map (
            O => \N__52970\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n126\
        );

    \I__10547\ : InMux
    port map (
            O => \N__52963\,
            I => \bfn_21_18_0_\
        );

    \I__10546\ : CascadeMux
    port map (
            O => \N__52960\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20596_cascade_\
        );

    \I__10545\ : CascadeMux
    port map (
            O => \N__52957\,
            I => \N__52954\
        );

    \I__10544\ : InMux
    port map (
            O => \N__52954\,
            I => \N__52951\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__52951\,
            I => \N__52948\
        );

    \I__10542\ : Span4Mux_v
    port map (
            O => \N__52948\,
            I => \N__52945\
        );

    \I__10541\ : Odrv4
    port map (
            O => \N__52945\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20604\
        );

    \I__10540\ : CascadeMux
    port map (
            O => \N__52942\,
            I => \N__52939\
        );

    \I__10539\ : InMux
    port map (
            O => \N__52939\,
            I => \N__52936\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__52936\,
            I => \N__52933\
        );

    \I__10537\ : Span4Mux_v
    port map (
            O => \N__52933\,
            I => \N__52930\
        );

    \I__10536\ : Sp12to4
    port map (
            O => \N__52930\,
            I => \N__52925\
        );

    \I__10535\ : InMux
    port map (
            O => \N__52929\,
            I => \N__52922\
        );

    \I__10534\ : InMux
    port map (
            O => \N__52928\,
            I => \N__52919\
        );

    \I__10533\ : Span12Mux_h
    port map (
            O => \N__52925\,
            I => \N__52912\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__52922\,
            I => \N__52912\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__52919\,
            I => \N__52912\
        );

    \I__10530\ : Odrv12
    port map (
            O => \N__52912\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_25\
        );

    \I__10529\ : InMux
    port map (
            O => \N__52909\,
            I => \N__52906\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__52906\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20588\
        );

    \I__10527\ : InMux
    port map (
            O => \N__52903\,
            I => \N__52900\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__52900\,
            I => \N__52897\
        );

    \I__10525\ : Span4Mux_h
    port map (
            O => \N__52897\,
            I => \N__52894\
        );

    \I__10524\ : Odrv4
    port map (
            O => \N__52894\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19896\
        );

    \I__10523\ : CascadeMux
    port map (
            O => \N__52891\,
            I => \foc.Out_31__N_333_cascade_\
        );

    \I__10522\ : InMux
    port map (
            O => \N__52888\,
            I => \N__52885\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__52885\,
            I => \N__52882\
        );

    \I__10520\ : Span4Mux_h
    port map (
            O => \N__52882\,
            I => \N__52879\
        );

    \I__10519\ : Odrv4
    port map (
            O => \N__52879\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19920\
        );

    \I__10518\ : InMux
    port map (
            O => \N__52876\,
            I => \N__52867\
        );

    \I__10517\ : InMux
    port map (
            O => \N__52875\,
            I => \N__52867\
        );

    \I__10516\ : InMux
    port map (
            O => \N__52874\,
            I => \N__52867\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__52867\,
            I => \N__52864\
        );

    \I__10514\ : Span12Mux_v
    port map (
            O => \N__52864\,
            I => \N__52861\
        );

    \I__10513\ : Odrv12
    port map (
            O => \N__52861\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_30\
        );

    \I__10512\ : CascadeMux
    port map (
            O => \N__52858\,
            I => \N__52854\
        );

    \I__10511\ : CascadeMux
    port map (
            O => \N__52857\,
            I => \N__52851\
        );

    \I__10510\ : InMux
    port map (
            O => \N__52854\,
            I => \N__52846\
        );

    \I__10509\ : InMux
    port map (
            O => \N__52851\,
            I => \N__52846\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__52846\,
            I => \N__52843\
        );

    \I__10507\ : Span4Mux_v
    port map (
            O => \N__52843\,
            I => \N__52839\
        );

    \I__10506\ : InMux
    port map (
            O => \N__52842\,
            I => \N__52836\
        );

    \I__10505\ : Sp12to4
    port map (
            O => \N__52839\,
            I => \N__52831\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__52836\,
            I => \N__52831\
        );

    \I__10503\ : Span12Mux_h
    port map (
            O => \N__52831\,
            I => \N__52828\
        );

    \I__10502\ : Odrv12
    port map (
            O => \N__52828\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_29\
        );

    \I__10501\ : InMux
    port map (
            O => \N__52825\,
            I => \N__52819\
        );

    \I__10500\ : InMux
    port map (
            O => \N__52824\,
            I => \N__52819\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__52819\,
            I => \N__52816\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__52816\,
            I => \N__52813\
        );

    \I__10497\ : Span4Mux_v
    port map (
            O => \N__52813\,
            I => \N__52810\
        );

    \I__10496\ : Span4Mux_v
    port map (
            O => \N__52810\,
            I => \N__52807\
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__52807\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Voltage_1_31\
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__52804\,
            I => \foc.Out_31__N_332_cascade_\
        );

    \I__10493\ : InMux
    port map (
            O => \N__52801\,
            I => \N__52798\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__52798\,
            I => \foc.qVoltage_9\
        );

    \I__10491\ : InMux
    port map (
            O => \N__52795\,
            I => \N__52789\
        );

    \I__10490\ : InMux
    port map (
            O => \N__52794\,
            I => \N__52789\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__52789\,
            I => \N__52786\
        );

    \I__10488\ : Span4Mux_h
    port map (
            O => \N__52786\,
            I => \N__52782\
        );

    \I__10487\ : InMux
    port map (
            O => \N__52785\,
            I => \N__52779\
        );

    \I__10486\ : Span4Mux_v
    port map (
            O => \N__52782\,
            I => \N__52776\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__52779\,
            I => \N__52773\
        );

    \I__10484\ : Sp12to4
    port map (
            O => \N__52776\,
            I => \N__52767\
        );

    \I__10483\ : Span12Mux_h
    port map (
            O => \N__52773\,
            I => \N__52767\
        );

    \I__10482\ : InMux
    port map (
            O => \N__52772\,
            I => \N__52764\
        );

    \I__10481\ : Odrv12
    port map (
            O => \N__52767\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__52764\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18\
        );

    \I__10479\ : CascadeMux
    port map (
            O => \N__52759\,
            I => \foc.qVoltage_14_cascade_\
        );

    \I__10478\ : InMux
    port map (
            O => \N__52756\,
            I => \N__52750\
        );

    \I__10477\ : InMux
    port map (
            O => \N__52755\,
            I => \N__52750\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__52750\,
            I => \N__52747\
        );

    \I__10475\ : Span4Mux_h
    port map (
            O => \N__52747\,
            I => \N__52742\
        );

    \I__10474\ : InMux
    port map (
            O => \N__52746\,
            I => \N__52739\
        );

    \I__10473\ : InMux
    port map (
            O => \N__52745\,
            I => \N__52736\
        );

    \I__10472\ : Sp12to4
    port map (
            O => \N__52742\,
            I => \N__52729\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__52739\,
            I => \N__52729\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__52736\,
            I => \N__52729\
        );

    \I__10469\ : Odrv12
    port map (
            O => \N__52729\,
            I => \foc.preSatVoltage_23\
        );

    \I__10468\ : InMux
    port map (
            O => \N__52726\,
            I => \N__52723\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__52723\,
            I => \N__52719\
        );

    \I__10466\ : InMux
    port map (
            O => \N__52722\,
            I => \N__52716\
        );

    \I__10465\ : Span4Mux_v
    port map (
            O => \N__52719\,
            I => \N__52713\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__52716\,
            I => \N__52710\
        );

    \I__10463\ : Span4Mux_h
    port map (
            O => \N__52713\,
            I => \N__52705\
        );

    \I__10462\ : Span4Mux_v
    port map (
            O => \N__52710\,
            I => \N__52705\
        );

    \I__10461\ : Span4Mux_h
    port map (
            O => \N__52705\,
            I => \N__52700\
        );

    \I__10460\ : InMux
    port map (
            O => \N__52704\,
            I => \N__52697\
        );

    \I__10459\ : InMux
    port map (
            O => \N__52703\,
            I => \N__52694\
        );

    \I__10458\ : Sp12to4
    port map (
            O => \N__52700\,
            I => \N__52687\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__52697\,
            I => \N__52687\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__52694\,
            I => \N__52687\
        );

    \I__10455\ : Odrv12
    port map (
            O => \N__52687\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_24\
        );

    \I__10454\ : InMux
    port map (
            O => \N__52684\,
            I => \N__52681\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__52681\,
            I => \foc.qVoltage_15\
        );

    \I__10452\ : CascadeMux
    port map (
            O => \N__52678\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20548_cascade_\
        );

    \I__10451\ : InMux
    port map (
            O => \N__52675\,
            I => \N__52672\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__52672\,
            I => \foc.dVoltage_15\
        );

    \I__10449\ : CascadeMux
    port map (
            O => \N__52669\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20562_cascade_\
        );

    \I__10448\ : InMux
    port map (
            O => \N__52666\,
            I => \N__52663\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__52663\,
            I => \foc.dVoltage_10\
        );

    \I__10446\ : CascadeMux
    port map (
            O => \N__52660\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20574_cascade_\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__52657\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19727_cascade_\
        );

    \I__10444\ : CascadeMux
    port map (
            O => \N__52654\,
            I => \foc.qVoltage_5_cascade_\
        );

    \I__10443\ : InMux
    port map (
            O => \N__52651\,
            I => \N__52645\
        );

    \I__10442\ : InMux
    port map (
            O => \N__52650\,
            I => \N__52645\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__52645\,
            I => \N__52642\
        );

    \I__10440\ : Span12Mux_v
    port map (
            O => \N__52642\,
            I => \N__52637\
        );

    \I__10439\ : InMux
    port map (
            O => \N__52641\,
            I => \N__52634\
        );

    \I__10438\ : InMux
    port map (
            O => \N__52640\,
            I => \N__52631\
        );

    \I__10437\ : Odrv12
    port map (
            O => \N__52637\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14\
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__52634\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__52631\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14\
        );

    \I__10434\ : InMux
    port map (
            O => \N__52624\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17560\
        );

    \I__10433\ : CascadeMux
    port map (
            O => \N__52621\,
            I => \N__52618\
        );

    \I__10432\ : InMux
    port map (
            O => \N__52618\,
            I => \N__52615\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__52615\,
            I => \N__52612\
        );

    \I__10430\ : Odrv12
    port map (
            O => \N__52612\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n550_adj_441\
        );

    \I__10429\ : InMux
    port map (
            O => \N__52609\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17561\
        );

    \I__10428\ : InMux
    port map (
            O => \N__52606\,
            I => \N__52603\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52600\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__52600\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n599_adj_376\
        );

    \I__10425\ : InMux
    port map (
            O => \N__52597\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17562\
        );

    \I__10424\ : CascadeMux
    port map (
            O => \N__52594\,
            I => \N__52591\
        );

    \I__10423\ : InMux
    port map (
            O => \N__52591\,
            I => \N__52588\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__52588\,
            I => \N__52585\
        );

    \I__10421\ : Odrv4
    port map (
            O => \N__52585\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n648\
        );

    \I__10420\ : InMux
    port map (
            O => \N__52582\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17563\
        );

    \I__10419\ : InMux
    port map (
            O => \N__52579\,
            I => \N__52576\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__52576\,
            I => \N__52573\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__52573\,
            I => \N__52569\
        );

    \I__10416\ : InMux
    port map (
            O => \N__52572\,
            I => \N__52566\
        );

    \I__10415\ : Span4Mux_v
    port map (
            O => \N__52569\,
            I => \N__52561\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__52566\,
            I => \N__52561\
        );

    \I__10413\ : Odrv4
    port map (
            O => \N__52561\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n745\
        );

    \I__10412\ : CascadeMux
    port map (
            O => \N__52558\,
            I => \N__52555\
        );

    \I__10411\ : InMux
    port map (
            O => \N__52555\,
            I => \N__52552\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__52552\,
            I => \N__52549\
        );

    \I__10409\ : Odrv4
    port map (
            O => \N__52549\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n697_adj_444\
        );

    \I__10408\ : CascadeMux
    port map (
            O => \N__52546\,
            I => \N__52543\
        );

    \I__10407\ : InMux
    port map (
            O => \N__52543\,
            I => \N__52540\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__52540\,
            I => \N__52537\
        );

    \I__10405\ : Odrv4
    port map (
            O => \N__52537\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n746_adj_409\
        );

    \I__10404\ : InMux
    port map (
            O => \N__52534\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17564\
        );

    \I__10403\ : InMux
    port map (
            O => \N__52531\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408\
        );

    \I__10402\ : CascadeMux
    port map (
            O => \N__52528\,
            I => \N__52525\
        );

    \I__10401\ : InMux
    port map (
            O => \N__52525\,
            I => \N__52522\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__52522\,
            I => \N__52519\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__52519\,
            I => \N__52516\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__52516\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_CO\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__52513\,
            I => \foc.dVoltage_2_cascade_\
        );

    \I__10396\ : InMux
    port map (
            O => \N__52510\,
            I => \N__52507\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__52507\,
            I => \N__52504\
        );

    \I__10394\ : Odrv4
    port map (
            O => \N__52504\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n109\
        );

    \I__10393\ : InMux
    port map (
            O => \N__52501\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17552\
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__52498\,
            I => \N__52495\
        );

    \I__10391\ : InMux
    port map (
            O => \N__52495\,
            I => \N__52492\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__52492\,
            I => \N__52489\
        );

    \I__10389\ : Odrv12
    port map (
            O => \N__52489\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n158\
        );

    \I__10388\ : InMux
    port map (
            O => \N__52486\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17553\
        );

    \I__10387\ : InMux
    port map (
            O => \N__52483\,
            I => \N__52480\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__52480\,
            I => \N__52477\
        );

    \I__10385\ : Odrv4
    port map (
            O => \N__52477\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n207_adj_394\
        );

    \I__10384\ : InMux
    port map (
            O => \N__52474\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17554\
        );

    \I__10383\ : CascadeMux
    port map (
            O => \N__52471\,
            I => \N__52468\
        );

    \I__10382\ : InMux
    port map (
            O => \N__52468\,
            I => \N__52465\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__52465\,
            I => \N__52462\
        );

    \I__10380\ : Odrv4
    port map (
            O => \N__52462\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n256_adj_392\
        );

    \I__10379\ : InMux
    port map (
            O => \N__52459\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17555\
        );

    \I__10378\ : InMux
    port map (
            O => \N__52456\,
            I => \N__52453\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__52453\,
            I => \N__52450\
        );

    \I__10376\ : Odrv12
    port map (
            O => \N__52450\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n305_adj_390\
        );

    \I__10375\ : InMux
    port map (
            O => \N__52447\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17556\
        );

    \I__10374\ : CascadeMux
    port map (
            O => \N__52444\,
            I => \N__52441\
        );

    \I__10373\ : InMux
    port map (
            O => \N__52441\,
            I => \N__52438\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__52438\,
            I => \N__52435\
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__52435\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n354\
        );

    \I__10370\ : InMux
    port map (
            O => \N__52432\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17557\
        );

    \I__10369\ : InMux
    port map (
            O => \N__52429\,
            I => \N__52426\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__52426\,
            I => \N__52423\
        );

    \I__10367\ : Odrv12
    port map (
            O => \N__52423\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n403\
        );

    \I__10366\ : InMux
    port map (
            O => \N__52420\,
            I => \bfn_21_12_0_\
        );

    \I__10365\ : CascadeMux
    port map (
            O => \N__52417\,
            I => \N__52414\
        );

    \I__10364\ : InMux
    port map (
            O => \N__52414\,
            I => \N__52411\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__52411\,
            I => \N__52408\
        );

    \I__10362\ : Odrv12
    port map (
            O => \N__52408\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n452\
        );

    \I__10361\ : InMux
    port map (
            O => \N__52405\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17559\
        );

    \I__10360\ : InMux
    port map (
            O => \N__52402\,
            I => \N__52399\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__52399\,
            I => \N__52396\
        );

    \I__10358\ : Odrv4
    port map (
            O => \N__52396\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n501_adj_481\
        );

    \I__10357\ : InMux
    port map (
            O => \N__52393\,
            I => \N__52390\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__52390\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n504_adj_467\
        );

    \I__10355\ : InMux
    port map (
            O => \N__52387\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17575\
        );

    \I__10354\ : CascadeMux
    port map (
            O => \N__52384\,
            I => \N__52381\
        );

    \I__10353\ : InMux
    port map (
            O => \N__52381\,
            I => \N__52378\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__52378\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n553_adj_446\
        );

    \I__10351\ : InMux
    port map (
            O => \N__52375\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17576\
        );

    \I__10350\ : InMux
    port map (
            O => \N__52372\,
            I => \N__52369\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__52369\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n602_adj_355\
        );

    \I__10348\ : InMux
    port map (
            O => \N__52366\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17577\
        );

    \I__10347\ : CascadeMux
    port map (
            O => \N__52363\,
            I => \N__52360\
        );

    \I__10346\ : InMux
    port map (
            O => \N__52360\,
            I => \N__52357\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__52357\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n651\
        );

    \I__10344\ : InMux
    port map (
            O => \N__52354\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17578\
        );

    \I__10343\ : InMux
    port map (
            O => \N__52351\,
            I => \N__52348\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__52348\,
            I => \N__52345\
        );

    \I__10341\ : Span4Mux_v
    port map (
            O => \N__52345\,
            I => \N__52341\
        );

    \I__10340\ : InMux
    port map (
            O => \N__52344\,
            I => \N__52338\
        );

    \I__10339\ : Odrv4
    port map (
            O => \N__52341\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n749\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__52338\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n749\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__52333\,
            I => \N__52330\
        );

    \I__10336\ : InMux
    port map (
            O => \N__52330\,
            I => \N__52327\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__52327\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n700\
        );

    \I__10334\ : InMux
    port map (
            O => \N__52324\,
            I => \N__52321\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__52321\,
            I => \N__52318\
        );

    \I__10332\ : Span4Mux_v
    port map (
            O => \N__52318\,
            I => \N__52315\
        );

    \I__10331\ : Odrv4
    port map (
            O => \N__52315\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n750_adj_407\
        );

    \I__10330\ : InMux
    port map (
            O => \N__52312\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17579\
        );

    \I__10329\ : InMux
    port map (
            O => \N__52309\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406\
        );

    \I__10328\ : CascadeMux
    port map (
            O => \N__52306\,
            I => \N__52303\
        );

    \I__10327\ : InMux
    port map (
            O => \N__52303\,
            I => \N__52300\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__52300\,
            I => \N__52297\
        );

    \I__10325\ : Span4Mux_v
    port map (
            O => \N__52297\,
            I => \N__52294\
        );

    \I__10324\ : Odrv4
    port map (
            O => \N__52294\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_CO\
        );

    \I__10323\ : CascadeMux
    port map (
            O => \N__52291\,
            I => \N__52288\
        );

    \I__10322\ : InMux
    port map (
            O => \N__52288\,
            I => \N__52285\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__52285\,
            I => \N__52282\
        );

    \I__10320\ : Odrv4
    port map (
            O => \N__52282\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n60_adj_495\
        );

    \I__10319\ : InMux
    port map (
            O => \N__52279\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17551\
        );

    \I__10318\ : CascadeMux
    port map (
            O => \N__52276\,
            I => \N__52273\
        );

    \I__10317\ : InMux
    port map (
            O => \N__52273\,
            I => \N__52270\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__52270\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n63\
        );

    \I__10315\ : InMux
    port map (
            O => \N__52267\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17566\
        );

    \I__10314\ : InMux
    port map (
            O => \N__52264\,
            I => \N__52261\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__52261\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n112_adj_442\
        );

    \I__10312\ : InMux
    port map (
            O => \N__52258\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17567\
        );

    \I__10311\ : InMux
    port map (
            O => \N__52255\,
            I => \N__52252\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__52252\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n161_adj_395\
        );

    \I__10309\ : InMux
    port map (
            O => \N__52249\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17568\
        );

    \I__10308\ : InMux
    port map (
            O => \N__52246\,
            I => \N__52243\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__52243\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n210_adj_393\
        );

    \I__10306\ : InMux
    port map (
            O => \N__52240\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17569\
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__52237\,
            I => \N__52234\
        );

    \I__10304\ : InMux
    port map (
            O => \N__52234\,
            I => \N__52231\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__52231\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n259_adj_391\
        );

    \I__10302\ : InMux
    port map (
            O => \N__52228\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17570\
        );

    \I__10301\ : InMux
    port map (
            O => \N__52225\,
            I => \N__52222\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__52222\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n308\
        );

    \I__10299\ : InMux
    port map (
            O => \N__52219\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17571\
        );

    \I__10298\ : CascadeMux
    port map (
            O => \N__52216\,
            I => \N__52213\
        );

    \I__10297\ : InMux
    port map (
            O => \N__52213\,
            I => \N__52210\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__52210\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n357\
        );

    \I__10295\ : InMux
    port map (
            O => \N__52207\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17572\
        );

    \I__10294\ : InMux
    port map (
            O => \N__52204\,
            I => \N__52201\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__52201\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n406\
        );

    \I__10292\ : InMux
    port map (
            O => \N__52198\,
            I => \bfn_21_10_0_\
        );

    \I__10291\ : CascadeMux
    port map (
            O => \N__52195\,
            I => \N__52192\
        );

    \I__10290\ : InMux
    port map (
            O => \N__52192\,
            I => \N__52189\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__52189\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n455\
        );

    \I__10288\ : InMux
    port map (
            O => \N__52186\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17574\
        );

    \I__10287\ : CascadeMux
    port map (
            O => \N__52183\,
            I => \N__52180\
        );

    \I__10286\ : InMux
    port map (
            O => \N__52180\,
            I => \N__52177\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__52177\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n461_adj_470\
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__52174\,
            I => \N__52171\
        );

    \I__10283\ : InMux
    port map (
            O => \N__52171\,
            I => \N__52168\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__52168\,
            I => \N__52165\
        );

    \I__10281\ : Odrv4
    port map (
            O => \N__52165\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n507_adj_447\
        );

    \I__10280\ : InMux
    port map (
            O => \N__52162\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17604\
        );

    \I__10279\ : InMux
    port map (
            O => \N__52159\,
            I => \N__52156\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__52156\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n510_adj_458\
        );

    \I__10277\ : InMux
    port map (
            O => \N__52153\,
            I => \N__52150\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__52150\,
            I => \N__52147\
        );

    \I__10275\ : Odrv4
    port map (
            O => \N__52147\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n556\
        );

    \I__10274\ : InMux
    port map (
            O => \N__52144\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17605\
        );

    \I__10273\ : CascadeMux
    port map (
            O => \N__52141\,
            I => \N__52138\
        );

    \I__10272\ : InMux
    port map (
            O => \N__52138\,
            I => \N__52135\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__52135\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n559\
        );

    \I__10270\ : CascadeMux
    port map (
            O => \N__52132\,
            I => \N__52129\
        );

    \I__10269\ : InMux
    port map (
            O => \N__52129\,
            I => \N__52126\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__52126\,
            I => \N__52123\
        );

    \I__10267\ : Odrv4
    port map (
            O => \N__52123\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n605\
        );

    \I__10266\ : InMux
    port map (
            O => \N__52120\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17606\
        );

    \I__10265\ : InMux
    port map (
            O => \N__52117\,
            I => \N__52114\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__52114\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n608\
        );

    \I__10263\ : InMux
    port map (
            O => \N__52111\,
            I => \N__52108\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__52108\,
            I => \N__52105\
        );

    \I__10261\ : Span4Mux_v
    port map (
            O => \N__52105\,
            I => \N__52102\
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__52102\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n654\
        );

    \I__10259\ : InMux
    port map (
            O => \N__52099\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17607\
        );

    \I__10258\ : CascadeMux
    port map (
            O => \N__52096\,
            I => \N__52093\
        );

    \I__10257\ : InMux
    port map (
            O => \N__52093\,
            I => \N__52090\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__52090\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n657\
        );

    \I__10255\ : CascadeMux
    port map (
            O => \N__52087\,
            I => \N__52084\
        );

    \I__10254\ : InMux
    port map (
            O => \N__52084\,
            I => \N__52081\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__52081\,
            I => \N__52078\
        );

    \I__10252\ : Sp12to4
    port map (
            O => \N__52078\,
            I => \N__52075\
        );

    \I__10251\ : Odrv12
    port map (
            O => \N__52075\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n703\
        );

    \I__10250\ : InMux
    port map (
            O => \N__52072\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17608\
        );

    \I__10249\ : InMux
    port map (
            O => \N__52069\,
            I => \N__52066\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__52066\,
            I => \N__52063\
        );

    \I__10247\ : Span4Mux_h
    port map (
            O => \N__52063\,
            I => \N__52059\
        );

    \I__10246\ : InMux
    port map (
            O => \N__52062\,
            I => \N__52056\
        );

    \I__10245\ : Odrv4
    port map (
            O => \N__52059\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n757\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__52056\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n757\
        );

    \I__10243\ : CascadeMux
    port map (
            O => \N__52051\,
            I => \N__52048\
        );

    \I__10242\ : InMux
    port map (
            O => \N__52048\,
            I => \N__52045\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__52045\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n706\
        );

    \I__10240\ : InMux
    port map (
            O => \N__52042\,
            I => \N__52039\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__52039\,
            I => \N__52036\
        );

    \I__10238\ : Span4Mux_v
    port map (
            O => \N__52036\,
            I => \N__52033\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__52033\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n758_adj_403\
        );

    \I__10236\ : InMux
    port map (
            O => \N__52030\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17609\
        );

    \I__10235\ : InMux
    port map (
            O => \N__52027\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n759\
        );

    \I__10234\ : CascadeMux
    port map (
            O => \N__52024\,
            I => \N__52021\
        );

    \I__10233\ : InMux
    port map (
            O => \N__52021\,
            I => \N__52018\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__52018\,
            I => \N__52015\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__52015\,
            I => \N__52012\
        );

    \I__10230\ : Odrv4
    port map (
            O => \N__52012\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_CO\
        );

    \I__10229\ : InMux
    port map (
            O => \N__52009\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17596\
        );

    \I__10228\ : CascadeMux
    port map (
            O => \N__52006\,
            I => \N__52003\
        );

    \I__10227\ : InMux
    port map (
            O => \N__52003\,
            I => \N__52000\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__52000\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n118_adj_487\
        );

    \I__10225\ : InMux
    port map (
            O => \N__51997\,
            I => \N__51994\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__51994\,
            I => \N__51991\
        );

    \I__10223\ : Odrv4
    port map (
            O => \N__51991\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n164_adj_466\
        );

    \I__10222\ : InMux
    port map (
            O => \N__51988\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17597\
        );

    \I__10221\ : InMux
    port map (
            O => \N__51985\,
            I => \N__51982\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__51982\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n167_adj_486\
        );

    \I__10219\ : CascadeMux
    port map (
            O => \N__51979\,
            I => \N__51976\
        );

    \I__10218\ : InMux
    port map (
            O => \N__51976\,
            I => \N__51973\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__51973\,
            I => \N__51970\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__51970\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n213_adj_445\
        );

    \I__10215\ : InMux
    port map (
            O => \N__51967\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17598\
        );

    \I__10214\ : InMux
    port map (
            O => \N__51964\,
            I => \N__51961\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__51961\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n216_adj_485\
        );

    \I__10212\ : CascadeMux
    port map (
            O => \N__51958\,
            I => \N__51955\
        );

    \I__10211\ : InMux
    port map (
            O => \N__51955\,
            I => \N__51952\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__51952\,
            I => \N__51949\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__51949\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n262\
        );

    \I__10208\ : InMux
    port map (
            O => \N__51946\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17599\
        );

    \I__10207\ : InMux
    port map (
            O => \N__51943\,
            I => \N__51940\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__51940\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n265_adj_471\
        );

    \I__10205\ : InMux
    port map (
            O => \N__51937\,
            I => \N__51934\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__51934\,
            I => \N__51931\
        );

    \I__10203\ : Odrv4
    port map (
            O => \N__51931\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n311\
        );

    \I__10202\ : InMux
    port map (
            O => \N__51928\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17600\
        );

    \I__10201\ : InMux
    port map (
            O => \N__51925\,
            I => \N__51922\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__51922\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n314\
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__51919\,
            I => \N__51916\
        );

    \I__10198\ : InMux
    port map (
            O => \N__51916\,
            I => \N__51913\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__51913\,
            I => \N__51910\
        );

    \I__10196\ : Odrv4
    port map (
            O => \N__51910\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n360_adj_484\
        );

    \I__10195\ : InMux
    port map (
            O => \N__51907\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17601\
        );

    \I__10194\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51901\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__51901\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n363\
        );

    \I__10192\ : InMux
    port map (
            O => \N__51898\,
            I => \N__51895\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__51895\,
            I => \N__51892\
        );

    \I__10190\ : Odrv4
    port map (
            O => \N__51892\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n409_adj_483\
        );

    \I__10189\ : InMux
    port map (
            O => \N__51889\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17602\
        );

    \I__10188\ : InMux
    port map (
            O => \N__51886\,
            I => \N__51883\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__51883\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n412_adj_482\
        );

    \I__10186\ : InMux
    port map (
            O => \N__51880\,
            I => \N__51877\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__51877\,
            I => \N__51874\
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__51874\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n458_adj_468\
        );

    \I__10183\ : InMux
    port map (
            O => \N__51871\,
            I => \bfn_21_8_0_\
        );

    \I__10182\ : InMux
    port map (
            O => \N__51868\,
            I => \N__51865\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__51865\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n476\
        );

    \I__10180\ : InMux
    port map (
            O => \N__51862\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18317\
        );

    \I__10179\ : InMux
    port map (
            O => \N__51859\,
            I => \N__51856\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__51856\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n525\
        );

    \I__10177\ : InMux
    port map (
            O => \N__51853\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18318\
        );

    \I__10176\ : InMux
    port map (
            O => \N__51850\,
            I => \N__51847\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__51847\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n574\
        );

    \I__10174\ : InMux
    port map (
            O => \N__51844\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18319\
        );

    \I__10173\ : InMux
    port map (
            O => \N__51841\,
            I => \N__51838\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__51838\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n623\
        );

    \I__10171\ : InMux
    port map (
            O => \N__51835\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18320\
        );

    \I__10170\ : CascadeMux
    port map (
            O => \N__51832\,
            I => \N__51829\
        );

    \I__10169\ : InMux
    port map (
            O => \N__51829\,
            I => \N__51826\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__51826\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n672\
        );

    \I__10167\ : InMux
    port map (
            O => \N__51823\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18321\
        );

    \I__10166\ : CascadeMux
    port map (
            O => \N__51820\,
            I => \N__51817\
        );

    \I__10165\ : InMux
    port map (
            O => \N__51817\,
            I => \N__51814\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__51814\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n721\
        );

    \I__10163\ : InMux
    port map (
            O => \N__51811\,
            I => \N__51808\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__51808\,
            I => \N__51805\
        );

    \I__10161\ : Span4Mux_v
    port map (
            O => \N__51805\,
            I => \N__51802\
        );

    \I__10160\ : Sp12to4
    port map (
            O => \N__51802\,
            I => \N__51799\
        );

    \I__10159\ : Odrv12
    port map (
            O => \N__51799\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n778\
        );

    \I__10158\ : InMux
    port map (
            O => \N__51796\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18322\
        );

    \I__10157\ : InMux
    port map (
            O => \N__51793\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779\
        );

    \I__10156\ : CascadeMux
    port map (
            O => \N__51790\,
            I => \N__51787\
        );

    \I__10155\ : InMux
    port map (
            O => \N__51787\,
            I => \N__51784\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__51784\,
            I => \N__51781\
        );

    \I__10153\ : Span4Mux_h
    port map (
            O => \N__51781\,
            I => \N__51778\
        );

    \I__10152\ : Span4Mux_v
    port map (
            O => \N__51778\,
            I => \N__51775\
        );

    \I__10151\ : Odrv4
    port map (
            O => \N__51775\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_CO\
        );

    \I__10150\ : InMux
    port map (
            O => \N__51772\,
            I => \N__51769\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__51769\,
            I => \N__51766\
        );

    \I__10148\ : Odrv4
    port map (
            O => \N__51766\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n66\
        );

    \I__10147\ : CascadeMux
    port map (
            O => \N__51763\,
            I => \N__51760\
        );

    \I__10146\ : InMux
    port map (
            O => \N__51760\,
            I => \N__51757\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__51757\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n69_adj_489\
        );

    \I__10144\ : CascadeMux
    port map (
            O => \N__51754\,
            I => \N__51751\
        );

    \I__10143\ : InMux
    port map (
            O => \N__51751\,
            I => \N__51748\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__51748\,
            I => \N__51745\
        );

    \I__10141\ : Odrv4
    port map (
            O => \N__51745\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n115_adj_488\
        );

    \I__10140\ : InMux
    port map (
            O => \N__51742\,
            I => \N__51739\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__51739\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n84\
        );

    \I__10138\ : InMux
    port map (
            O => \N__51736\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18309\
        );

    \I__10137\ : InMux
    port map (
            O => \N__51733\,
            I => \N__51730\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__51730\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n133\
        );

    \I__10135\ : InMux
    port map (
            O => \N__51727\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18310\
        );

    \I__10134\ : InMux
    port map (
            O => \N__51724\,
            I => \N__51721\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__51721\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n182\
        );

    \I__10132\ : InMux
    port map (
            O => \N__51718\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18311\
        );

    \I__10131\ : InMux
    port map (
            O => \N__51715\,
            I => \N__51712\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__51712\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n231\
        );

    \I__10129\ : InMux
    port map (
            O => \N__51709\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18312\
        );

    \I__10128\ : InMux
    port map (
            O => \N__51706\,
            I => \N__51703\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__51703\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n280\
        );

    \I__10126\ : InMux
    port map (
            O => \N__51700\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18313\
        );

    \I__10125\ : InMux
    port map (
            O => \N__51697\,
            I => \N__51694\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__51694\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n329\
        );

    \I__10123\ : InMux
    port map (
            O => \N__51691\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18314\
        );

    \I__10122\ : InMux
    port map (
            O => \N__51688\,
            I => \N__51685\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__51685\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n378\
        );

    \I__10120\ : InMux
    port map (
            O => \N__51682\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18315\
        );

    \I__10119\ : InMux
    port map (
            O => \N__51679\,
            I => \N__51676\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__51676\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n427\
        );

    \I__10117\ : InMux
    port map (
            O => \N__51673\,
            I => \bfn_20_29_0_\
        );

    \I__10116\ : InMux
    port map (
            O => \N__51670\,
            I => \N__51667\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__51667\,
            I => \N__51664\
        );

    \I__10114\ : Odrv4
    port map (
            O => \N__51664\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n455\
        );

    \I__10113\ : InMux
    port map (
            O => \N__51661\,
            I => \bfn_20_26_0_\
        );

    \I__10112\ : InMux
    port map (
            O => \N__51658\,
            I => \N__51655\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__51655\,
            I => \N__51652\
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__51652\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n504\
        );

    \I__10109\ : InMux
    port map (
            O => \N__51649\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18227\
        );

    \I__10108\ : InMux
    port map (
            O => \N__51646\,
            I => \N__51643\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__51643\,
            I => \N__51640\
        );

    \I__10106\ : Odrv12
    port map (
            O => \N__51640\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n553\
        );

    \I__10105\ : InMux
    port map (
            O => \N__51637\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18228\
        );

    \I__10104\ : CascadeMux
    port map (
            O => \N__51634\,
            I => \N__51631\
        );

    \I__10103\ : InMux
    port map (
            O => \N__51631\,
            I => \N__51628\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__51628\,
            I => \N__51625\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__51625\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n602\
        );

    \I__10100\ : InMux
    port map (
            O => \N__51622\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18229\
        );

    \I__10099\ : CascadeMux
    port map (
            O => \N__51619\,
            I => \N__51616\
        );

    \I__10098\ : InMux
    port map (
            O => \N__51616\,
            I => \N__51613\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__51613\,
            I => \N__51610\
        );

    \I__10096\ : Span4Mux_h
    port map (
            O => \N__51610\,
            I => \N__51607\
        );

    \I__10095\ : Odrv4
    port map (
            O => \N__51607\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n651\
        );

    \I__10094\ : InMux
    port map (
            O => \N__51604\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18230\
        );

    \I__10093\ : CascadeMux
    port map (
            O => \N__51601\,
            I => \N__51598\
        );

    \I__10092\ : InMux
    port map (
            O => \N__51598\,
            I => \N__51595\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__51595\,
            I => \N__51592\
        );

    \I__10090\ : Odrv4
    port map (
            O => \N__51592\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n700\
        );

    \I__10089\ : InMux
    port map (
            O => \N__51589\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18231\
        );

    \I__10088\ : InMux
    port map (
            O => \N__51586\,
            I => \N__51583\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__51583\,
            I => \N__51580\
        );

    \I__10086\ : Span4Mux_v
    port map (
            O => \N__51580\,
            I => \N__51577\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__51577\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n754\
        );

    \I__10084\ : InMux
    port map (
            O => \N__51574\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18232\
        );

    \I__10083\ : InMux
    port map (
            O => \N__51571\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755\
        );

    \I__10082\ : CascadeMux
    port map (
            O => \N__51568\,
            I => \N__51565\
        );

    \I__10081\ : InMux
    port map (
            O => \N__51565\,
            I => \N__51562\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__51562\,
            I => \N__51559\
        );

    \I__10079\ : Span4Mux_v
    port map (
            O => \N__51559\,
            I => \N__51556\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__51556\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_CO\
        );

    \I__10077\ : CascadeMux
    port map (
            O => \N__51553\,
            I => \N__51550\
        );

    \I__10076\ : InMux
    port map (
            O => \N__51550\,
            I => \N__51547\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__51547\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n66\
        );

    \I__10074\ : InMux
    port map (
            O => \N__51544\,
            I => \N__51541\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__51541\,
            I => \N__51538\
        );

    \I__10072\ : Odrv4
    port map (
            O => \N__51538\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n112\
        );

    \I__10071\ : InMux
    port map (
            O => \N__51535\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18219\
        );

    \I__10070\ : InMux
    port map (
            O => \N__51532\,
            I => \N__51529\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__51529\,
            I => \N__51526\
        );

    \I__10068\ : Odrv4
    port map (
            O => \N__51526\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n161\
        );

    \I__10067\ : InMux
    port map (
            O => \N__51523\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18220\
        );

    \I__10066\ : InMux
    port map (
            O => \N__51520\,
            I => \N__51517\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__51517\,
            I => \N__51514\
        );

    \I__10064\ : Odrv4
    port map (
            O => \N__51514\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n210\
        );

    \I__10063\ : InMux
    port map (
            O => \N__51511\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18221\
        );

    \I__10062\ : InMux
    port map (
            O => \N__51508\,
            I => \N__51505\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__51505\,
            I => \N__51502\
        );

    \I__10060\ : Odrv4
    port map (
            O => \N__51502\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n259\
        );

    \I__10059\ : InMux
    port map (
            O => \N__51499\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18222\
        );

    \I__10058\ : CascadeMux
    port map (
            O => \N__51496\,
            I => \N__51493\
        );

    \I__10057\ : InMux
    port map (
            O => \N__51493\,
            I => \N__51490\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__51490\,
            I => \N__51487\
        );

    \I__10055\ : Odrv4
    port map (
            O => \N__51487\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n308\
        );

    \I__10054\ : InMux
    port map (
            O => \N__51484\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18223\
        );

    \I__10053\ : CascadeMux
    port map (
            O => \N__51481\,
            I => \N__51478\
        );

    \I__10052\ : InMux
    port map (
            O => \N__51478\,
            I => \N__51475\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__51475\,
            I => \N__51472\
        );

    \I__10050\ : Odrv12
    port map (
            O => \N__51472\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n357\
        );

    \I__10049\ : InMux
    port map (
            O => \N__51469\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18224\
        );

    \I__10048\ : InMux
    port map (
            O => \N__51466\,
            I => \N__51463\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__51463\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n406\
        );

    \I__10046\ : InMux
    port map (
            O => \N__51460\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18225\
        );

    \I__10045\ : InMux
    port map (
            O => \N__51457\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18210\
        );

    \I__10044\ : InMux
    port map (
            O => \N__51454\,
            I => \N__51451\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__51451\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n452\
        );

    \I__10042\ : InMux
    port map (
            O => \N__51448\,
            I => \bfn_20_24_0_\
        );

    \I__10041\ : InMux
    port map (
            O => \N__51445\,
            I => \N__51442\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__51442\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n501\
        );

    \I__10039\ : InMux
    port map (
            O => \N__51439\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18212\
        );

    \I__10038\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51433\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__51433\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n550\
        );

    \I__10036\ : InMux
    port map (
            O => \N__51430\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18213\
        );

    \I__10035\ : InMux
    port map (
            O => \N__51427\,
            I => \N__51424\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__51424\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n599\
        );

    \I__10033\ : InMux
    port map (
            O => \N__51421\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18214\
        );

    \I__10032\ : CascadeMux
    port map (
            O => \N__51418\,
            I => \N__51415\
        );

    \I__10031\ : InMux
    port map (
            O => \N__51415\,
            I => \N__51412\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__51412\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n648\
        );

    \I__10029\ : InMux
    port map (
            O => \N__51409\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18215\
        );

    \I__10028\ : CascadeMux
    port map (
            O => \N__51406\,
            I => \N__51403\
        );

    \I__10027\ : InMux
    port map (
            O => \N__51403\,
            I => \N__51400\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__51400\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n697\
        );

    \I__10025\ : InMux
    port map (
            O => \N__51397\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18216\
        );

    \I__10024\ : InMux
    port map (
            O => \N__51394\,
            I => \N__51391\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__51391\,
            I => \N__51388\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__51388\,
            I => \N__51385\
        );

    \I__10021\ : Odrv4
    port map (
            O => \N__51385\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n750\
        );

    \I__10020\ : InMux
    port map (
            O => \N__51382\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18217\
        );

    \I__10019\ : InMux
    port map (
            O => \N__51379\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751\
        );

    \I__10018\ : CascadeMux
    port map (
            O => \N__51376\,
            I => \N__51373\
        );

    \I__10017\ : InMux
    port map (
            O => \N__51373\,
            I => \N__51370\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__51370\,
            I => \N__51367\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__51367\,
            I => \N__51364\
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__51364\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_CO\
        );

    \I__10013\ : CascadeMux
    port map (
            O => \N__51361\,
            I => \N__51358\
        );

    \I__10012\ : InMux
    port map (
            O => \N__51358\,
            I => \N__51355\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__51355\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n63\
        );

    \I__10010\ : CascadeMux
    port map (
            O => \N__51352\,
            I => \N__51349\
        );

    \I__10009\ : InMux
    port map (
            O => \N__51349\,
            I => \N__51346\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__51346\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n109\
        );

    \I__10007\ : InMux
    port map (
            O => \N__51343\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18204\
        );

    \I__10006\ : InMux
    port map (
            O => \N__51340\,
            I => \N__51337\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__51337\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n158\
        );

    \I__10004\ : InMux
    port map (
            O => \N__51334\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18205\
        );

    \I__10003\ : InMux
    port map (
            O => \N__51331\,
            I => \N__51328\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__51328\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n207\
        );

    \I__10001\ : InMux
    port map (
            O => \N__51325\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18206\
        );

    \I__10000\ : InMux
    port map (
            O => \N__51322\,
            I => \N__51319\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__51319\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n256\
        );

    \I__9998\ : InMux
    port map (
            O => \N__51316\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18207\
        );

    \I__9997\ : InMux
    port map (
            O => \N__51313\,
            I => \N__51310\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__51310\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n305\
        );

    \I__9995\ : InMux
    port map (
            O => \N__51307\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18208\
        );

    \I__9994\ : InMux
    port map (
            O => \N__51304\,
            I => \N__51301\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__51301\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n354\
        );

    \I__9992\ : InMux
    port map (
            O => \N__51298\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18209\
        );

    \I__9991\ : InMux
    port map (
            O => \N__51295\,
            I => \N__51292\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__51292\,
            I => \N__51289\
        );

    \I__9989\ : Odrv4
    port map (
            O => \N__51289\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n403\
        );

    \I__9988\ : CascadeMux
    port map (
            O => \N__51286\,
            I => \Saturate_out1_31__N_267_adj_2418_cascade_\
        );

    \I__9987\ : CascadeMux
    port map (
            O => \N__51283\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n22_adj_762_cascade_\
        );

    \I__9986\ : CascadeMux
    port map (
            O => \N__51280\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20694_cascade_\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__51277\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19729_cascade_\
        );

    \I__9984\ : InMux
    port map (
            O => \N__51274\,
            I => \N__51271\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__51271\,
            I => \N__51268\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__51268\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20676\
        );

    \I__9981\ : CascadeMux
    port map (
            O => \N__51265\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20664_cascade_\
        );

    \I__9980\ : CascadeMux
    port map (
            O => \N__51262\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20650_cascade_\
        );

    \I__9979\ : CascadeMux
    port map (
            O => \N__51259\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n58_cascade_\
        );

    \I__9978\ : CascadeMux
    port map (
            O => \N__51256\,
            I => \Saturate_out1_31__N_266_adj_2417_cascade_\
        );

    \I__9977\ : InMux
    port map (
            O => \N__51253\,
            I => \N__51250\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__51250\,
            I => \N__51247\
        );

    \I__9975\ : Odrv4
    port map (
            O => \N__51247\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20620\
        );

    \I__9974\ : InMux
    port map (
            O => \N__51244\,
            I => \N__51241\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__51241\,
            I => \N__51238\
        );

    \I__9972\ : Odrv12
    port map (
            O => \N__51238\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20608\
        );

    \I__9971\ : InMux
    port map (
            O => \N__51235\,
            I => \N__51232\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__51232\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18\
        );

    \I__9969\ : InMux
    port map (
            O => \N__51229\,
            I => \N__51226\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__51226\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n27\
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__51223\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20586_cascade_\
        );

    \I__9966\ : InMux
    port map (
            O => \N__51220\,
            I => \N__51217\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__51217\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20590\
        );

    \I__9964\ : InMux
    port map (
            O => \N__51214\,
            I => \N__51211\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__51211\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20614\
        );

    \I__9962\ : InMux
    port map (
            O => \N__51208\,
            I => \N__51205\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__51205\,
            I => \N__51201\
        );

    \I__9960\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51198\
        );

    \I__9959\ : Span4Mux_h
    port map (
            O => \N__51201\,
            I => \N__51194\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__51198\,
            I => \N__51191\
        );

    \I__9957\ : CascadeMux
    port map (
            O => \N__51197\,
            I => \N__51187\
        );

    \I__9956\ : Sp12to4
    port map (
            O => \N__51194\,
            I => \N__51182\
        );

    \I__9955\ : Span12Mux_h
    port map (
            O => \N__51191\,
            I => \N__51182\
        );

    \I__9954\ : InMux
    port map (
            O => \N__51190\,
            I => \N__51179\
        );

    \I__9953\ : InMux
    port map (
            O => \N__51187\,
            I => \N__51176\
        );

    \I__9952\ : Odrv12
    port map (
            O => \N__51182\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__51179\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__51176\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16\
        );

    \I__9949\ : CascadeMux
    port map (
            O => \N__51169\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20602_cascade_\
        );

    \I__9948\ : InMux
    port map (
            O => \N__51166\,
            I => \N__51163\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__51163\,
            I => \foc.qVoltage_7\
        );

    \I__9946\ : InMux
    port map (
            O => \N__51160\,
            I => \N__51153\
        );

    \I__9945\ : InMux
    port map (
            O => \N__51159\,
            I => \N__51153\
        );

    \I__9944\ : CascadeMux
    port map (
            O => \N__51158\,
            I => \N__51150\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__51153\,
            I => \N__51146\
        );

    \I__9942\ : InMux
    port map (
            O => \N__51150\,
            I => \N__51143\
        );

    \I__9941\ : InMux
    port map (
            O => \N__51149\,
            I => \N__51140\
        );

    \I__9940\ : Span4Mux_v
    port map (
            O => \N__51146\,
            I => \N__51132\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__51143\,
            I => \N__51132\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__51140\,
            I => \N__51132\
        );

    \I__9937\ : InMux
    port map (
            O => \N__51139\,
            I => \N__51129\
        );

    \I__9936\ : Span4Mux_v
    port map (
            O => \N__51132\,
            I => \N__51122\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__51129\,
            I => \N__51122\
        );

    \I__9934\ : InMux
    port map (
            O => \N__51128\,
            I => \N__51119\
        );

    \I__9933\ : InMux
    port map (
            O => \N__51127\,
            I => \N__51116\
        );

    \I__9932\ : Span4Mux_v
    port map (
            O => \N__51122\,
            I => \N__51113\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__51119\,
            I => \N__51108\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__51116\,
            I => \N__51108\
        );

    \I__9929\ : Span4Mux_h
    port map (
            O => \N__51113\,
            I => \N__51105\
        );

    \I__9928\ : Span4Mux_v
    port map (
            O => \N__51108\,
            I => \N__51102\
        );

    \I__9927\ : Odrv4
    port map (
            O => \N__51105\,
            I => \Error_sub_temp_31\
        );

    \I__9926\ : Odrv4
    port map (
            O => \N__51102\,
            I => \Error_sub_temp_31\
        );

    \I__9925\ : CascadeMux
    port map (
            O => \N__51097\,
            I => \N__51094\
        );

    \I__9924\ : InMux
    port map (
            O => \N__51094\,
            I => \N__51090\
        );

    \I__9923\ : InMux
    port map (
            O => \N__51093\,
            I => \N__51087\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__51090\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__51087\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424\
        );

    \I__9920\ : InMux
    port map (
            O => \N__51082\,
            I => \N__51079\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__51079\,
            I => \N__51075\
        );

    \I__9918\ : InMux
    port map (
            O => \N__51078\,
            I => \N__51072\
        );

    \I__9917\ : Span4Mux_v
    port map (
            O => \N__51075\,
            I => \N__51069\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__51072\,
            I => \N__51066\
        );

    \I__9915\ : Odrv4
    port map (
            O => \N__51069\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17\
        );

    \I__9914\ : Odrv12
    port map (
            O => \N__51066\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17\
        );

    \I__9913\ : InMux
    port map (
            O => \N__51061\,
            I => \N__51058\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__51058\,
            I => \foc.qVoltage_3\
        );

    \I__9911\ : InMux
    port map (
            O => \N__51055\,
            I => \N__51049\
        );

    \I__9910\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51049\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__51049\,
            I => \N__51046\
        );

    \I__9908\ : Span4Mux_h
    port map (
            O => \N__51046\,
            I => \N__51043\
        );

    \I__9907\ : Span4Mux_v
    port map (
            O => \N__51043\,
            I => \N__51038\
        );

    \I__9906\ : InMux
    port map (
            O => \N__51042\,
            I => \N__51035\
        );

    \I__9905\ : InMux
    port map (
            O => \N__51041\,
            I => \N__51032\
        );

    \I__9904\ : Odrv4
    port map (
            O => \N__51038\,
            I => \foc.preSatVoltage_13\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__51035\,
            I => \foc.preSatVoltage_13\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__51032\,
            I => \foc.preSatVoltage_13\
        );

    \I__9901\ : CascadeMux
    port map (
            O => \N__51025\,
            I => \foc.qVoltage_4_cascade_\
        );

    \I__9900\ : InMux
    port map (
            O => \N__51022\,
            I => \N__51018\
        );

    \I__9899\ : InMux
    port map (
            O => \N__51021\,
            I => \N__51015\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__51018\,
            I => \N__51010\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__51015\,
            I => \N__51010\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__51010\,
            I => \N__51005\
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__51009\,
            I => \N__51002\
        );

    \I__9894\ : CascadeMux
    port map (
            O => \N__51008\,
            I => \N__50999\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__51005\,
            I => \N__50996\
        );

    \I__9892\ : InMux
    port map (
            O => \N__51002\,
            I => \N__50993\
        );

    \I__9891\ : InMux
    port map (
            O => \N__50999\,
            I => \N__50990\
        );

    \I__9890\ : Odrv4
    port map (
            O => \N__50996\,
            I => \foc.preSatVoltage_12\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__50993\,
            I => \foc.preSatVoltage_12\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__50990\,
            I => \foc.preSatVoltage_12\
        );

    \I__9887\ : InMux
    port map (
            O => \N__50983\,
            I => \N__50980\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__50980\,
            I => \N__50977\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__50977\,
            I => \N__50972\
        );

    \I__9884\ : InMux
    port map (
            O => \N__50976\,
            I => \N__50967\
        );

    \I__9883\ : InMux
    port map (
            O => \N__50975\,
            I => \N__50967\
        );

    \I__9882\ : Sp12to4
    port map (
            O => \N__50972\,
            I => \N__50962\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__50967\,
            I => \N__50962\
        );

    \I__9880\ : Odrv12
    port map (
            O => \N__50962\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_26\
        );

    \I__9879\ : CascadeMux
    port map (
            O => \N__50959\,
            I => \N__50956\
        );

    \I__9878\ : InMux
    port map (
            O => \N__50956\,
            I => \N__50953\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__50953\,
            I => \N__50950\
        );

    \I__9876\ : Span4Mux_h
    port map (
            O => \N__50950\,
            I => \N__50945\
        );

    \I__9875\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50940\
        );

    \I__9874\ : InMux
    port map (
            O => \N__50948\,
            I => \N__50940\
        );

    \I__9873\ : Sp12to4
    port map (
            O => \N__50945\,
            I => \N__50935\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__50940\,
            I => \N__50935\
        );

    \I__9871\ : Odrv12
    port map (
            O => \N__50935\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_28\
        );

    \I__9870\ : InMux
    port map (
            O => \N__50932\,
            I => \N__50926\
        );

    \I__9869\ : InMux
    port map (
            O => \N__50931\,
            I => \N__50926\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__50926\,
            I => \N__50923\
        );

    \I__9867\ : Span4Mux_h
    port map (
            O => \N__50923\,
            I => \N__50919\
        );

    \I__9866\ : InMux
    port map (
            O => \N__50922\,
            I => \N__50916\
        );

    \I__9865\ : Span4Mux_v
    port map (
            O => \N__50919\,
            I => \N__50912\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__50916\,
            I => \N__50909\
        );

    \I__9863\ : InMux
    port map (
            O => \N__50915\,
            I => \N__50906\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__50912\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17\
        );

    \I__9861\ : Odrv4
    port map (
            O => \N__50909\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__50906\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17\
        );

    \I__9859\ : CascadeMux
    port map (
            O => \N__50899\,
            I => \foc.qVoltage_8_cascade_\
        );

    \I__9858\ : InMux
    port map (
            O => \N__50896\,
            I => \N__50893\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__50893\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n8265\
        );

    \I__9856\ : InMux
    port map (
            O => \N__50890\,
            I => \N__50887\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__50887\,
            I => \N__50884\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__50884\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19884\
        );

    \I__9853\ : InMux
    port map (
            O => \N__50881\,
            I => \N__50878\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__50878\,
            I => \N__50874\
        );

    \I__9851\ : CascadeMux
    port map (
            O => \N__50877\,
            I => \N__50870\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__50874\,
            I => \N__50867\
        );

    \I__9849\ : InMux
    port map (
            O => \N__50873\,
            I => \N__50862\
        );

    \I__9848\ : InMux
    port map (
            O => \N__50870\,
            I => \N__50862\
        );

    \I__9847\ : Span4Mux_v
    port map (
            O => \N__50867\,
            I => \N__50859\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__50862\,
            I => \N__50856\
        );

    \I__9845\ : Odrv4
    port map (
            O => \N__50859\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27\
        );

    \I__9844\ : Odrv12
    port map (
            O => \N__50856\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27\
        );

    \I__9843\ : CascadeMux
    port map (
            O => \N__50851\,
            I => \N__50848\
        );

    \I__9842\ : InMux
    port map (
            O => \N__50848\,
            I => \N__50845\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__50845\,
            I => \N__50842\
        );

    \I__9840\ : Span4Mux_v
    port map (
            O => \N__50842\,
            I => \N__50839\
        );

    \I__9839\ : Span4Mux_v
    port map (
            O => \N__50839\,
            I => \N__50836\
        );

    \I__9838\ : Span4Mux_v
    port map (
            O => \N__50836\,
            I => \N__50833\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__50833\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_CO\
        );

    \I__9836\ : InMux
    port map (
            O => \N__50830\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17516\
        );

    \I__9835\ : InMux
    port map (
            O => \N__50827\,
            I => \N__50824\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__50824\,
            I => \N__50821\
        );

    \I__9833\ : Span4Mux_v
    port map (
            O => \N__50821\,
            I => \N__50818\
        );

    \I__9832\ : Span4Mux_v
    port map (
            O => \N__50818\,
            I => \N__50815\
        );

    \I__9831\ : Odrv4
    port map (
            O => \N__50815\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n786_adj_348\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__50812\,
            I => \N__50809\
        );

    \I__9829\ : InMux
    port map (
            O => \N__50809\,
            I => \N__50806\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__50806\,
            I => \N__50803\
        );

    \I__9827\ : Span12Mux_h
    port map (
            O => \N__50803\,
            I => \N__50800\
        );

    \I__9826\ : Odrv12
    port map (
            O => \N__50800\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_CO\
        );

    \I__9825\ : InMux
    port map (
            O => \N__50797\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17517\
        );

    \I__9824\ : InMux
    port map (
            O => \N__50794\,
            I => \N__50791\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__50791\,
            I => \N__50788\
        );

    \I__9822\ : Span4Mux_v
    port map (
            O => \N__50788\,
            I => \N__50785\
        );

    \I__9821\ : Odrv4
    port map (
            O => \N__50785\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n790\
        );

    \I__9820\ : CascadeMux
    port map (
            O => \N__50782\,
            I => \N__50779\
        );

    \I__9819\ : InMux
    port map (
            O => \N__50779\,
            I => \N__50776\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__50776\,
            I => \N__50773\
        );

    \I__9817\ : Span4Mux_v
    port map (
            O => \N__50773\,
            I => \N__50770\
        );

    \I__9816\ : Span4Mux_v
    port map (
            O => \N__50770\,
            I => \N__50767\
        );

    \I__9815\ : Odrv4
    port map (
            O => \N__50767\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_CO\
        );

    \I__9814\ : InMux
    port map (
            O => \N__50764\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17518\
        );

    \I__9813\ : InMux
    port map (
            O => \N__50761\,
            I => \N__50758\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__50758\,
            I => \N__50755\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__50755\,
            I => n794_adj_2420
        );

    \I__9810\ : CascadeMux
    port map (
            O => \N__50752\,
            I => \N__50749\
        );

    \I__9809\ : InMux
    port map (
            O => \N__50749\,
            I => \N__50746\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__50746\,
            I => \N__50743\
        );

    \I__9807\ : Span4Mux_v
    port map (
            O => \N__50743\,
            I => \N__50740\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__50740\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n791\
        );

    \I__9805\ : InMux
    port map (
            O => \N__50737\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17519\
        );

    \I__9804\ : InMux
    port map (
            O => \N__50734\,
            I => \N__50731\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__50731\,
            I => \N__50727\
        );

    \I__9802\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50724\
        );

    \I__9801\ : Span4Mux_v
    port map (
            O => \N__50727\,
            I => \N__50719\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__50724\,
            I => \N__50719\
        );

    \I__9799\ : Odrv4
    port map (
            O => \N__50719\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n796\
        );

    \I__9798\ : InMux
    port map (
            O => \N__50716\,
            I => \bfn_20_16_0_\
        );

    \I__9797\ : CascadeMux
    port map (
            O => \N__50713\,
            I => \N__50709\
        );

    \I__9796\ : InMux
    port map (
            O => \N__50712\,
            I => \N__50703\
        );

    \I__9795\ : InMux
    port map (
            O => \N__50709\,
            I => \N__50703\
        );

    \I__9794\ : CascadeMux
    port map (
            O => \N__50708\,
            I => \N__50700\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__50703\,
            I => \N__50697\
        );

    \I__9792\ : InMux
    port map (
            O => \N__50700\,
            I => \N__50694\
        );

    \I__9791\ : Span4Mux_h
    port map (
            O => \N__50697\,
            I => \N__50690\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__50694\,
            I => \N__50687\
        );

    \I__9789\ : InMux
    port map (
            O => \N__50693\,
            I => \N__50684\
        );

    \I__9788\ : Span4Mux_v
    port map (
            O => \N__50690\,
            I => \N__50681\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__50687\,
            I => \N__50676\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__50684\,
            I => \N__50676\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__50681\,
            I => \foc.preSatVoltage_19\
        );

    \I__9784\ : Odrv4
    port map (
            O => \N__50676\,
            I => \foc.preSatVoltage_19\
        );

    \I__9783\ : InMux
    port map (
            O => \N__50671\,
            I => \N__50668\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__50668\,
            I => \foc.qVoltage_10\
        );

    \I__9781\ : InMux
    port map (
            O => \N__50665\,
            I => \N__50659\
        );

    \I__9780\ : InMux
    port map (
            O => \N__50664\,
            I => \N__50659\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__50659\,
            I => \N__50656\
        );

    \I__9778\ : Span4Mux_v
    port map (
            O => \N__50656\,
            I => \N__50651\
        );

    \I__9777\ : CascadeMux
    port map (
            O => \N__50655\,
            I => \N__50648\
        );

    \I__9776\ : CascadeMux
    port map (
            O => \N__50654\,
            I => \N__50645\
        );

    \I__9775\ : Sp12to4
    port map (
            O => \N__50651\,
            I => \N__50642\
        );

    \I__9774\ : InMux
    port map (
            O => \N__50648\,
            I => \N__50639\
        );

    \I__9773\ : InMux
    port map (
            O => \N__50645\,
            I => \N__50636\
        );

    \I__9772\ : Span12Mux_h
    port map (
            O => \N__50642\,
            I => \N__50629\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__50639\,
            I => \N__50629\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__50636\,
            I => \N__50629\
        );

    \I__9769\ : Odrv12
    port map (
            O => \N__50629\,
            I => \foc.preSatVoltage_22\
        );

    \I__9768\ : InMux
    port map (
            O => \N__50626\,
            I => \N__50623\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__50623\,
            I => \foc.qVoltage_13\
        );

    \I__9766\ : InMux
    port map (
            O => \N__50620\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17508\
        );

    \I__9765\ : InMux
    port map (
            O => \N__50617\,
            I => \N__50614\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__50614\,
            I => \N__50611\
        );

    \I__9763\ : Odrv12
    port map (
            O => \N__50611\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n754_adj_405\
        );

    \I__9762\ : InMux
    port map (
            O => \N__50608\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17509\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__50605\,
            I => \N__50602\
        );

    \I__9760\ : InMux
    port map (
            O => \N__50602\,
            I => \N__50599\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__50599\,
            I => \N__50596\
        );

    \I__9758\ : Odrv12
    port map (
            O => \N__50596\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_CO\
        );

    \I__9757\ : InMux
    port map (
            O => \N__50593\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17510\
        );

    \I__9756\ : InMux
    port map (
            O => \N__50590\,
            I => \N__50587\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__50587\,
            I => \N__50584\
        );

    \I__9754\ : Odrv12
    port map (
            O => \N__50584\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n762_adj_402\
        );

    \I__9753\ : InMux
    port map (
            O => \N__50581\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17511\
        );

    \I__9752\ : InMux
    port map (
            O => \N__50578\,
            I => \N__50575\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__50575\,
            I => \N__50572\
        );

    \I__9750\ : Span4Mux_v
    port map (
            O => \N__50572\,
            I => \N__50569\
        );

    \I__9749\ : Odrv4
    port map (
            O => \N__50569\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n766_adj_385\
        );

    \I__9748\ : CascadeMux
    port map (
            O => \N__50566\,
            I => \N__50563\
        );

    \I__9747\ : InMux
    port map (
            O => \N__50563\,
            I => \N__50560\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__50560\,
            I => \N__50557\
        );

    \I__9745\ : Odrv12
    port map (
            O => \N__50557\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_CO\
        );

    \I__9744\ : InMux
    port map (
            O => \N__50554\,
            I => \bfn_20_15_0_\
        );

    \I__9743\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50548\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__50548\,
            I => \N__50545\
        );

    \I__9741\ : Span4Mux_v
    port map (
            O => \N__50545\,
            I => \N__50542\
        );

    \I__9740\ : Span4Mux_v
    port map (
            O => \N__50542\,
            I => \N__50539\
        );

    \I__9739\ : Odrv4
    port map (
            O => \N__50539\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n770_adj_381\
        );

    \I__9738\ : CascadeMux
    port map (
            O => \N__50536\,
            I => \N__50533\
        );

    \I__9737\ : InMux
    port map (
            O => \N__50533\,
            I => \N__50530\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__50530\,
            I => \N__50527\
        );

    \I__9735\ : Span12Mux_v
    port map (
            O => \N__50527\,
            I => \N__50524\
        );

    \I__9734\ : Odrv12
    port map (
            O => \N__50524\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_CO\
        );

    \I__9733\ : InMux
    port map (
            O => \N__50521\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17513\
        );

    \I__9732\ : InMux
    port map (
            O => \N__50518\,
            I => \N__50515\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__50515\,
            I => \N__50512\
        );

    \I__9730\ : Span12Mux_v
    port map (
            O => \N__50512\,
            I => \N__50509\
        );

    \I__9729\ : Odrv12
    port map (
            O => \N__50509\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n774_adj_374\
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__50506\,
            I => \N__50503\
        );

    \I__9727\ : InMux
    port map (
            O => \N__50503\,
            I => \N__50500\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__50500\,
            I => \N__50497\
        );

    \I__9725\ : Span12Mux_v
    port map (
            O => \N__50497\,
            I => \N__50494\
        );

    \I__9724\ : Odrv12
    port map (
            O => \N__50494\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_CO\
        );

    \I__9723\ : InMux
    port map (
            O => \N__50491\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17514\
        );

    \I__9722\ : InMux
    port map (
            O => \N__50488\,
            I => \N__50485\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__50485\,
            I => \N__50482\
        );

    \I__9720\ : Span4Mux_h
    port map (
            O => \N__50482\,
            I => \N__50479\
        );

    \I__9719\ : Span4Mux_v
    port map (
            O => \N__50479\,
            I => \N__50476\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__50476\,
            I => \N__50473\
        );

    \I__9717\ : Odrv4
    port map (
            O => \N__50473\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n778_adj_356\
        );

    \I__9716\ : CascadeMux
    port map (
            O => \N__50470\,
            I => \N__50467\
        );

    \I__9715\ : InMux
    port map (
            O => \N__50467\,
            I => \N__50464\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__50464\,
            I => \N__50461\
        );

    \I__9713\ : Span12Mux_v
    port map (
            O => \N__50461\,
            I => \N__50458\
        );

    \I__9712\ : Odrv12
    port map (
            O => \N__50458\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_CO\
        );

    \I__9711\ : InMux
    port map (
            O => \N__50455\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17515\
        );

    \I__9710\ : InMux
    port map (
            O => \N__50452\,
            I => \N__50449\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__50449\,
            I => \N__50446\
        );

    \I__9708\ : Span4Mux_v
    port map (
            O => \N__50446\,
            I => \N__50443\
        );

    \I__9707\ : Span4Mux_v
    port map (
            O => \N__50443\,
            I => \N__50440\
        );

    \I__9706\ : Span4Mux_v
    port map (
            O => \N__50440\,
            I => \N__50437\
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__50437\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n782_adj_351\
        );

    \I__9704\ : CascadeMux
    port map (
            O => \N__50434\,
            I => \N__50431\
        );

    \I__9703\ : InMux
    port map (
            O => \N__50431\,
            I => \N__50428\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__50428\,
            I => \N__50425\
        );

    \I__9701\ : Sp12to4
    port map (
            O => \N__50425\,
            I => \N__50422\
        );

    \I__9700\ : Span12Mux_s11_v
    port map (
            O => \N__50422\,
            I => \N__50419\
        );

    \I__9699\ : Odrv12
    port map (
            O => \N__50419\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n721\
        );

    \I__9698\ : InMux
    port map (
            O => \N__50416\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17909\
        );

    \I__9697\ : CascadeMux
    port map (
            O => \N__50413\,
            I => \N__50410\
        );

    \I__9696\ : InMux
    port map (
            O => \N__50410\,
            I => \N__50407\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__50407\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n724\
        );

    \I__9694\ : InMux
    port map (
            O => \N__50404\,
            I => \N__50401\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__50401\,
            I => \N__50398\
        );

    \I__9692\ : Span4Mux_v
    port map (
            O => \N__50398\,
            I => \N__50395\
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__50395\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n782\
        );

    \I__9690\ : InMux
    port map (
            O => \N__50392\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17910\
        );

    \I__9689\ : InMux
    port map (
            O => \N__50389\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n783\
        );

    \I__9688\ : CascadeMux
    port map (
            O => \N__50386\,
            I => \N__50383\
        );

    \I__9687\ : InMux
    port map (
            O => \N__50383\,
            I => \N__50380\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__50380\,
            I => \N__50377\
        );

    \I__9685\ : Span4Mux_v
    port map (
            O => \N__50377\,
            I => \N__50374\
        );

    \I__9684\ : Odrv4
    port map (
            O => \N__50374\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_CO\
        );

    \I__9683\ : InMux
    port map (
            O => \N__50371\,
            I => \N__50368\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__50368\,
            I => \N__50365\
        );

    \I__9681\ : Span4Mux_v
    port map (
            O => \N__50365\,
            I => \N__50359\
        );

    \I__9680\ : InMux
    port map (
            O => \N__50364\,
            I => \N__50354\
        );

    \I__9679\ : InMux
    port map (
            O => \N__50363\,
            I => \N__50354\
        );

    \I__9678\ : InMux
    port map (
            O => \N__50362\,
            I => \N__50351\
        );

    \I__9677\ : Span4Mux_h
    port map (
            O => \N__50359\,
            I => \N__50344\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__50354\,
            I => \N__50344\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__50351\,
            I => \N__50344\
        );

    \I__9674\ : Span4Mux_v
    port map (
            O => \N__50344\,
            I => \N__50339\
        );

    \I__9673\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50336\
        );

    \I__9672\ : InMux
    port map (
            O => \N__50342\,
            I => \N__50333\
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__50339\,
            I => \Error_sub_temp_30\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__50336\,
            I => \Error_sub_temp_30\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__50333\,
            I => \Error_sub_temp_30\
        );

    \I__9668\ : InMux
    port map (
            O => \N__50326\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17505\
        );

    \I__9667\ : InMux
    port map (
            O => \N__50323\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17506\
        );

    \I__9666\ : InMux
    port map (
            O => \N__50320\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17507\
        );

    \I__9665\ : InMux
    port map (
            O => \N__50317\,
            I => \N__50314\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__50314\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n332_adj_513\
        );

    \I__9663\ : InMux
    port map (
            O => \N__50311\,
            I => \N__50308\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__50308\,
            I => \N__50305\
        );

    \I__9661\ : Span4Mux_v
    port map (
            O => \N__50305\,
            I => \N__50302\
        );

    \I__9660\ : Odrv4
    port map (
            O => \N__50302\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n378_adj_436\
        );

    \I__9659\ : InMux
    port map (
            O => \N__50299\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17902\
        );

    \I__9658\ : InMux
    port map (
            O => \N__50296\,
            I => \N__50293\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__50293\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n381\
        );

    \I__9656\ : InMux
    port map (
            O => \N__50290\,
            I => \N__50287\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__50287\,
            I => \N__50284\
        );

    \I__9654\ : Odrv4
    port map (
            O => \N__50284\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n427_adj_432\
        );

    \I__9653\ : InMux
    port map (
            O => \N__50281\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17903\
        );

    \I__9652\ : InMux
    port map (
            O => \N__50278\,
            I => \N__50275\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__50275\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n430\
        );

    \I__9650\ : InMux
    port map (
            O => \N__50272\,
            I => \N__50269\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__50269\,
            I => \N__50266\
        );

    \I__9648\ : Span4Mux_v
    port map (
            O => \N__50266\,
            I => \N__50263\
        );

    \I__9647\ : Odrv4
    port map (
            O => \N__50263\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n476\
        );

    \I__9646\ : InMux
    port map (
            O => \N__50260\,
            I => \bfn_20_12_0_\
        );

    \I__9645\ : InMux
    port map (
            O => \N__50257\,
            I => \N__50254\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__50254\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n479\
        );

    \I__9643\ : InMux
    port map (
            O => \N__50251\,
            I => \N__50248\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__50248\,
            I => \N__50245\
        );

    \I__9641\ : Span4Mux_v
    port map (
            O => \N__50245\,
            I => \N__50242\
        );

    \I__9640\ : Odrv4
    port map (
            O => \N__50242\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n525\
        );

    \I__9639\ : InMux
    port map (
            O => \N__50239\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17905\
        );

    \I__9638\ : InMux
    port map (
            O => \N__50236\,
            I => \N__50233\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__50233\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n528\
        );

    \I__9636\ : InMux
    port map (
            O => \N__50230\,
            I => \N__50227\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__50227\,
            I => \N__50224\
        );

    \I__9634\ : Span4Mux_h
    port map (
            O => \N__50224\,
            I => \N__50221\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__50221\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n574\
        );

    \I__9632\ : InMux
    port map (
            O => \N__50218\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17906\
        );

    \I__9631\ : InMux
    port map (
            O => \N__50215\,
            I => \N__50212\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__50212\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n577\
        );

    \I__9629\ : InMux
    port map (
            O => \N__50209\,
            I => \N__50206\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__50206\,
            I => \N__50203\
        );

    \I__9627\ : Span4Mux_v
    port map (
            O => \N__50203\,
            I => \N__50200\
        );

    \I__9626\ : Odrv4
    port map (
            O => \N__50200\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n623\
        );

    \I__9625\ : InMux
    port map (
            O => \N__50197\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17907\
        );

    \I__9624\ : InMux
    port map (
            O => \N__50194\,
            I => \N__50191\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__50191\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n626\
        );

    \I__9622\ : CascadeMux
    port map (
            O => \N__50188\,
            I => \N__50185\
        );

    \I__9621\ : InMux
    port map (
            O => \N__50185\,
            I => \N__50182\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__50182\,
            I => \N__50179\
        );

    \I__9619\ : Span4Mux_h
    port map (
            O => \N__50179\,
            I => \N__50176\
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__50176\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n672\
        );

    \I__9617\ : InMux
    port map (
            O => \N__50173\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17908\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__50170\,
            I => \N__50167\
        );

    \I__9615\ : InMux
    port map (
            O => \N__50167\,
            I => \N__50164\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__50164\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n675\
        );

    \I__9613\ : InMux
    port map (
            O => \N__50161\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17593\
        );

    \I__9612\ : InMux
    port map (
            O => \N__50158\,
            I => \N__50155\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__50155\,
            I => \N__50151\
        );

    \I__9610\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50148\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__50151\,
            I => \N__50143\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__50148\,
            I => \N__50143\
        );

    \I__9607\ : Span4Mux_h
    port map (
            O => \N__50143\,
            I => \N__50140\
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__50140\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n753\
        );

    \I__9605\ : InMux
    port map (
            O => \N__50137\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17594\
        );

    \I__9604\ : InMux
    port map (
            O => \N__50134\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404\
        );

    \I__9603\ : InMux
    port map (
            O => \N__50131\,
            I => \N__50128\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__50128\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n87\
        );

    \I__9601\ : InMux
    port map (
            O => \N__50125\,
            I => \N__50122\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__50122\,
            I => \N__50119\
        );

    \I__9599\ : Span4Mux_v
    port map (
            O => \N__50119\,
            I => \N__50116\
        );

    \I__9598\ : Odrv4
    port map (
            O => \N__50116\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n133_adj_388\
        );

    \I__9597\ : InMux
    port map (
            O => \N__50113\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17897\
        );

    \I__9596\ : InMux
    port map (
            O => \N__50110\,
            I => \N__50107\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__50107\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n136\
        );

    \I__9594\ : InMux
    port map (
            O => \N__50104\,
            I => \N__50101\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__50101\,
            I => \N__50098\
        );

    \I__9592\ : Span4Mux_h
    port map (
            O => \N__50098\,
            I => \N__50095\
        );

    \I__9591\ : Odrv4
    port map (
            O => \N__50095\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n182_adj_451\
        );

    \I__9590\ : InMux
    port map (
            O => \N__50092\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17898\
        );

    \I__9589\ : InMux
    port map (
            O => \N__50089\,
            I => \N__50086\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__50086\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n185\
        );

    \I__9587\ : InMux
    port map (
            O => \N__50083\,
            I => \N__50080\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__50080\,
            I => \N__50077\
        );

    \I__9585\ : Span12Mux_h
    port map (
            O => \N__50077\,
            I => \N__50074\
        );

    \I__9584\ : Odrv12
    port map (
            O => \N__50074\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n231_adj_387\
        );

    \I__9583\ : InMux
    port map (
            O => \N__50071\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17899\
        );

    \I__9582\ : InMux
    port map (
            O => \N__50068\,
            I => \N__50065\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__50065\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n234\
        );

    \I__9580\ : InMux
    port map (
            O => \N__50062\,
            I => \N__50059\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__50059\,
            I => \N__50056\
        );

    \I__9578\ : Span4Mux_h
    port map (
            O => \N__50056\,
            I => \N__50053\
        );

    \I__9577\ : Odrv4
    port map (
            O => \N__50053\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n280_adj_379\
        );

    \I__9576\ : InMux
    port map (
            O => \N__50050\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17900\
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__50047\,
            I => \N__50044\
        );

    \I__9574\ : InMux
    port map (
            O => \N__50044\,
            I => \N__50041\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__50041\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n283_adj_514\
        );

    \I__9572\ : InMux
    port map (
            O => \N__50038\,
            I => \N__50035\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__50035\,
            I => \N__50032\
        );

    \I__9570\ : Span4Mux_h
    port map (
            O => \N__50032\,
            I => \N__50029\
        );

    \I__9569\ : Odrv4
    port map (
            O => \N__50029\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n329_adj_439\
        );

    \I__9568\ : InMux
    port map (
            O => \N__50026\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17901\
        );

    \I__9567\ : InMux
    port map (
            O => \N__50023\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17584\
        );

    \I__9566\ : InMux
    port map (
            O => \N__50020\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17585\
        );

    \I__9565\ : InMux
    port map (
            O => \N__50017\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17586\
        );

    \I__9564\ : InMux
    port map (
            O => \N__50014\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17587\
        );

    \I__9563\ : InMux
    port map (
            O => \N__50011\,
            I => \bfn_20_10_0_\
        );

    \I__9562\ : InMux
    port map (
            O => \N__50008\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17589\
        );

    \I__9561\ : InMux
    port map (
            O => \N__50005\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17590\
        );

    \I__9560\ : InMux
    port map (
            O => \N__50002\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17591\
        );

    \I__9559\ : InMux
    port map (
            O => \N__49999\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17592\
        );

    \I__9558\ : InMux
    port map (
            O => \N__49996\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17621\
        );

    \I__9557\ : InMux
    port map (
            O => \N__49993\,
            I => \N__49990\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__49990\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n611\
        );

    \I__9555\ : InMux
    port map (
            O => \N__49987\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17622\
        );

    \I__9554\ : CascadeMux
    port map (
            O => \N__49984\,
            I => \N__49981\
        );

    \I__9553\ : InMux
    port map (
            O => \N__49981\,
            I => \N__49978\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__49978\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n660\
        );

    \I__9551\ : InMux
    port map (
            O => \N__49975\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17623\
        );

    \I__9550\ : InMux
    port map (
            O => \N__49972\,
            I => \N__49969\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__49969\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n709_adj_512\
        );

    \I__9548\ : CascadeMux
    port map (
            O => \N__49966\,
            I => \N__49963\
        );

    \I__9547\ : InMux
    port map (
            O => \N__49963\,
            I => \N__49960\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__49960\,
            I => \N__49957\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__49957\,
            I => \N__49953\
        );

    \I__9544\ : InMux
    port map (
            O => \N__49956\,
            I => \N__49950\
        );

    \I__9543\ : Odrv4
    port map (
            O => \N__49953\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n761\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__49950\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n761\
        );

    \I__9541\ : InMux
    port map (
            O => \N__49945\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17624\
        );

    \I__9540\ : InMux
    port map (
            O => \N__49942\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386\
        );

    \I__9539\ : InMux
    port map (
            O => \N__49939\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17581\
        );

    \I__9538\ : InMux
    port map (
            O => \N__49936\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17582\
        );

    \I__9537\ : InMux
    port map (
            O => \N__49933\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17583\
        );

    \I__9536\ : InMux
    port map (
            O => \N__49930\,
            I => \N__49927\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__49927\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n170_adj_490\
        );

    \I__9534\ : InMux
    port map (
            O => \N__49924\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17613\
        );

    \I__9533\ : InMux
    port map (
            O => \N__49921\,
            I => \N__49918\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__49918\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n219_adj_472\
        );

    \I__9531\ : InMux
    port map (
            O => \N__49915\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17614\
        );

    \I__9530\ : InMux
    port map (
            O => \N__49912\,
            I => \N__49909\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__49909\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n268\
        );

    \I__9528\ : InMux
    port map (
            O => \N__49906\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17615\
        );

    \I__9527\ : InMux
    port map (
            O => \N__49903\,
            I => \N__49900\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__49900\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n317\
        );

    \I__9525\ : InMux
    port map (
            O => \N__49897\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17616\
        );

    \I__9524\ : InMux
    port map (
            O => \N__49894\,
            I => \N__49891\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__49891\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n366\
        );

    \I__9522\ : InMux
    port map (
            O => \N__49888\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17617\
        );

    \I__9521\ : InMux
    port map (
            O => \N__49885\,
            I => \N__49882\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__49882\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n415_adj_449\
        );

    \I__9519\ : InMux
    port map (
            O => \N__49879\,
            I => \bfn_20_8_0_\
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__49876\,
            I => \N__49873\
        );

    \I__9517\ : InMux
    port map (
            O => \N__49873\,
            I => \N__49870\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__49870\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n464\
        );

    \I__9515\ : InMux
    port map (
            O => \N__49867\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17619\
        );

    \I__9514\ : InMux
    port map (
            O => \N__49864\,
            I => \N__49861\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__49861\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n513\
        );

    \I__9512\ : InMux
    port map (
            O => \N__49858\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17620\
        );

    \I__9511\ : CascadeMux
    port map (
            O => \N__49855\,
            I => \N__49852\
        );

    \I__9510\ : InMux
    port map (
            O => \N__49852\,
            I => \N__49849\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__49849\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n562\
        );

    \I__9508\ : InMux
    port map (
            O => \N__49846\,
            I => \N__49843\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__49843\,
            I => \N__49840\
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__49840\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n473\
        );

    \I__9505\ : CascadeMux
    port map (
            O => \N__49837\,
            I => \N__49834\
        );

    \I__9504\ : InMux
    port map (
            O => \N__49834\,
            I => \N__49831\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__49831\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n519\
        );

    \I__9502\ : InMux
    port map (
            O => \N__49828\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18130\
        );

    \I__9501\ : InMux
    port map (
            O => \N__49825\,
            I => \N__49822\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__49822\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n568\
        );

    \I__9499\ : InMux
    port map (
            O => \N__49819\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18131\
        );

    \I__9498\ : CascadeMux
    port map (
            O => \N__49816\,
            I => \N__49811\
        );

    \I__9497\ : InMux
    port map (
            O => \N__49815\,
            I => \N__49808\
        );

    \I__9496\ : InMux
    port map (
            O => \N__49814\,
            I => \N__49803\
        );

    \I__9495\ : InMux
    port map (
            O => \N__49811\,
            I => \N__49803\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__49808\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n617\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__49803\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n617\
        );

    \I__9492\ : InMux
    port map (
            O => \N__49798\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18132\
        );

    \I__9491\ : InMux
    port map (
            O => \N__49795\,
            I => \N__49791\
        );

    \I__9490\ : InMux
    port map (
            O => \N__49794\,
            I => \N__49788\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__49791\,
            I => \N__49785\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__49788\,
            I => \N__49782\
        );

    \I__9487\ : Span4Mux_h
    port map (
            O => \N__49785\,
            I => \N__49779\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__49782\,
            I => \N__49776\
        );

    \I__9485\ : Odrv4
    port map (
            O => \N__49779\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n773\
        );

    \I__9484\ : Odrv4
    port map (
            O => \N__49776\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n773\
        );

    \I__9483\ : CascadeMux
    port map (
            O => \N__49771\,
            I => \N__49767\
        );

    \I__9482\ : CascadeMux
    port map (
            O => \N__49770\,
            I => \N__49764\
        );

    \I__9481\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49760\
        );

    \I__9480\ : InMux
    port map (
            O => \N__49764\,
            I => \N__49755\
        );

    \I__9479\ : InMux
    port map (
            O => \N__49763\,
            I => \N__49755\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__49760\,
            I => \N__49750\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__49755\,
            I => \N__49750\
        );

    \I__9476\ : Odrv4
    port map (
            O => \N__49750\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n522\
        );

    \I__9475\ : InMux
    port map (
            O => \N__49747\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18133\
        );

    \I__9474\ : InMux
    port map (
            O => \N__49744\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357\
        );

    \I__9473\ : InMux
    port map (
            O => \N__49741\,
            I => \N__49738\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__49738\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n72_adj_508\
        );

    \I__9471\ : InMux
    port map (
            O => \N__49735\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17611\
        );

    \I__9470\ : CascadeMux
    port map (
            O => \N__49732\,
            I => \N__49729\
        );

    \I__9469\ : InMux
    port map (
            O => \N__49729\,
            I => \N__49726\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__49726\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n121_adj_504\
        );

    \I__9467\ : InMux
    port map (
            O => \N__49723\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17612\
        );

    \I__9466\ : CascadeMux
    port map (
            O => \N__49720\,
            I => \N__49717\
        );

    \I__9465\ : InMux
    port map (
            O => \N__49717\,
            I => \N__49714\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__49714\,
            I => \N__49711\
        );

    \I__9463\ : Odrv12
    port map (
            O => \N__49711\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n81\
        );

    \I__9462\ : InMux
    port map (
            O => \N__49708\,
            I => \N__49705\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__49705\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n127\
        );

    \I__9460\ : InMux
    port map (
            O => \N__49702\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18122\
        );

    \I__9459\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49696\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__49696\,
            I => \N__49693\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__49693\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n130\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__49690\,
            I => \N__49687\
        );

    \I__9455\ : InMux
    port map (
            O => \N__49687\,
            I => \N__49684\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__49684\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n176\
        );

    \I__9453\ : InMux
    port map (
            O => \N__49681\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18123\
        );

    \I__9452\ : CascadeMux
    port map (
            O => \N__49678\,
            I => \N__49675\
        );

    \I__9451\ : InMux
    port map (
            O => \N__49675\,
            I => \N__49672\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__49672\,
            I => \N__49669\
        );

    \I__9449\ : Odrv12
    port map (
            O => \N__49669\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n179\
        );

    \I__9448\ : InMux
    port map (
            O => \N__49666\,
            I => \N__49663\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__49663\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n225\
        );

    \I__9446\ : InMux
    port map (
            O => \N__49660\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18124\
        );

    \I__9445\ : InMux
    port map (
            O => \N__49657\,
            I => \N__49654\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__49654\,
            I => \N__49651\
        );

    \I__9443\ : Odrv12
    port map (
            O => \N__49651\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n228\
        );

    \I__9442\ : InMux
    port map (
            O => \N__49648\,
            I => \N__49645\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__49645\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n274\
        );

    \I__9440\ : InMux
    port map (
            O => \N__49642\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18125\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__49639\,
            I => \N__49636\
        );

    \I__9438\ : InMux
    port map (
            O => \N__49636\,
            I => \N__49633\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__49633\,
            I => \N__49630\
        );

    \I__9436\ : Odrv4
    port map (
            O => \N__49630\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n277\
        );

    \I__9435\ : InMux
    port map (
            O => \N__49627\,
            I => \N__49624\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__49624\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n323\
        );

    \I__9433\ : InMux
    port map (
            O => \N__49621\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18126\
        );

    \I__9432\ : CascadeMux
    port map (
            O => \N__49618\,
            I => \N__49615\
        );

    \I__9431\ : InMux
    port map (
            O => \N__49615\,
            I => \N__49612\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__49612\,
            I => \N__49609\
        );

    \I__9429\ : Odrv12
    port map (
            O => \N__49609\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n326\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__49606\,
            I => \N__49603\
        );

    \I__9427\ : InMux
    port map (
            O => \N__49603\,
            I => \N__49600\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__49600\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n372\
        );

    \I__9425\ : InMux
    port map (
            O => \N__49597\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18127\
        );

    \I__9424\ : InMux
    port map (
            O => \N__49594\,
            I => \N__49591\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__49591\,
            I => \N__49588\
        );

    \I__9422\ : Odrv12
    port map (
            O => \N__49588\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n375\
        );

    \I__9421\ : CascadeMux
    port map (
            O => \N__49585\,
            I => \N__49582\
        );

    \I__9420\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49579\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__49579\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n421\
        );

    \I__9418\ : InMux
    port map (
            O => \N__49576\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18128\
        );

    \I__9417\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49570\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__49570\,
            I => \N__49567\
        );

    \I__9415\ : Span4Mux_h
    port map (
            O => \N__49567\,
            I => \N__49564\
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__49564\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n424\
        );

    \I__9413\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49558\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__49558\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n470\
        );

    \I__9411\ : InMux
    port map (
            O => \N__49555\,
            I => \bfn_20_6_0_\
        );

    \I__9410\ : InMux
    port map (
            O => \N__49552\,
            I => \bfn_19_29_0_\
        );

    \I__9409\ : InMux
    port map (
            O => \N__49549\,
            I => \N__49546\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__49546\,
            I => \N__49543\
        );

    \I__9407\ : Odrv4
    port map (
            O => \N__49543\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n479\
        );

    \I__9406\ : InMux
    port map (
            O => \N__49540\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18332\
        );

    \I__9405\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49534\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__49534\,
            I => \N__49531\
        );

    \I__9403\ : Odrv4
    port map (
            O => \N__49531\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n528\
        );

    \I__9402\ : InMux
    port map (
            O => \N__49528\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18333\
        );

    \I__9401\ : InMux
    port map (
            O => \N__49525\,
            I => \N__49522\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__49522\,
            I => \N__49519\
        );

    \I__9399\ : Odrv12
    port map (
            O => \N__49519\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n577\
        );

    \I__9398\ : InMux
    port map (
            O => \N__49516\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18334\
        );

    \I__9397\ : InMux
    port map (
            O => \N__49513\,
            I => \N__49510\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__49510\,
            I => \N__49507\
        );

    \I__9395\ : Odrv12
    port map (
            O => \N__49507\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n626\
        );

    \I__9394\ : InMux
    port map (
            O => \N__49504\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18335\
        );

    \I__9393\ : CascadeMux
    port map (
            O => \N__49501\,
            I => \N__49498\
        );

    \I__9392\ : InMux
    port map (
            O => \N__49498\,
            I => \N__49495\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__49495\,
            I => \N__49492\
        );

    \I__9390\ : Span4Mux_v
    port map (
            O => \N__49492\,
            I => \N__49489\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__49489\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n675\
        );

    \I__9388\ : InMux
    port map (
            O => \N__49486\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18336\
        );

    \I__9387\ : InMux
    port map (
            O => \N__49483\,
            I => \N__49480\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__49480\,
            I => \N__49477\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__49477\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n724\
        );

    \I__9384\ : InMux
    port map (
            O => \N__49474\,
            I => \N__49471\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__49471\,
            I => \N__49468\
        );

    \I__9382\ : Span12Mux_v
    port map (
            O => \N__49468\,
            I => \N__49465\
        );

    \I__9381\ : Odrv12
    port map (
            O => \N__49465\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n782\
        );

    \I__9380\ : InMux
    port map (
            O => \N__49462\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18337\
        );

    \I__9379\ : InMux
    port map (
            O => \N__49459\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__49456\,
            I => \N__49453\
        );

    \I__9377\ : InMux
    port map (
            O => \N__49453\,
            I => \N__49450\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__49450\,
            I => \N__49447\
        );

    \I__9375\ : Span12Mux_v
    port map (
            O => \N__49447\,
            I => \N__49444\
        );

    \I__9374\ : Odrv12
    port map (
            O => \N__49444\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_CO\
        );

    \I__9373\ : CascadeMux
    port map (
            O => \N__49441\,
            I => \N__49438\
        );

    \I__9372\ : InMux
    port map (
            O => \N__49438\,
            I => \N__49435\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__49435\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n78\
        );

    \I__9370\ : CascadeMux
    port map (
            O => \N__49432\,
            I => \N__49429\
        );

    \I__9369\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49426\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__49426\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n87\
        );

    \I__9367\ : InMux
    port map (
            O => \N__49423\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18324\
        );

    \I__9366\ : InMux
    port map (
            O => \N__49420\,
            I => \N__49417\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__49417\,
            I => \N__49414\
        );

    \I__9364\ : Odrv4
    port map (
            O => \N__49414\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n136\
        );

    \I__9363\ : InMux
    port map (
            O => \N__49411\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18325\
        );

    \I__9362\ : CascadeMux
    port map (
            O => \N__49408\,
            I => \N__49405\
        );

    \I__9361\ : InMux
    port map (
            O => \N__49405\,
            I => \N__49402\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__49402\,
            I => \N__49399\
        );

    \I__9359\ : Odrv4
    port map (
            O => \N__49399\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n185\
        );

    \I__9358\ : InMux
    port map (
            O => \N__49396\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18326\
        );

    \I__9357\ : InMux
    port map (
            O => \N__49393\,
            I => \N__49390\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__49390\,
            I => \N__49387\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__49387\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n234\
        );

    \I__9354\ : InMux
    port map (
            O => \N__49384\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18327\
        );

    \I__9353\ : InMux
    port map (
            O => \N__49381\,
            I => \N__49378\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__49378\,
            I => \N__49375\
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__49375\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n283\
        );

    \I__9350\ : InMux
    port map (
            O => \N__49372\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18328\
        );

    \I__9349\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49366\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__49366\,
            I => \N__49363\
        );

    \I__9347\ : Odrv4
    port map (
            O => \N__49363\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n332\
        );

    \I__9346\ : InMux
    port map (
            O => \N__49360\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18329\
        );

    \I__9345\ : InMux
    port map (
            O => \N__49357\,
            I => \N__49354\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__49354\,
            I => \N__49351\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__49351\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n381\
        );

    \I__9342\ : InMux
    port map (
            O => \N__49348\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18330\
        );

    \I__9341\ : InMux
    port map (
            O => \N__49345\,
            I => \N__49342\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__49342\,
            I => \N__49339\
        );

    \I__9339\ : Odrv12
    port map (
            O => \N__49339\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n430\
        );

    \I__9338\ : CascadeMux
    port map (
            O => \N__49336\,
            I => \N__49333\
        );

    \I__9337\ : InMux
    port map (
            O => \N__49333\,
            I => \N__49330\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__49330\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n433\
        );

    \I__9335\ : InMux
    port map (
            O => \N__49327\,
            I => \bfn_19_27_0_\
        );

    \I__9334\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49321\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__49321\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n482\
        );

    \I__9332\ : InMux
    port map (
            O => \N__49318\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18347\
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__49315\,
            I => \N__49312\
        );

    \I__9330\ : InMux
    port map (
            O => \N__49312\,
            I => \N__49309\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__49309\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n531\
        );

    \I__9328\ : InMux
    port map (
            O => \N__49306\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18348\
        );

    \I__9327\ : InMux
    port map (
            O => \N__49303\,
            I => \N__49300\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__49300\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n580\
        );

    \I__9325\ : InMux
    port map (
            O => \N__49297\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18349\
        );

    \I__9324\ : InMux
    port map (
            O => \N__49294\,
            I => \N__49291\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__49291\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n629\
        );

    \I__9322\ : InMux
    port map (
            O => \N__49288\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18350\
        );

    \I__9321\ : InMux
    port map (
            O => \N__49285\,
            I => \N__49282\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__49282\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n678\
        );

    \I__9319\ : InMux
    port map (
            O => \N__49279\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18351\
        );

    \I__9318\ : CascadeMux
    port map (
            O => \N__49276\,
            I => \N__49273\
        );

    \I__9317\ : InMux
    port map (
            O => \N__49273\,
            I => \N__49270\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__49270\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n727\
        );

    \I__9315\ : InMux
    port map (
            O => \N__49267\,
            I => \N__49264\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__49264\,
            I => \N__49261\
        );

    \I__9313\ : Odrv12
    port map (
            O => \N__49261\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n786\
        );

    \I__9312\ : InMux
    port map (
            O => \N__49258\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18352\
        );

    \I__9311\ : InMux
    port map (
            O => \N__49255\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__49252\,
            I => \N__49249\
        );

    \I__9309\ : InMux
    port map (
            O => \N__49249\,
            I => \N__49246\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__49246\,
            I => \N__49243\
        );

    \I__9307\ : Span4Mux_v
    port map (
            O => \N__49243\,
            I => \N__49240\
        );

    \I__9306\ : Odrv4
    port map (
            O => \N__49240\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_CO\
        );

    \I__9305\ : InMux
    port map (
            O => \N__49237\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__49234\,
            I => \N__49231\
        );

    \I__9303\ : InMux
    port map (
            O => \N__49231\,
            I => \N__49228\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__49228\,
            I => \N__49225\
        );

    \I__9301\ : Odrv12
    port map (
            O => \N__49225\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_CO\
        );

    \I__9300\ : InMux
    port map (
            O => \N__49222\,
            I => \N__49219\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__49219\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n90\
        );

    \I__9298\ : InMux
    port map (
            O => \N__49216\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18339\
        );

    \I__9297\ : CascadeMux
    port map (
            O => \N__49213\,
            I => \N__49210\
        );

    \I__9296\ : InMux
    port map (
            O => \N__49210\,
            I => \N__49207\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__49207\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n139\
        );

    \I__9294\ : InMux
    port map (
            O => \N__49204\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18340\
        );

    \I__9293\ : InMux
    port map (
            O => \N__49201\,
            I => \N__49198\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__49198\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n188\
        );

    \I__9291\ : InMux
    port map (
            O => \N__49195\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18341\
        );

    \I__9290\ : InMux
    port map (
            O => \N__49192\,
            I => \N__49189\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__49189\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n237\
        );

    \I__9288\ : InMux
    port map (
            O => \N__49186\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18342\
        );

    \I__9287\ : InMux
    port map (
            O => \N__49183\,
            I => \N__49180\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__49180\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n286\
        );

    \I__9285\ : InMux
    port map (
            O => \N__49177\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18343\
        );

    \I__9284\ : InMux
    port map (
            O => \N__49174\,
            I => \N__49171\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__49171\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n335\
        );

    \I__9282\ : InMux
    port map (
            O => \N__49168\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18344\
        );

    \I__9281\ : InMux
    port map (
            O => \N__49165\,
            I => \N__49162\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__49162\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n384\
        );

    \I__9279\ : InMux
    port map (
            O => \N__49159\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18345\
        );

    \I__9278\ : InMux
    port map (
            O => \N__49156\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18194\
        );

    \I__9277\ : InMux
    port map (
            O => \N__49153\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18195\
        );

    \I__9276\ : InMux
    port map (
            O => \N__49150\,
            I => \bfn_19_25_0_\
        );

    \I__9275\ : InMux
    port map (
            O => \N__49147\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18197\
        );

    \I__9274\ : InMux
    port map (
            O => \N__49144\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18198\
        );

    \I__9273\ : InMux
    port map (
            O => \N__49141\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18199\
        );

    \I__9272\ : InMux
    port map (
            O => \N__49138\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18200\
        );

    \I__9271\ : InMux
    port map (
            O => \N__49135\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18201\
        );

    \I__9270\ : InMux
    port map (
            O => \N__49132\,
            I => \N__49129\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__49129\,
            I => \N__49126\
        );

    \I__9268\ : Odrv12
    port map (
            O => \N__49126\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n746\
        );

    \I__9267\ : InMux
    port map (
            O => \N__49123\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18202\
        );

    \I__9266\ : InMux
    port map (
            O => \N__49120\,
            I => \N__49117\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__49117\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n60\
        );

    \I__9264\ : InMux
    port map (
            O => \N__49114\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18189\
        );

    \I__9263\ : InMux
    port map (
            O => \N__49111\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18190\
        );

    \I__9262\ : InMux
    port map (
            O => \N__49108\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18191\
        );

    \I__9261\ : InMux
    port map (
            O => \N__49105\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18192\
        );

    \I__9260\ : InMux
    port map (
            O => \N__49102\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18193\
        );

    \I__9259\ : InMux
    port map (
            O => \N__49099\,
            I => \bfn_19_22_0_\
        );

    \I__9258\ : InMux
    port map (
            O => \N__49096\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18152\
        );

    \I__9257\ : InMux
    port map (
            O => \N__49093\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18153\
        );

    \I__9256\ : InMux
    port map (
            O => \N__49090\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18154\
        );

    \I__9255\ : InMux
    port map (
            O => \N__49087\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18155\
        );

    \I__9254\ : InMux
    port map (
            O => \N__49084\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18156\
        );

    \I__9253\ : InMux
    port map (
            O => \N__49081\,
            I => \N__49078\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__49078\,
            I => \N__49075\
        );

    \I__9251\ : Span4Mux_v
    port map (
            O => \N__49075\,
            I => \N__49072\
        );

    \I__9250\ : Odrv4
    port map (
            O => \N__49072\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n790\
        );

    \I__9249\ : InMux
    port map (
            O => \N__49069\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18157\
        );

    \I__9248\ : InMux
    port map (
            O => \N__49066\,
            I => \N__49063\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__49063\,
            I => \N__49060\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__49060\,
            I => \N__49057\
        );

    \I__9245\ : Span4Mux_v
    port map (
            O => \N__49057\,
            I => \N__49054\
        );

    \I__9244\ : Odrv4
    port map (
            O => \N__49054\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n794\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__49051\,
            I => \N__49048\
        );

    \I__9242\ : InMux
    port map (
            O => \N__49048\,
            I => \N__49045\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__49045\,
            I => \N__49042\
        );

    \I__9240\ : Span12Mux_h
    port map (
            O => \N__49042\,
            I => \N__49039\
        );

    \I__9239\ : Odrv12
    port map (
            O => \N__49039\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_CO\
        );

    \I__9238\ : InMux
    port map (
            O => \N__49036\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18158\
        );

    \I__9237\ : InMux
    port map (
            O => \N__49033\,
            I => \N__49030\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__49030\,
            I => \N__49027\
        );

    \I__9235\ : Span4Mux_h
    port map (
            O => \N__49027\,
            I => \N__49024\
        );

    \I__9234\ : Odrv4
    port map (
            O => \N__49024\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_CO\
        );

    \I__9233\ : CascadeMux
    port map (
            O => \N__49021\,
            I => \N__49018\
        );

    \I__9232\ : InMux
    port map (
            O => \N__49018\,
            I => \N__49015\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__49015\,
            I => \N__49012\
        );

    \I__9230\ : Span4Mux_v
    port map (
            O => \N__49012\,
            I => \N__49008\
        );

    \I__9229\ : InMux
    port map (
            O => \N__49011\,
            I => \N__49005\
        );

    \I__9228\ : Span4Mux_h
    port map (
            O => \N__49008\,
            I => \N__49002\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48999\
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__49002\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n796\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__48999\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n796\
        );

    \I__9224\ : InMux
    port map (
            O => \N__48994\,
            I => \bfn_19_23_0_\
        );

    \I__9223\ : CascadeMux
    port map (
            O => \N__48991\,
            I => \N__48988\
        );

    \I__9222\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48984\
        );

    \I__9221\ : InMux
    port map (
            O => \N__48987\,
            I => \N__48981\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__48984\,
            I => \N__48976\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__48981\,
            I => \N__48976\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__48976\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n738\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__48973\,
            I => \N__48970\
        );

    \I__9216\ : InMux
    port map (
            O => \N__48970\,
            I => \N__48962\
        );

    \I__9215\ : InMux
    port map (
            O => \N__48969\,
            I => \N__48962\
        );

    \I__9214\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48959\
        );

    \I__9213\ : InMux
    port map (
            O => \N__48967\,
            I => \N__48956\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__48962\,
            I => \N__48953\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__48959\,
            I => \N__48947\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__48956\,
            I => \N__48947\
        );

    \I__9209\ : Sp12to4
    port map (
            O => \N__48953\,
            I => \N__48944\
        );

    \I__9208\ : InMux
    port map (
            O => \N__48952\,
            I => \N__48941\
        );

    \I__9207\ : Span4Mux_v
    port map (
            O => \N__48947\,
            I => \N__48936\
        );

    \I__9206\ : Span12Mux_v
    port map (
            O => \N__48944\,
            I => \N__48931\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__48941\,
            I => \N__48931\
        );

    \I__9204\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48926\
        );

    \I__9203\ : InMux
    port map (
            O => \N__48939\,
            I => \N__48926\
        );

    \I__9202\ : Odrv4
    port map (
            O => \N__48936\,
            I => \Error_sub_temp_31_adj_2384\
        );

    \I__9201\ : Odrv12
    port map (
            O => \N__48931\,
            I => \Error_sub_temp_31_adj_2384\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__48926\,
            I => \Error_sub_temp_31_adj_2384\
        );

    \I__9199\ : InMux
    port map (
            O => \N__48919\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18144\
        );

    \I__9198\ : InMux
    port map (
            O => \N__48916\,
            I => \N__48913\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__48913\,
            I => \N__48910\
        );

    \I__9196\ : Odrv4
    port map (
            O => \N__48910\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n8356\
        );

    \I__9195\ : InMux
    port map (
            O => \N__48907\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18145\
        );

    \I__9194\ : InMux
    port map (
            O => \N__48904\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18146\
        );

    \I__9193\ : InMux
    port map (
            O => \N__48901\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18147\
        );

    \I__9192\ : InMux
    port map (
            O => \N__48898\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18148\
        );

    \I__9191\ : InMux
    port map (
            O => \N__48895\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18149\
        );

    \I__9190\ : InMux
    port map (
            O => \N__48892\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18150\
        );

    \I__9189\ : InMux
    port map (
            O => \N__48889\,
            I => \N__48886\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__48886\,
            I => \N__48883\
        );

    \I__9187\ : Span4Mux_v
    port map (
            O => \N__48883\,
            I => \N__48880\
        );

    \I__9186\ : Span4Mux_v
    port map (
            O => \N__48880\,
            I => \N__48877\
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__48877\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_CO\
        );

    \I__9184\ : InMux
    port map (
            O => \N__48874\,
            I => \bfn_19_19_0_\
        );

    \I__9183\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48868\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__48868\,
            I => \N__48864\
        );

    \I__9181\ : InMux
    port map (
            O => \N__48867\,
            I => \N__48861\
        );

    \I__9180\ : Odrv4
    port map (
            O => \N__48864\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__48861\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8\
        );

    \I__9178\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48853\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__48853\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20870\
        );

    \I__9176\ : CascadeMux
    port map (
            O => \N__48850\,
            I => \N__48847\
        );

    \I__9175\ : InMux
    port map (
            O => \N__48847\,
            I => \N__48844\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__48844\,
            I => \N__48841\
        );

    \I__9173\ : Span12Mux_h
    port map (
            O => \N__48841\,
            I => \N__48836\
        );

    \I__9172\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48833\
        );

    \I__9171\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48830\
        );

    \I__9170\ : Odrv12
    port map (
            O => \N__48836\,
            I => \foc.preSatVoltage_10\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__48833\,
            I => \foc.preSatVoltage_10\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__48830\,
            I => \foc.preSatVoltage_10\
        );

    \I__9167\ : InMux
    port map (
            O => \N__48823\,
            I => \N__48820\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__48820\,
            I => \N__48816\
        );

    \I__9165\ : InMux
    port map (
            O => \N__48819\,
            I => \N__48813\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__48816\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__48813\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9\
        );

    \I__9162\ : InMux
    port map (
            O => \N__48808\,
            I => \N__48805\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__48805\,
            I => \N__48802\
        );

    \I__9160\ : Odrv12
    port map (
            O => \N__48802\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_CO\
        );

    \I__9159\ : CascadeMux
    port map (
            O => \N__48799\,
            I => \N__48796\
        );

    \I__9158\ : InMux
    port map (
            O => \N__48796\,
            I => \N__48793\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__48793\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n766\
        );

    \I__9156\ : InMux
    port map (
            O => \N__48790\,
            I => \bfn_19_18_0_\
        );

    \I__9155\ : InMux
    port map (
            O => \N__48787\,
            I => \N__48784\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__48784\,
            I => \N__48781\
        );

    \I__9153\ : Odrv4
    port map (
            O => \N__48781\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n770\
        );

    \I__9152\ : CascadeMux
    port map (
            O => \N__48778\,
            I => \N__48775\
        );

    \I__9151\ : InMux
    port map (
            O => \N__48775\,
            I => \N__48772\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__48772\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_CO\
        );

    \I__9149\ : InMux
    port map (
            O => \N__48769\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17719\
        );

    \I__9148\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48763\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__48763\,
            I => \N__48760\
        );

    \I__9146\ : Span4Mux_v
    port map (
            O => \N__48760\,
            I => \N__48757\
        );

    \I__9145\ : Odrv4
    port map (
            O => \N__48757\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n774\
        );

    \I__9144\ : CascadeMux
    port map (
            O => \N__48754\,
            I => \N__48751\
        );

    \I__9143\ : InMux
    port map (
            O => \N__48751\,
            I => \N__48748\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__48748\,
            I => \N__48745\
        );

    \I__9141\ : Span4Mux_v
    port map (
            O => \N__48745\,
            I => \N__48742\
        );

    \I__9140\ : Odrv4
    port map (
            O => \N__48742\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_CO\
        );

    \I__9139\ : InMux
    port map (
            O => \N__48739\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17720\
        );

    \I__9138\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48733\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__48733\,
            I => \N__48730\
        );

    \I__9136\ : Sp12to4
    port map (
            O => \N__48730\,
            I => \N__48727\
        );

    \I__9135\ : Span12Mux_v
    port map (
            O => \N__48727\,
            I => \N__48724\
        );

    \I__9134\ : Odrv12
    port map (
            O => \N__48724\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n778\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__48721\,
            I => \N__48718\
        );

    \I__9132\ : InMux
    port map (
            O => \N__48718\,
            I => \N__48715\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__48715\,
            I => \N__48712\
        );

    \I__9130\ : Span4Mux_v
    port map (
            O => \N__48712\,
            I => \N__48709\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__48709\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_CO\
        );

    \I__9128\ : InMux
    port map (
            O => \N__48706\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17721\
        );

    \I__9127\ : CascadeMux
    port map (
            O => \N__48703\,
            I => \N__48700\
        );

    \I__9126\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48697\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__48697\,
            I => \N__48694\
        );

    \I__9124\ : Span12Mux_v
    port map (
            O => \N__48694\,
            I => \N__48691\
        );

    \I__9123\ : Odrv12
    port map (
            O => \N__48691\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_CO\
        );

    \I__9122\ : InMux
    port map (
            O => \N__48688\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17722\
        );

    \I__9121\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48682\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__48682\,
            I => \N__48679\
        );

    \I__9119\ : Odrv12
    port map (
            O => \N__48679\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n786\
        );

    \I__9118\ : InMux
    port map (
            O => \N__48676\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17723\
        );

    \I__9117\ : InMux
    port map (
            O => \N__48673\,
            I => \N__48670\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__48670\,
            I => \N__48667\
        );

    \I__9115\ : Span12Mux_v
    port map (
            O => \N__48667\,
            I => \N__48664\
        );

    \I__9114\ : Odrv12
    port map (
            O => \N__48664\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n790_adj_415\
        );

    \I__9113\ : CascadeMux
    port map (
            O => \N__48661\,
            I => \N__48658\
        );

    \I__9112\ : InMux
    port map (
            O => \N__48658\,
            I => \N__48655\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__48655\,
            I => \N__48652\
        );

    \I__9110\ : Span4Mux_v
    port map (
            O => \N__48652\,
            I => \N__48649\
        );

    \I__9109\ : Odrv4
    port map (
            O => \N__48649\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_CO\
        );

    \I__9108\ : InMux
    port map (
            O => \N__48646\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17724\
        );

    \I__9107\ : InMux
    port map (
            O => \N__48643\,
            I => \N__48640\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__48640\,
            I => \N__48637\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__48637\,
            I => \N__48634\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__48634\,
            I => \N__48631\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__48631\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n794_adj_413\
        );

    \I__9102\ : CascadeMux
    port map (
            O => \N__48628\,
            I => \N__48625\
        );

    \I__9101\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48622\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__48622\,
            I => \N__48619\
        );

    \I__9099\ : Sp12to4
    port map (
            O => \N__48619\,
            I => \N__48616\
        );

    \I__9098\ : Odrv12
    port map (
            O => \N__48616\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_CO\
        );

    \I__9097\ : InMux
    port map (
            O => \N__48613\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17725\
        );

    \I__9096\ : InMux
    port map (
            O => \N__48610\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17711\
        );

    \I__9095\ : InMux
    port map (
            O => \N__48607\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17712\
        );

    \I__9094\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48601\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__48601\,
            I => \N__48598\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__48598\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n746\
        );

    \I__9091\ : InMux
    port map (
            O => \N__48595\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17713\
        );

    \I__9090\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48589\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__48589\,
            I => \N__48586\
        );

    \I__9088\ : Span4Mux_v
    port map (
            O => \N__48586\,
            I => \N__48583\
        );

    \I__9087\ : Odrv4
    port map (
            O => \N__48583\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n750\
        );

    \I__9086\ : CascadeMux
    port map (
            O => \N__48580\,
            I => \N__48577\
        );

    \I__9085\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48574\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__48574\,
            I => \N__48571\
        );

    \I__9083\ : Span4Mux_v
    port map (
            O => \N__48571\,
            I => \N__48568\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__48568\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_CO\
        );

    \I__9081\ : InMux
    port map (
            O => \N__48565\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17714\
        );

    \I__9080\ : InMux
    port map (
            O => \N__48562\,
            I => \N__48559\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__48559\,
            I => \N__48556\
        );

    \I__9078\ : Span4Mux_v
    port map (
            O => \N__48556\,
            I => \N__48553\
        );

    \I__9077\ : Span4Mux_h
    port map (
            O => \N__48553\,
            I => \N__48550\
        );

    \I__9076\ : Odrv4
    port map (
            O => \N__48550\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n754\
        );

    \I__9075\ : CascadeMux
    port map (
            O => \N__48547\,
            I => \N__48544\
        );

    \I__9074\ : InMux
    port map (
            O => \N__48544\,
            I => \N__48541\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__48541\,
            I => \N__48538\
        );

    \I__9072\ : Span4Mux_v
    port map (
            O => \N__48538\,
            I => \N__48535\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__48535\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_CO\
        );

    \I__9070\ : InMux
    port map (
            O => \N__48532\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17715\
        );

    \I__9069\ : InMux
    port map (
            O => \N__48529\,
            I => \N__48526\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__48526\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n758\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__48523\,
            I => \N__48520\
        );

    \I__9066\ : InMux
    port map (
            O => \N__48520\,
            I => \N__48517\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48514\
        );

    \I__9064\ : Span4Mux_h
    port map (
            O => \N__48514\,
            I => \N__48511\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__48511\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_CO\
        );

    \I__9062\ : InMux
    port map (
            O => \N__48508\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17716\
        );

    \I__9061\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48502\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__48502\,
            I => \N__48499\
        );

    \I__9059\ : Odrv4
    port map (
            O => \N__48499\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n762\
        );

    \I__9058\ : CascadeMux
    port map (
            O => \N__48496\,
            I => \N__48493\
        );

    \I__9057\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48490\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__48490\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_CO\
        );

    \I__9055\ : InMux
    port map (
            O => \N__48487\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17717\
        );

    \I__9054\ : CascadeMux
    port map (
            O => \N__48484\,
            I => \N__48481\
        );

    \I__9053\ : InMux
    port map (
            O => \N__48481\,
            I => \N__48478\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__48478\,
            I => \N__48475\
        );

    \I__9051\ : Odrv4
    port map (
            O => \N__48475\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n412\
        );

    \I__9050\ : InMux
    port map (
            O => \N__48472\,
            I => \N__48469\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48466\
        );

    \I__9048\ : Odrv4
    port map (
            O => \N__48466\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n458\
        );

    \I__9047\ : InMux
    port map (
            O => \N__48463\,
            I => \bfn_19_16_0_\
        );

    \I__9046\ : InMux
    port map (
            O => \N__48460\,
            I => \N__48457\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__48457\,
            I => \N__48454\
        );

    \I__9044\ : Odrv12
    port map (
            O => \N__48454\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n461\
        );

    \I__9043\ : InMux
    port map (
            O => \N__48451\,
            I => \N__48448\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__48448\,
            I => \N__48445\
        );

    \I__9041\ : Odrv12
    port map (
            O => \N__48445\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n507\
        );

    \I__9040\ : InMux
    port map (
            O => \N__48442\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17804\
        );

    \I__9039\ : InMux
    port map (
            O => \N__48439\,
            I => \N__48436\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__48436\,
            I => \N__48433\
        );

    \I__9037\ : Odrv4
    port map (
            O => \N__48433\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n510\
        );

    \I__9036\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48427\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__48427\,
            I => \N__48424\
        );

    \I__9034\ : Odrv4
    port map (
            O => \N__48424\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n556_adj_370\
        );

    \I__9033\ : InMux
    port map (
            O => \N__48421\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17805\
        );

    \I__9032\ : InMux
    port map (
            O => \N__48418\,
            I => \N__48415\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__48415\,
            I => \N__48412\
        );

    \I__9030\ : Odrv12
    port map (
            O => \N__48412\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n559_adj_358\
        );

    \I__9029\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48406\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__48406\,
            I => \N__48403\
        );

    \I__9027\ : Odrv12
    port map (
            O => \N__48403\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n605_adj_462\
        );

    \I__9026\ : InMux
    port map (
            O => \N__48400\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17806\
        );

    \I__9025\ : InMux
    port map (
            O => \N__48397\,
            I => \N__48394\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__48394\,
            I => \N__48391\
        );

    \I__9023\ : Odrv4
    port map (
            O => \N__48391\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n608_adj_377\
        );

    \I__9022\ : CascadeMux
    port map (
            O => \N__48388\,
            I => \N__48385\
        );

    \I__9021\ : InMux
    port map (
            O => \N__48385\,
            I => \N__48382\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__48382\,
            I => \N__48379\
        );

    \I__9019\ : Odrv4
    port map (
            O => \N__48379\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n654_adj_456\
        );

    \I__9018\ : InMux
    port map (
            O => \N__48376\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17807\
        );

    \I__9017\ : CascadeMux
    port map (
            O => \N__48373\,
            I => \N__48370\
        );

    \I__9016\ : InMux
    port map (
            O => \N__48370\,
            I => \N__48367\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48364\
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__48364\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n657_adj_360\
        );

    \I__9013\ : CascadeMux
    port map (
            O => \N__48361\,
            I => \N__48358\
        );

    \I__9012\ : InMux
    port map (
            O => \N__48358\,
            I => \N__48355\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__48355\,
            I => \N__48352\
        );

    \I__9010\ : Odrv12
    port map (
            O => \N__48352\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n703_adj_359\
        );

    \I__9009\ : InMux
    port map (
            O => \N__48349\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17808\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__48346\,
            I => \N__48343\
        );

    \I__9007\ : InMux
    port map (
            O => \N__48343\,
            I => \N__48340\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__48340\,
            I => \N__48337\
        );

    \I__9005\ : Odrv12
    port map (
            O => \N__48337\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n706_adj_371\
        );

    \I__9004\ : InMux
    port map (
            O => \N__48334\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17809\
        );

    \I__9003\ : InMux
    port map (
            O => \N__48331\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354\
        );

    \I__9002\ : InMux
    port map (
            O => \N__48328\,
            I => \N__48325\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__48325\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n69\
        );

    \I__9000\ : InMux
    port map (
            O => \N__48322\,
            I => \N__48319\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__48319\,
            I => \N__48316\
        );

    \I__8998\ : Odrv12
    port map (
            O => \N__48316\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n115\
        );

    \I__8997\ : InMux
    port map (
            O => \N__48313\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17796\
        );

    \I__8996\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48307\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__48307\,
            I => \N__48304\
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__48304\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n118\
        );

    \I__8993\ : InMux
    port map (
            O => \N__48301\,
            I => \N__48298\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__48298\,
            I => \N__48295\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__48295\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n164\
        );

    \I__8990\ : InMux
    port map (
            O => \N__48292\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17797\
        );

    \I__8989\ : CascadeMux
    port map (
            O => \N__48289\,
            I => \N__48286\
        );

    \I__8988\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48283\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__48283\,
            I => \N__48280\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__48280\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n167\
        );

    \I__8985\ : InMux
    port map (
            O => \N__48277\,
            I => \N__48274\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__48274\,
            I => \N__48271\
        );

    \I__8983\ : Odrv12
    port map (
            O => \N__48271\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n213\
        );

    \I__8982\ : InMux
    port map (
            O => \N__48268\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17798\
        );

    \I__8981\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48262\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__48262\,
            I => \N__48259\
        );

    \I__8979\ : Odrv4
    port map (
            O => \N__48259\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n216\
        );

    \I__8978\ : InMux
    port map (
            O => \N__48256\,
            I => \N__48253\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__48253\,
            I => \N__48250\
        );

    \I__8976\ : Odrv4
    port map (
            O => \N__48250\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n262_adj_425\
        );

    \I__8975\ : InMux
    port map (
            O => \N__48247\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17799\
        );

    \I__8974\ : InMux
    port map (
            O => \N__48244\,
            I => \N__48241\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__48241\,
            I => \N__48238\
        );

    \I__8972\ : Odrv4
    port map (
            O => \N__48238\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n265\
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__48235\,
            I => \N__48232\
        );

    \I__8970\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48229\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__48229\,
            I => \N__48226\
        );

    \I__8968\ : Odrv4
    port map (
            O => \N__48226\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n311_adj_422\
        );

    \I__8967\ : InMux
    port map (
            O => \N__48223\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17800\
        );

    \I__8966\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48217\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__48217\,
            I => \N__48214\
        );

    \I__8964\ : Odrv12
    port map (
            O => \N__48214\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n314_adj_401\
        );

    \I__8963\ : CascadeMux
    port map (
            O => \N__48211\,
            I => \N__48208\
        );

    \I__8962\ : InMux
    port map (
            O => \N__48208\,
            I => \N__48205\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__48205\,
            I => \N__48202\
        );

    \I__8960\ : Odrv12
    port map (
            O => \N__48202\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n360\
        );

    \I__8959\ : InMux
    port map (
            O => \N__48199\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17801\
        );

    \I__8958\ : InMux
    port map (
            O => \N__48196\,
            I => \N__48193\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__48193\,
            I => \N__48190\
        );

    \I__8956\ : Odrv4
    port map (
            O => \N__48190\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n363_adj_380\
        );

    \I__8955\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48184\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__48184\,
            I => \N__48181\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__48181\,
            I => \N__48178\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__48178\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n409\
        );

    \I__8951\ : InMux
    port map (
            O => \N__48175\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17802\
        );

    \I__8950\ : InMux
    port map (
            O => \N__48172\,
            I => \N__48169\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__48169\,
            I => \N__48166\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__48166\,
            I => \N__48163\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__48163\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n366_adj_426\
        );

    \I__8946\ : InMux
    port map (
            O => \N__48160\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17817\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__48157\,
            I => \N__48154\
        );

    \I__8944\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48151\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__48151\,
            I => \N__48148\
        );

    \I__8942\ : Odrv4
    port map (
            O => \N__48148\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n415\
        );

    \I__8941\ : InMux
    port map (
            O => \N__48145\,
            I => \bfn_19_14_0_\
        );

    \I__8940\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48139\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__48139\,
            I => \N__48136\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__48136\,
            I => \N__48133\
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__48133\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n464_adj_423\
        );

    \I__8936\ : InMux
    port map (
            O => \N__48130\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17819\
        );

    \I__8935\ : InMux
    port map (
            O => \N__48127\,
            I => \N__48124\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__48124\,
            I => \N__48121\
        );

    \I__8933\ : Odrv4
    port map (
            O => \N__48121\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n513_adj_412\
        );

    \I__8932\ : InMux
    port map (
            O => \N__48118\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17820\
        );

    \I__8931\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48112\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__48112\,
            I => \N__48109\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__48109\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n562_adj_378\
        );

    \I__8928\ : InMux
    port map (
            O => \N__48106\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17821\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__48103\,
            I => \N__48100\
        );

    \I__8926\ : InMux
    port map (
            O => \N__48100\,
            I => \N__48097\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__48097\,
            I => \N__48094\
        );

    \I__8924\ : Odrv4
    port map (
            O => \N__48094\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n611_adj_373\
        );

    \I__8923\ : InMux
    port map (
            O => \N__48091\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17822\
        );

    \I__8922\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48085\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__48085\,
            I => \N__48082\
        );

    \I__8920\ : Span4Mux_v
    port map (
            O => \N__48082\,
            I => \N__48079\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__48079\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n660_adj_372\
        );

    \I__8918\ : InMux
    port map (
            O => \N__48076\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17823\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__48073\,
            I => \N__48070\
        );

    \I__8916\ : InMux
    port map (
            O => \N__48070\,
            I => \N__48067\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__48067\,
            I => \N__48064\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__48064\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n709\
        );

    \I__8913\ : InMux
    port map (
            O => \N__48061\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17824\
        );

    \I__8912\ : InMux
    port map (
            O => \N__48058\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n763\
        );

    \I__8911\ : InMux
    port map (
            O => \N__48055\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421\
        );

    \I__8910\ : CascadeMux
    port map (
            O => \N__48052\,
            I => \N__48049\
        );

    \I__8909\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48046\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__48046\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n72\
        );

    \I__8907\ : InMux
    port map (
            O => \N__48043\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17811\
        );

    \I__8906\ : InMux
    port map (
            O => \N__48040\,
            I => \N__48037\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__48037\,
            I => \N__48034\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__48034\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n121\
        );

    \I__8903\ : InMux
    port map (
            O => \N__48031\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17812\
        );

    \I__8902\ : InMux
    port map (
            O => \N__48028\,
            I => \N__48025\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__48025\,
            I => \N__48022\
        );

    \I__8900\ : Odrv4
    port map (
            O => \N__48022\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n170\
        );

    \I__8899\ : InMux
    port map (
            O => \N__48019\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17813\
        );

    \I__8898\ : InMux
    port map (
            O => \N__48016\,
            I => \N__48013\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__48013\,
            I => \N__48010\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__48010\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n219\
        );

    \I__8895\ : InMux
    port map (
            O => \N__48007\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17814\
        );

    \I__8894\ : InMux
    port map (
            O => \N__48004\,
            I => \N__48001\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__48001\,
            I => \N__47998\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__47998\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n268_adj_437\
        );

    \I__8891\ : InMux
    port map (
            O => \N__47995\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17815\
        );

    \I__8890\ : CascadeMux
    port map (
            O => \N__47992\,
            I => \N__47989\
        );

    \I__8889\ : InMux
    port map (
            O => \N__47989\,
            I => \N__47986\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__47986\,
            I => \N__47983\
        );

    \I__8887\ : Odrv4
    port map (
            O => \N__47983\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n317_adj_428\
        );

    \I__8886\ : InMux
    port map (
            O => \N__47980\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17816\
        );

    \I__8885\ : InMux
    port map (
            O => \N__47977\,
            I => \N__47974\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__47974\,
            I => \N__47971\
        );

    \I__8883\ : Odrv12
    port map (
            O => \N__47971\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n335\
        );

    \I__8882\ : InMux
    port map (
            O => \N__47968\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17917\
        );

    \I__8881\ : InMux
    port map (
            O => \N__47965\,
            I => \N__47962\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__47962\,
            I => \N__47959\
        );

    \I__8879\ : Odrv4
    port map (
            O => \N__47959\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n384\
        );

    \I__8878\ : InMux
    port map (
            O => \N__47956\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17918\
        );

    \I__8877\ : InMux
    port map (
            O => \N__47953\,
            I => \N__47950\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__47950\,
            I => \N__47947\
        );

    \I__8875\ : Odrv12
    port map (
            O => \N__47947\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n433\
        );

    \I__8874\ : InMux
    port map (
            O => \N__47944\,
            I => \bfn_19_12_0_\
        );

    \I__8873\ : InMux
    port map (
            O => \N__47941\,
            I => \N__47938\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__47938\,
            I => \N__47935\
        );

    \I__8871\ : Odrv4
    port map (
            O => \N__47935\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n482\
        );

    \I__8870\ : InMux
    port map (
            O => \N__47932\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17920\
        );

    \I__8869\ : InMux
    port map (
            O => \N__47929\,
            I => \N__47926\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__47926\,
            I => \N__47923\
        );

    \I__8867\ : Odrv4
    port map (
            O => \N__47923\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n531\
        );

    \I__8866\ : InMux
    port map (
            O => \N__47920\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17921\
        );

    \I__8865\ : InMux
    port map (
            O => \N__47917\,
            I => \N__47914\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__47914\,
            I => \N__47911\
        );

    \I__8863\ : Odrv12
    port map (
            O => \N__47911\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n580\
        );

    \I__8862\ : InMux
    port map (
            O => \N__47908\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17922\
        );

    \I__8861\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47902\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__47902\,
            I => \N__47899\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__47899\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n629\
        );

    \I__8858\ : InMux
    port map (
            O => \N__47896\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17923\
        );

    \I__8857\ : CascadeMux
    port map (
            O => \N__47893\,
            I => \N__47890\
        );

    \I__8856\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47887\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__47887\,
            I => \N__47884\
        );

    \I__8854\ : Span4Mux_v
    port map (
            O => \N__47884\,
            I => \N__47881\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__47881\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n678\
        );

    \I__8852\ : InMux
    port map (
            O => \N__47878\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17924\
        );

    \I__8851\ : CascadeMux
    port map (
            O => \N__47875\,
            I => \N__47872\
        );

    \I__8850\ : InMux
    port map (
            O => \N__47872\,
            I => \N__47869\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__47869\,
            I => \N__47866\
        );

    \I__8848\ : Odrv4
    port map (
            O => \N__47866\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n727\
        );

    \I__8847\ : InMux
    port map (
            O => \N__47863\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17925\
        );

    \I__8846\ : CascadeMux
    port map (
            O => \N__47860\,
            I => \N__47857\
        );

    \I__8845\ : InMux
    port map (
            O => \N__47857\,
            I => \N__47854\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__47854\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n730\
        );

    \I__8843\ : InMux
    port map (
            O => \N__47851\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17940\
        );

    \I__8842\ : InMux
    port map (
            O => \N__47848\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416\
        );

    \I__8841\ : CascadeMux
    port map (
            O => \N__47845\,
            I => \N__47842\
        );

    \I__8840\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47839\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__47839\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n90_adj_420\
        );

    \I__8838\ : InMux
    port map (
            O => \N__47836\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17912\
        );

    \I__8837\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47830\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__47830\,
            I => \N__47827\
        );

    \I__8835\ : Odrv4
    port map (
            O => \N__47827\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n139_adj_419\
        );

    \I__8834\ : InMux
    port map (
            O => \N__47824\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17913\
        );

    \I__8833\ : InMux
    port map (
            O => \N__47821\,
            I => \N__47818\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__47818\,
            I => \N__47815\
        );

    \I__8831\ : Odrv12
    port map (
            O => \N__47815\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n188_adj_418\
        );

    \I__8830\ : InMux
    port map (
            O => \N__47812\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17914\
        );

    \I__8829\ : InMux
    port map (
            O => \N__47809\,
            I => \N__47806\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__47806\,
            I => \N__47803\
        );

    \I__8827\ : Odrv4
    port map (
            O => \N__47803\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n237_adj_417\
        );

    \I__8826\ : InMux
    port map (
            O => \N__47800\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17915\
        );

    \I__8825\ : InMux
    port map (
            O => \N__47797\,
            I => \N__47794\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__47794\,
            I => \N__47791\
        );

    \I__8823\ : Odrv4
    port map (
            O => \N__47791\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n286\
        );

    \I__8822\ : InMux
    port map (
            O => \N__47788\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17916\
        );

    \I__8821\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47782\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__47782\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n289\
        );

    \I__8819\ : InMux
    port map (
            O => \N__47779\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17931\
        );

    \I__8818\ : InMux
    port map (
            O => \N__47776\,
            I => \N__47773\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__47773\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n338\
        );

    \I__8816\ : InMux
    port map (
            O => \N__47770\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17932\
        );

    \I__8815\ : InMux
    port map (
            O => \N__47767\,
            I => \N__47764\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__47764\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n387\
        );

    \I__8813\ : InMux
    port map (
            O => \N__47761\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17933\
        );

    \I__8812\ : CascadeMux
    port map (
            O => \N__47758\,
            I => \N__47755\
        );

    \I__8811\ : InMux
    port map (
            O => \N__47755\,
            I => \N__47752\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__47752\,
            I => \N__47749\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__47749\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n436\
        );

    \I__8808\ : InMux
    port map (
            O => \N__47746\,
            I => \bfn_19_10_0_\
        );

    \I__8807\ : InMux
    port map (
            O => \N__47743\,
            I => \N__47740\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__47740\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n485\
        );

    \I__8805\ : InMux
    port map (
            O => \N__47737\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17935\
        );

    \I__8804\ : InMux
    port map (
            O => \N__47734\,
            I => \N__47731\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__47731\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n534\
        );

    \I__8802\ : InMux
    port map (
            O => \N__47728\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17936\
        );

    \I__8801\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47722\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__47722\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n583\
        );

    \I__8799\ : InMux
    port map (
            O => \N__47719\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17937\
        );

    \I__8798\ : InMux
    port map (
            O => \N__47716\,
            I => \N__47713\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__47713\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n632\
        );

    \I__8796\ : InMux
    port map (
            O => \N__47710\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17938\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__47707\,
            I => \N__47704\
        );

    \I__8794\ : InMux
    port map (
            O => \N__47704\,
            I => \N__47701\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__47701\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n681\
        );

    \I__8792\ : InMux
    port map (
            O => \N__47698\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17939\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__47695\,
            I => \N__47692\
        );

    \I__8790\ : InMux
    port map (
            O => \N__47692\,
            I => \N__47689\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__47689\,
            I => \N__47686\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__47686\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n663\
        );

    \I__8787\ : InMux
    port map (
            O => \N__47683\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17638\
        );

    \I__8786\ : InMux
    port map (
            O => \N__47680\,
            I => \N__47676\
        );

    \I__8785\ : InMux
    port map (
            O => \N__47679\,
            I => \N__47673\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__47676\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n765\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__47673\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n765\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__47668\,
            I => \N__47665\
        );

    \I__8781\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47662\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__47662\,
            I => \N__47659\
        );

    \I__8779\ : Odrv4
    port map (
            O => \N__47659\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n712\
        );

    \I__8778\ : InMux
    port map (
            O => \N__47656\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17639\
        );

    \I__8777\ : InMux
    port map (
            O => \N__47653\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382\
        );

    \I__8776\ : InMux
    port map (
            O => \N__47650\,
            I => \N__47647\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__47647\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n93\
        );

    \I__8774\ : InMux
    port map (
            O => \N__47644\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17927\
        );

    \I__8773\ : InMux
    port map (
            O => \N__47641\,
            I => \N__47638\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__47638\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n142_adj_414\
        );

    \I__8771\ : InMux
    port map (
            O => \N__47635\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17928\
        );

    \I__8770\ : CascadeMux
    port map (
            O => \N__47632\,
            I => \N__47629\
        );

    \I__8769\ : InMux
    port map (
            O => \N__47629\,
            I => \N__47626\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__47626\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n191\
        );

    \I__8767\ : InMux
    port map (
            O => \N__47623\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17929\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__47620\,
            I => \N__47617\
        );

    \I__8765\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47614\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__47614\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n240\
        );

    \I__8763\ : InMux
    port map (
            O => \N__47611\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17930\
        );

    \I__8762\ : InMux
    port map (
            O => \N__47608\,
            I => \N__47605\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__47605\,
            I => \N__47602\
        );

    \I__8760\ : Odrv4
    port map (
            O => \N__47602\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n222\
        );

    \I__8759\ : InMux
    port map (
            O => \N__47599\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17629\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__47596\,
            I => \N__47593\
        );

    \I__8757\ : InMux
    port map (
            O => \N__47593\,
            I => \N__47590\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__47590\,
            I => \N__47587\
        );

    \I__8755\ : Odrv4
    port map (
            O => \N__47587\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n271\
        );

    \I__8754\ : InMux
    port map (
            O => \N__47584\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17630\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__47581\,
            I => \N__47578\
        );

    \I__8752\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47575\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__47575\,
            I => \N__47572\
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__47572\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n320\
        );

    \I__8749\ : InMux
    port map (
            O => \N__47569\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17631\
        );

    \I__8748\ : InMux
    port map (
            O => \N__47566\,
            I => \N__47563\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__47563\,
            I => \N__47560\
        );

    \I__8746\ : Odrv4
    port map (
            O => \N__47560\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n369\
        );

    \I__8745\ : InMux
    port map (
            O => \N__47557\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17632\
        );

    \I__8744\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47551\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__47551\,
            I => \N__47548\
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__47548\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n418\
        );

    \I__8741\ : InMux
    port map (
            O => \N__47545\,
            I => \bfn_19_8_0_\
        );

    \I__8740\ : CascadeMux
    port map (
            O => \N__47542\,
            I => \N__47539\
        );

    \I__8739\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47536\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__47536\,
            I => \N__47533\
        );

    \I__8737\ : Odrv12
    port map (
            O => \N__47533\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n467\
        );

    \I__8736\ : InMux
    port map (
            O => \N__47530\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17634\
        );

    \I__8735\ : InMux
    port map (
            O => \N__47527\,
            I => \N__47524\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__47524\,
            I => \N__47521\
        );

    \I__8733\ : Odrv4
    port map (
            O => \N__47521\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n516\
        );

    \I__8732\ : InMux
    port map (
            O => \N__47518\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17635\
        );

    \I__8731\ : CascadeMux
    port map (
            O => \N__47515\,
            I => \N__47512\
        );

    \I__8730\ : InMux
    port map (
            O => \N__47512\,
            I => \N__47509\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__47509\,
            I => \N__47506\
        );

    \I__8728\ : Odrv12
    port map (
            O => \N__47506\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n565\
        );

    \I__8727\ : InMux
    port map (
            O => \N__47503\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17636\
        );

    \I__8726\ : InMux
    port map (
            O => \N__47500\,
            I => \N__47497\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__47497\,
            I => \N__47494\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__47494\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n614\
        );

    \I__8723\ : InMux
    port map (
            O => \N__47491\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17637\
        );

    \I__8722\ : InMux
    port map (
            O => \N__47488\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17651\
        );

    \I__8721\ : InMux
    port map (
            O => \N__47485\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17652\
        );

    \I__8720\ : InMux
    port map (
            O => \N__47482\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17653\
        );

    \I__8719\ : CascadeMux
    port map (
            O => \N__47479\,
            I => \N__47476\
        );

    \I__8718\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47473\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__47473\,
            I => \N__47469\
        );

    \I__8716\ : InMux
    port map (
            O => \N__47472\,
            I => \N__47466\
        );

    \I__8715\ : Span4Mux_v
    port map (
            O => \N__47469\,
            I => \N__47463\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__47466\,
            I => \N__47460\
        );

    \I__8713\ : Odrv4
    port map (
            O => \N__47463\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n769\
        );

    \I__8712\ : Odrv12
    port map (
            O => \N__47460\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n769\
        );

    \I__8711\ : InMux
    port map (
            O => \N__47455\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17654\
        );

    \I__8710\ : InMux
    port map (
            O => \N__47452\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n771\
        );

    \I__8709\ : CascadeMux
    port map (
            O => \N__47449\,
            I => \N__47446\
        );

    \I__8708\ : InMux
    port map (
            O => \N__47446\,
            I => \N__47443\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__47443\,
            I => \N__47440\
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__47440\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n75_adj_510\
        );

    \I__8705\ : InMux
    port map (
            O => \N__47437\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17626\
        );

    \I__8704\ : InMux
    port map (
            O => \N__47434\,
            I => \N__47431\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__47431\,
            I => \N__47428\
        );

    \I__8702\ : Odrv4
    port map (
            O => \N__47428\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n124\
        );

    \I__8701\ : InMux
    port map (
            O => \N__47425\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17627\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__47422\,
            I => \N__47419\
        );

    \I__8699\ : InMux
    port map (
            O => \N__47419\,
            I => \N__47416\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__47416\,
            I => \N__47413\
        );

    \I__8697\ : Odrv12
    port map (
            O => \N__47413\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n173\
        );

    \I__8696\ : InMux
    port map (
            O => \N__47410\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17628\
        );

    \I__8695\ : InMux
    port map (
            O => \N__47407\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17642\
        );

    \I__8694\ : InMux
    port map (
            O => \N__47404\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17643\
        );

    \I__8693\ : InMux
    port map (
            O => \N__47401\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17644\
        );

    \I__8692\ : InMux
    port map (
            O => \N__47398\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17645\
        );

    \I__8691\ : InMux
    port map (
            O => \N__47395\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17646\
        );

    \I__8690\ : InMux
    port map (
            O => \N__47392\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17647\
        );

    \I__8689\ : InMux
    port map (
            O => \N__47389\,
            I => \bfn_19_6_0_\
        );

    \I__8688\ : InMux
    port map (
            O => \N__47386\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17649\
        );

    \I__8687\ : InMux
    port map (
            O => \N__47383\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17650\
        );

    \I__8686\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47377\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__47377\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n534\
        );

    \I__8684\ : InMux
    port map (
            O => \N__47374\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18363\
        );

    \I__8683\ : InMux
    port map (
            O => \N__47371\,
            I => \N__47368\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__47368\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n583\
        );

    \I__8681\ : InMux
    port map (
            O => \N__47365\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18364\
        );

    \I__8680\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47359\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__47359\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n632\
        );

    \I__8678\ : InMux
    port map (
            O => \N__47356\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18365\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__47353\,
            I => \N__47350\
        );

    \I__8676\ : InMux
    port map (
            O => \N__47350\,
            I => \N__47347\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__47347\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n681\
        );

    \I__8674\ : InMux
    port map (
            O => \N__47344\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18366\
        );

    \I__8673\ : InMux
    port map (
            O => \N__47341\,
            I => \N__47338\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__47338\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n730\
        );

    \I__8671\ : InMux
    port map (
            O => \N__47335\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18367\
        );

    \I__8670\ : InMux
    port map (
            O => \N__47332\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n791\
        );

    \I__8669\ : InMux
    port map (
            O => \N__47329\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17641\
        );

    \I__8668\ : CascadeMux
    port map (
            O => \N__47326\,
            I => \N__47323\
        );

    \I__8667\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47320\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__47320\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n93\
        );

    \I__8665\ : InMux
    port map (
            O => \N__47317\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18354\
        );

    \I__8664\ : CascadeMux
    port map (
            O => \N__47314\,
            I => \N__47311\
        );

    \I__8663\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47308\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__47308\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n142\
        );

    \I__8661\ : InMux
    port map (
            O => \N__47305\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18355\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__47302\,
            I => \N__47299\
        );

    \I__8659\ : InMux
    port map (
            O => \N__47299\,
            I => \N__47296\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__47296\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n191\
        );

    \I__8657\ : InMux
    port map (
            O => \N__47293\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18356\
        );

    \I__8656\ : InMux
    port map (
            O => \N__47290\,
            I => \N__47287\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__47287\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n240\
        );

    \I__8654\ : InMux
    port map (
            O => \N__47284\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18357\
        );

    \I__8653\ : InMux
    port map (
            O => \N__47281\,
            I => \N__47278\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__47278\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n289\
        );

    \I__8651\ : InMux
    port map (
            O => \N__47275\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18358\
        );

    \I__8650\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47269\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__47269\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n338\
        );

    \I__8648\ : InMux
    port map (
            O => \N__47266\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18359\
        );

    \I__8647\ : InMux
    port map (
            O => \N__47263\,
            I => \N__47260\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__47260\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n387\
        );

    \I__8645\ : InMux
    port map (
            O => \N__47257\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18360\
        );

    \I__8644\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47251\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__47251\,
            I => \N__47248\
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__47248\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n436\
        );

    \I__8641\ : InMux
    port map (
            O => \N__47245\,
            I => \bfn_18_27_0_\
        );

    \I__8640\ : InMux
    port map (
            O => \N__47242\,
            I => \N__47239\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__47239\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n485\
        );

    \I__8638\ : InMux
    port map (
            O => \N__47236\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18362\
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__47233\,
            I => \N__47230\
        );

    \I__8636\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47227\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__47227\,
            I => \N__47224\
        );

    \I__8634\ : Span12Mux_h
    port map (
            O => \N__47224\,
            I => \N__47221\
        );

    \I__8633\ : Odrv12
    port map (
            O => \N__47221\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_24\
        );

    \I__8632\ : InMux
    port map (
            O => \N__47218\,
            I => \bfn_18_25_0_\
        );

    \I__8631\ : InMux
    port map (
            O => \N__47215\,
            I => \N__47212\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47209\
        );

    \I__8629\ : Span12Mux_s9_v
    port map (
            O => \N__47209\,
            I => \N__47206\
        );

    \I__8628\ : Odrv12
    port map (
            O => \N__47206\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_25\
        );

    \I__8627\ : InMux
    port map (
            O => \N__47203\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15907\
        );

    \I__8626\ : CascadeMux
    port map (
            O => \N__47200\,
            I => \N__47197\
        );

    \I__8625\ : InMux
    port map (
            O => \N__47197\,
            I => \N__47194\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__47194\,
            I => \N__47191\
        );

    \I__8623\ : Span4Mux_v
    port map (
            O => \N__47191\,
            I => \N__47188\
        );

    \I__8622\ : Sp12to4
    port map (
            O => \N__47188\,
            I => \N__47185\
        );

    \I__8621\ : Odrv12
    port map (
            O => \N__47185\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_26\
        );

    \I__8620\ : InMux
    port map (
            O => \N__47182\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15908\
        );

    \I__8619\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47176\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__47176\,
            I => \N__47173\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__47173\,
            I => \N__47170\
        );

    \I__8616\ : Span4Mux_h
    port map (
            O => \N__47170\,
            I => \N__47167\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__47167\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_27\
        );

    \I__8614\ : InMux
    port map (
            O => \N__47164\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15909\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__47161\,
            I => \N__47158\
        );

    \I__8612\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47155\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__47155\,
            I => \N__47152\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__47152\,
            I => \N__47149\
        );

    \I__8609\ : Span4Mux_h
    port map (
            O => \N__47149\,
            I => \N__47146\
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__47146\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_28\
        );

    \I__8607\ : InMux
    port map (
            O => \N__47143\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15910\
        );

    \I__8606\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47137\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47134\
        );

    \I__8604\ : Span4Mux_v
    port map (
            O => \N__47134\,
            I => \N__47131\
        );

    \I__8603\ : Span4Mux_h
    port map (
            O => \N__47131\,
            I => \N__47128\
        );

    \I__8602\ : Odrv4
    port map (
            O => \N__47128\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_29\
        );

    \I__8601\ : InMux
    port map (
            O => \N__47125\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15911\
        );

    \I__8600\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47119\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__47119\,
            I => \N__47116\
        );

    \I__8598\ : Span4Mux_v
    port map (
            O => \N__47116\,
            I => \N__47113\
        );

    \I__8597\ : Span4Mux_h
    port map (
            O => \N__47113\,
            I => \N__47110\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__47110\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_30\
        );

    \I__8595\ : InMux
    port map (
            O => \N__47107\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15912\
        );

    \I__8594\ : CascadeMux
    port map (
            O => \N__47104\,
            I => \N__47101\
        );

    \I__8593\ : InMux
    port map (
            O => \N__47101\,
            I => \N__47098\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__47098\,
            I => \N__47095\
        );

    \I__8591\ : Span12Mux_h
    port map (
            O => \N__47095\,
            I => \N__47092\
        );

    \I__8590\ : Odrv12
    port map (
            O => \N__47092\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_15\
        );

    \I__8589\ : InMux
    port map (
            O => \N__47089\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15897\
        );

    \I__8588\ : InMux
    port map (
            O => \N__47086\,
            I => \N__47083\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__47083\,
            I => \N__47080\
        );

    \I__8586\ : Span12Mux_h
    port map (
            O => \N__47080\,
            I => \N__47077\
        );

    \I__8585\ : Odrv12
    port map (
            O => \N__47077\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_16\
        );

    \I__8584\ : InMux
    port map (
            O => \N__47074\,
            I => \bfn_18_24_0_\
        );

    \I__8583\ : CascadeMux
    port map (
            O => \N__47071\,
            I => \N__47068\
        );

    \I__8582\ : InMux
    port map (
            O => \N__47068\,
            I => \N__47065\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__47065\,
            I => \N__47062\
        );

    \I__8580\ : Span4Mux_v
    port map (
            O => \N__47062\,
            I => \N__47059\
        );

    \I__8579\ : Span4Mux_h
    port map (
            O => \N__47059\,
            I => \N__47056\
        );

    \I__8578\ : Odrv4
    port map (
            O => \N__47056\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_17\
        );

    \I__8577\ : InMux
    port map (
            O => \N__47053\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15899\
        );

    \I__8576\ : CascadeMux
    port map (
            O => \N__47050\,
            I => \N__47047\
        );

    \I__8575\ : InMux
    port map (
            O => \N__47047\,
            I => \N__47044\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__47044\,
            I => \N__47041\
        );

    \I__8573\ : Span4Mux_v
    port map (
            O => \N__47041\,
            I => \N__47038\
        );

    \I__8572\ : Span4Mux_h
    port map (
            O => \N__47038\,
            I => \N__47035\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__47035\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_18\
        );

    \I__8570\ : InMux
    port map (
            O => \N__47032\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15900\
        );

    \I__8569\ : InMux
    port map (
            O => \N__47029\,
            I => \N__47026\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__47026\,
            I => \N__47023\
        );

    \I__8567\ : Span4Mux_h
    port map (
            O => \N__47023\,
            I => \N__47020\
        );

    \I__8566\ : Span4Mux_h
    port map (
            O => \N__47020\,
            I => \N__47017\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__47017\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_19\
        );

    \I__8564\ : InMux
    port map (
            O => \N__47014\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15901\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__47011\,
            I => \N__47008\
        );

    \I__8562\ : InMux
    port map (
            O => \N__47008\,
            I => \N__47005\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__47005\,
            I => \N__47002\
        );

    \I__8560\ : Span4Mux_v
    port map (
            O => \N__47002\,
            I => \N__46999\
        );

    \I__8559\ : Span4Mux_h
    port map (
            O => \N__46999\,
            I => \N__46996\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__46996\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_20\
        );

    \I__8557\ : InMux
    port map (
            O => \N__46993\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15902\
        );

    \I__8556\ : CascadeMux
    port map (
            O => \N__46990\,
            I => \N__46987\
        );

    \I__8555\ : InMux
    port map (
            O => \N__46987\,
            I => \N__46984\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__46984\,
            I => \N__46981\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__46981\,
            I => \N__46978\
        );

    \I__8552\ : Span4Mux_h
    port map (
            O => \N__46978\,
            I => \N__46975\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__46975\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_21\
        );

    \I__8550\ : InMux
    port map (
            O => \N__46972\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15903\
        );

    \I__8549\ : CascadeMux
    port map (
            O => \N__46969\,
            I => \N__46966\
        );

    \I__8548\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46963\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__46963\,
            I => \N__46960\
        );

    \I__8546\ : Span4Mux_v
    port map (
            O => \N__46960\,
            I => \N__46957\
        );

    \I__8545\ : Span4Mux_h
    port map (
            O => \N__46957\,
            I => \N__46954\
        );

    \I__8544\ : Odrv4
    port map (
            O => \N__46954\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_22\
        );

    \I__8543\ : InMux
    port map (
            O => \N__46951\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15904\
        );

    \I__8542\ : CascadeMux
    port map (
            O => \N__46948\,
            I => \N__46945\
        );

    \I__8541\ : InMux
    port map (
            O => \N__46945\,
            I => \N__46942\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__46942\,
            I => \N__46939\
        );

    \I__8539\ : Span4Mux_v
    port map (
            O => \N__46939\,
            I => \N__46936\
        );

    \I__8538\ : Span4Mux_h
    port map (
            O => \N__46936\,
            I => \N__46933\
        );

    \I__8537\ : Odrv4
    port map (
            O => \N__46933\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_23\
        );

    \I__8536\ : InMux
    port map (
            O => \N__46930\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15905\
        );

    \I__8535\ : CascadeMux
    port map (
            O => \N__46927\,
            I => \N__46924\
        );

    \I__8534\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46921\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__46921\,
            I => \N__46918\
        );

    \I__8532\ : Span4Mux_h
    port map (
            O => \N__46918\,
            I => \N__46915\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__46915\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_7\
        );

    \I__8530\ : InMux
    port map (
            O => \N__46912\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15889\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__46909\,
            I => \N__46906\
        );

    \I__8528\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46903\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__46903\,
            I => \N__46900\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__46900\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_8\
        );

    \I__8525\ : InMux
    port map (
            O => \N__46897\,
            I => \bfn_18_23_0_\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__46894\,
            I => \N__46891\
        );

    \I__8523\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46888\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46885\
        );

    \I__8521\ : Span4Mux_v
    port map (
            O => \N__46885\,
            I => \N__46882\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__46882\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_9\
        );

    \I__8519\ : InMux
    port map (
            O => \N__46879\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15891\
        );

    \I__8518\ : CascadeMux
    port map (
            O => \N__46876\,
            I => \N__46873\
        );

    \I__8517\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46870\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__46870\,
            I => \N__46867\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__46867\,
            I => \N__46864\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__46864\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_10\
        );

    \I__8513\ : InMux
    port map (
            O => \N__46861\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15892\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__46858\,
            I => \N__46855\
        );

    \I__8511\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46852\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__46852\,
            I => \N__46849\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__46849\,
            I => \N__46846\
        );

    \I__8508\ : Odrv4
    port map (
            O => \N__46846\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_11\
        );

    \I__8507\ : InMux
    port map (
            O => \N__46843\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15893\
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__46840\,
            I => \N__46837\
        );

    \I__8505\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46834\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__46834\,
            I => \N__46831\
        );

    \I__8503\ : Span4Mux_h
    port map (
            O => \N__46831\,
            I => \N__46828\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__46828\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_12\
        );

    \I__8501\ : InMux
    port map (
            O => \N__46825\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15894\
        );

    \I__8500\ : CascadeMux
    port map (
            O => \N__46822\,
            I => \N__46819\
        );

    \I__8499\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46816\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__46816\,
            I => \N__46813\
        );

    \I__8497\ : Span4Mux_h
    port map (
            O => \N__46813\,
            I => \N__46810\
        );

    \I__8496\ : Odrv4
    port map (
            O => \N__46810\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_13\
        );

    \I__8495\ : InMux
    port map (
            O => \N__46807\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15895\
        );

    \I__8494\ : InMux
    port map (
            O => \N__46804\,
            I => \N__46801\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__46801\,
            I => \N__46798\
        );

    \I__8492\ : Span4Mux_h
    port map (
            O => \N__46798\,
            I => \N__46795\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__46795\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_14\
        );

    \I__8490\ : InMux
    port map (
            O => \N__46792\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15896\
        );

    \I__8489\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46786\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__46786\,
            I => \N__46782\
        );

    \I__8487\ : InMux
    port map (
            O => \N__46785\,
            I => \N__46779\
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__46782\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__46779\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28\
        );

    \I__8484\ : InMux
    port map (
            O => \N__46774\,
            I => \N__46770\
        );

    \I__8483\ : InMux
    port map (
            O => \N__46773\,
            I => \N__46767\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__46770\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20174\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__46767\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20174\
        );

    \I__8480\ : CascadeMux
    port map (
            O => \N__46762\,
            I => \N__46759\
        );

    \I__8479\ : InMux
    port map (
            O => \N__46759\,
            I => \N__46756\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__46756\,
            I => \N__46753\
        );

    \I__8477\ : Span4Mux_v
    port map (
            O => \N__46753\,
            I => \N__46750\
        );

    \I__8476\ : Odrv4
    port map (
            O => \N__46750\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_1\
        );

    \I__8475\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46743\
        );

    \I__8474\ : InMux
    port map (
            O => \N__46746\,
            I => \N__46740\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__46743\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__46740\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2\
        );

    \I__8471\ : InMux
    port map (
            O => \N__46735\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15883\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__46732\,
            I => \N__46729\
        );

    \I__8469\ : InMux
    port map (
            O => \N__46729\,
            I => \N__46726\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__46726\,
            I => \N__46723\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__46723\,
            I => \N__46720\
        );

    \I__8466\ : Odrv4
    port map (
            O => \N__46720\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_2\
        );

    \I__8465\ : CascadeMux
    port map (
            O => \N__46717\,
            I => \N__46713\
        );

    \I__8464\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46710\
        );

    \I__8463\ : InMux
    port map (
            O => \N__46713\,
            I => \N__46707\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__46710\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__46707\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3\
        );

    \I__8460\ : InMux
    port map (
            O => \N__46702\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15884\
        );

    \I__8459\ : InMux
    port map (
            O => \N__46699\,
            I => \N__46696\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__46696\,
            I => \N__46693\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__46693\,
            I => \N__46690\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__46690\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_3\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__46687\,
            I => \N__46684\
        );

    \I__8454\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46680\
        );

    \I__8453\ : InMux
    port map (
            O => \N__46683\,
            I => \N__46677\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__46680\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__46677\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4\
        );

    \I__8450\ : InMux
    port map (
            O => \N__46672\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15885\
        );

    \I__8449\ : CascadeMux
    port map (
            O => \N__46669\,
            I => \N__46666\
        );

    \I__8448\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46663\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__46663\,
            I => \N__46660\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__46660\,
            I => \N__46657\
        );

    \I__8445\ : Span4Mux_v
    port map (
            O => \N__46657\,
            I => \N__46654\
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__46654\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_4\
        );

    \I__8443\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46647\
        );

    \I__8442\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46644\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__46647\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__46644\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5\
        );

    \I__8439\ : InMux
    port map (
            O => \N__46639\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15886\
        );

    \I__8438\ : CascadeMux
    port map (
            O => \N__46636\,
            I => \N__46633\
        );

    \I__8437\ : InMux
    port map (
            O => \N__46633\,
            I => \N__46630\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__46630\,
            I => \N__46627\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__46627\,
            I => \N__46624\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__46624\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_5\
        );

    \I__8433\ : InMux
    port map (
            O => \N__46621\,
            I => \N__46617\
        );

    \I__8432\ : InMux
    port map (
            O => \N__46620\,
            I => \N__46614\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__46617\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__46614\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6\
        );

    \I__8429\ : InMux
    port map (
            O => \N__46609\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15887\
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__46606\,
            I => \N__46603\
        );

    \I__8427\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46600\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__46600\,
            I => \N__46597\
        );

    \I__8425\ : Span4Mux_h
    port map (
            O => \N__46597\,
            I => \N__46594\
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__46594\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_6\
        );

    \I__8423\ : InMux
    port map (
            O => \N__46591\,
            I => \N__46587\
        );

    \I__8422\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46584\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__46587\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__46584\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7\
        );

    \I__8419\ : InMux
    port map (
            O => \N__46579\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15888\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__46576\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19914_cascade_\
        );

    \I__8417\ : InMux
    port map (
            O => \N__46573\,
            I => \N__46569\
        );

    \I__8416\ : InMux
    port map (
            O => \N__46572\,
            I => \N__46566\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__46569\,
            I => \N__46563\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__46566\,
            I => \N__46560\
        );

    \I__8413\ : Odrv4
    port map (
            O => \N__46563\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24\
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__46560\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24\
        );

    \I__8411\ : InMux
    port map (
            O => \N__46555\,
            I => \N__46551\
        );

    \I__8410\ : InMux
    port map (
            O => \N__46554\,
            I => \N__46548\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46545\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__46548\,
            I => \N__46542\
        );

    \I__8407\ : Odrv12
    port map (
            O => \N__46545\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26\
        );

    \I__8406\ : Odrv12
    port map (
            O => \N__46542\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26\
        );

    \I__8405\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46534\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__46534\,
            I => \N__46531\
        );

    \I__8403\ : Odrv4
    port map (
            O => \N__46531\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20102\
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__46528\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20086_cascade_\
        );

    \I__8401\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46522\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__46522\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19890\
        );

    \I__8399\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46515\
        );

    \I__8398\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46512\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46509\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__46512\,
            I => \N__46506\
        );

    \I__8395\ : Span4Mux_v
    port map (
            O => \N__46509\,
            I => \N__46503\
        );

    \I__8394\ : Odrv4
    port map (
            O => \N__46506\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21\
        );

    \I__8393\ : Odrv4
    port map (
            O => \N__46503\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__46498\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20858_cascade_\
        );

    \I__8391\ : InMux
    port map (
            O => \N__46495\,
            I => \N__46492\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__46492\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n452_adj_362\
        );

    \I__8389\ : InMux
    port map (
            O => \N__46489\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17759\
        );

    \I__8388\ : InMux
    port map (
            O => \N__46486\,
            I => \N__46483\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__46483\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n501\
        );

    \I__8386\ : InMux
    port map (
            O => \N__46480\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17760\
        );

    \I__8385\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46474\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__46474\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n550\
        );

    \I__8383\ : InMux
    port map (
            O => \N__46471\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17761\
        );

    \I__8382\ : InMux
    port map (
            O => \N__46468\,
            I => \N__46465\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__46465\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n599\
        );

    \I__8380\ : InMux
    port map (
            O => \N__46462\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17762\
        );

    \I__8379\ : CascadeMux
    port map (
            O => \N__46459\,
            I => \N__46456\
        );

    \I__8378\ : InMux
    port map (
            O => \N__46456\,
            I => \N__46453\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__46453\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n648_adj_347\
        );

    \I__8376\ : InMux
    port map (
            O => \N__46450\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17763\
        );

    \I__8375\ : CascadeMux
    port map (
            O => \N__46447\,
            I => \N__46444\
        );

    \I__8374\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46441\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__46441\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n697\
        );

    \I__8372\ : InMux
    port map (
            O => \N__46438\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17764\
        );

    \I__8371\ : InMux
    port map (
            O => \N__46435\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n747\
        );

    \I__8370\ : InMux
    port map (
            O => \N__46432\,
            I => \N__46429\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__46429\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20108\
        );

    \I__8368\ : CascadeMux
    port map (
            O => \N__46426\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20092_cascade_\
        );

    \I__8367\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46420\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__46420\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n60\
        );

    \I__8365\ : InMux
    port map (
            O => \N__46417\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17751\
        );

    \I__8364\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46411\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__46411\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n109_adj_383\
        );

    \I__8362\ : InMux
    port map (
            O => \N__46408\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17752\
        );

    \I__8361\ : CascadeMux
    port map (
            O => \N__46405\,
            I => \N__46402\
        );

    \I__8360\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46399\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__46399\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n158_adj_375\
        );

    \I__8358\ : InMux
    port map (
            O => \N__46396\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17753\
        );

    \I__8357\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46390\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__46390\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n207\
        );

    \I__8355\ : InMux
    port map (
            O => \N__46387\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17754\
        );

    \I__8354\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46381\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__46381\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n256\
        );

    \I__8352\ : InMux
    port map (
            O => \N__46378\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17755\
        );

    \I__8351\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46372\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__46372\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n305\
        );

    \I__8349\ : InMux
    port map (
            O => \N__46369\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17756\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__46366\,
            I => \N__46363\
        );

    \I__8347\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46360\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__46360\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n354_adj_367\
        );

    \I__8345\ : InMux
    port map (
            O => \N__46357\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17757\
        );

    \I__8344\ : InMux
    port map (
            O => \N__46354\,
            I => \N__46351\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__46351\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n403_adj_365\
        );

    \I__8342\ : InMux
    port map (
            O => \N__46348\,
            I => \bfn_18_19_0_\
        );

    \I__8341\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46342\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__46342\,
            I => \N__46339\
        );

    \I__8339\ : Odrv12
    port map (
            O => \N__46339\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n418_adj_500\
        );

    \I__8338\ : InMux
    port map (
            O => \N__46336\,
            I => \bfn_18_17_0_\
        );

    \I__8337\ : InMux
    port map (
            O => \N__46333\,
            I => \N__46330\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__46330\,
            I => \N__46327\
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__46327\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n467_adj_499\
        );

    \I__8334\ : InMux
    port map (
            O => \N__46324\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17834\
        );

    \I__8333\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46318\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__46318\,
            I => \N__46315\
        );

    \I__8331\ : Odrv4
    port map (
            O => \N__46315\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n516_adj_498\
        );

    \I__8330\ : InMux
    port map (
            O => \N__46312\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17835\
        );

    \I__8329\ : InMux
    port map (
            O => \N__46309\,
            I => \N__46306\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__46306\,
            I => \N__46303\
        );

    \I__8327\ : Odrv12
    port map (
            O => \N__46303\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n565_adj_497\
        );

    \I__8326\ : InMux
    port map (
            O => \N__46300\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17836\
        );

    \I__8325\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46294\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46291\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__46291\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n614_adj_496\
        );

    \I__8322\ : InMux
    port map (
            O => \N__46288\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17837\
        );

    \I__8321\ : InMux
    port map (
            O => \N__46285\,
            I => \N__46282\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__46282\,
            I => \N__46279\
        );

    \I__8319\ : Odrv4
    port map (
            O => \N__46279\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n663_adj_494\
        );

    \I__8318\ : InMux
    port map (
            O => \N__46276\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17838\
        );

    \I__8317\ : CascadeMux
    port map (
            O => \N__46273\,
            I => \N__46270\
        );

    \I__8316\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46267\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__46267\,
            I => \N__46264\
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__46264\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n712_adj_493\
        );

    \I__8313\ : InMux
    port map (
            O => \N__46261\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17839\
        );

    \I__8312\ : InMux
    port map (
            O => \N__46258\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n767\
        );

    \I__8311\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46252\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__46252\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n75\
        );

    \I__8309\ : InMux
    port map (
            O => \N__46249\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17826\
        );

    \I__8308\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46243\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__46243\,
            I => \N__46240\
        );

    \I__8306\ : Odrv4
    port map (
            O => \N__46240\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n124_adj_507\
        );

    \I__8305\ : InMux
    port map (
            O => \N__46237\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17827\
        );

    \I__8304\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46231\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__46231\,
            I => \N__46228\
        );

    \I__8302\ : Odrv12
    port map (
            O => \N__46228\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n173_adj_506\
        );

    \I__8301\ : InMux
    port map (
            O => \N__46225\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17828\
        );

    \I__8300\ : InMux
    port map (
            O => \N__46222\,
            I => \N__46219\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__46219\,
            I => \N__46216\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__46216\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n222_adj_505\
        );

    \I__8297\ : InMux
    port map (
            O => \N__46213\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17829\
        );

    \I__8296\ : InMux
    port map (
            O => \N__46210\,
            I => \N__46207\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__46207\,
            I => \N__46204\
        );

    \I__8294\ : Odrv4
    port map (
            O => \N__46204\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n271_adj_503\
        );

    \I__8293\ : InMux
    port map (
            O => \N__46201\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17830\
        );

    \I__8292\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46195\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__46195\,
            I => \N__46192\
        );

    \I__8290\ : Odrv12
    port map (
            O => \N__46192\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n320_adj_502\
        );

    \I__8289\ : InMux
    port map (
            O => \N__46189\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17831\
        );

    \I__8288\ : CascadeMux
    port map (
            O => \N__46186\,
            I => \N__46183\
        );

    \I__8287\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46180\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__46180\,
            I => \N__46177\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__46177\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n369_adj_501\
        );

    \I__8284\ : InMux
    port map (
            O => \N__46174\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17832\
        );

    \I__8283\ : InMux
    port map (
            O => \N__46171\,
            I => \N__46168\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__46168\,
            I => \N__46165\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__46165\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n372_adj_473\
        );

    \I__8280\ : InMux
    port map (
            O => \N__46162\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17847\
        );

    \I__8279\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46156\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__46156\,
            I => \N__46153\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__46153\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n421_adj_465\
        );

    \I__8276\ : InMux
    port map (
            O => \N__46150\,
            I => \bfn_18_15_0_\
        );

    \I__8275\ : InMux
    port map (
            O => \N__46147\,
            I => \N__46144\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__46144\,
            I => \N__46141\
        );

    \I__8273\ : Odrv4
    port map (
            O => \N__46141\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n470_adj_463\
        );

    \I__8272\ : InMux
    port map (
            O => \N__46138\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17849\
        );

    \I__8271\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46132\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__46132\,
            I => \N__46129\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__46129\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n519_adj_461\
        );

    \I__8268\ : InMux
    port map (
            O => \N__46126\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17850\
        );

    \I__8267\ : InMux
    port map (
            O => \N__46123\,
            I => \N__46120\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__46120\,
            I => \N__46117\
        );

    \I__8265\ : Odrv12
    port map (
            O => \N__46117\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n568_adj_460\
        );

    \I__8264\ : InMux
    port map (
            O => \N__46114\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17851\
        );

    \I__8263\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46108\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__46108\,
            I => \N__46105\
        );

    \I__8261\ : Odrv12
    port map (
            O => \N__46105\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n617_adj_459\
        );

    \I__8260\ : InMux
    port map (
            O => \N__46102\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17852\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__46099\,
            I => \N__46096\
        );

    \I__8258\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46093\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__46093\,
            I => \N__46090\
        );

    \I__8256\ : Span4Mux_v
    port map (
            O => \N__46090\,
            I => \N__46087\
        );

    \I__8255\ : Odrv4
    port map (
            O => \N__46087\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n666\
        );

    \I__8254\ : InMux
    port map (
            O => \N__46084\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17853\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__46081\,
            I => \N__46078\
        );

    \I__8252\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46075\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46072\
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__46072\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n715\
        );

    \I__8249\ : InMux
    port map (
            O => \N__46069\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17854\
        );

    \I__8248\ : InMux
    port map (
            O => \N__46066\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353\
        );

    \I__8247\ : InMux
    port map (
            O => \N__46063\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17880\
        );

    \I__8246\ : InMux
    port map (
            O => \N__46060\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n775\
        );

    \I__8245\ : InMux
    port map (
            O => \N__46057\,
            I => \N__46054\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__46054\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n78_adj_480\
        );

    \I__8243\ : InMux
    port map (
            O => \N__46051\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17841\
        );

    \I__8242\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46045\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__46045\,
            I => \N__46042\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__46042\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n127_adj_479\
        );

    \I__8239\ : InMux
    port map (
            O => \N__46039\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17842\
        );

    \I__8238\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46033\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__46033\,
            I => \N__46030\
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__46030\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n176_adj_478\
        );

    \I__8235\ : InMux
    port map (
            O => \N__46027\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17843\
        );

    \I__8234\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46021\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__46021\,
            I => \N__46018\
        );

    \I__8232\ : Odrv12
    port map (
            O => \N__46018\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n225_adj_477\
        );

    \I__8231\ : InMux
    port map (
            O => \N__46015\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17844\
        );

    \I__8230\ : InMux
    port map (
            O => \N__46012\,
            I => \N__46009\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__46009\,
            I => \N__46006\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__46006\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n274_adj_476\
        );

    \I__8227\ : InMux
    port map (
            O => \N__46003\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17845\
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__46000\,
            I => \N__45997\
        );

    \I__8225\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45994\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__45994\,
            I => \N__45991\
        );

    \I__8223\ : Odrv4
    port map (
            O => \N__45991\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n323_adj_475\
        );

    \I__8222\ : InMux
    port map (
            O => \N__45988\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17846\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__45985\,
            I => \N__45982\
        );

    \I__8220\ : InMux
    port map (
            O => \N__45982\,
            I => \N__45979\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__45979\,
            I => \N__45976\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__45976\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n326_adj_443\
        );

    \I__8217\ : InMux
    port map (
            O => \N__45973\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17872\
        );

    \I__8216\ : InMux
    port map (
            O => \N__45970\,
            I => \N__45967\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__45967\,
            I => \N__45964\
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__45964\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n375_adj_438\
        );

    \I__8213\ : InMux
    port map (
            O => \N__45961\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17873\
        );

    \I__8212\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45955\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__45955\,
            I => \N__45952\
        );

    \I__8210\ : Odrv4
    port map (
            O => \N__45952\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n424_adj_435\
        );

    \I__8209\ : InMux
    port map (
            O => \N__45949\,
            I => \bfn_18_13_0_\
        );

    \I__8208\ : InMux
    port map (
            O => \N__45946\,
            I => \N__45943\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__45943\,
            I => \N__45940\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__45940\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n473_adj_431\
        );

    \I__8205\ : InMux
    port map (
            O => \N__45937\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17875\
        );

    \I__8204\ : InMux
    port map (
            O => \N__45934\,
            I => \N__45931\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__45931\,
            I => \N__45928\
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__45928\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n522_adj_430\
        );

    \I__8201\ : InMux
    port map (
            O => \N__45925\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17876\
        );

    \I__8200\ : InMux
    port map (
            O => \N__45922\,
            I => \N__45919\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__45919\,
            I => \N__45916\
        );

    \I__8198\ : Odrv12
    port map (
            O => \N__45916\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n571\
        );

    \I__8197\ : InMux
    port map (
            O => \N__45913\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17877\
        );

    \I__8196\ : InMux
    port map (
            O => \N__45910\,
            I => \N__45907\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__45907\,
            I => \N__45904\
        );

    \I__8194\ : Odrv4
    port map (
            O => \N__45904\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n620\
        );

    \I__8193\ : InMux
    port map (
            O => \N__45901\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17878\
        );

    \I__8192\ : CascadeMux
    port map (
            O => \N__45898\,
            I => \N__45895\
        );

    \I__8191\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45892\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__45892\,
            I => \N__45889\
        );

    \I__8189\ : Span4Mux_v
    port map (
            O => \N__45889\,
            I => \N__45886\
        );

    \I__8188\ : Odrv4
    port map (
            O => \N__45886\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n669\
        );

    \I__8187\ : InMux
    port map (
            O => \N__45883\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17879\
        );

    \I__8186\ : InMux
    port map (
            O => \N__45880\,
            I => \N__45877\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__45877\,
            I => \N__45874\
        );

    \I__8184\ : Odrv12
    port map (
            O => \N__45874\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n718\
        );

    \I__8183\ : InMux
    port map (
            O => \N__45871\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17894\
        );

    \I__8182\ : InMux
    port map (
            O => \N__45868\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17895\
        );

    \I__8181\ : InMux
    port map (
            O => \N__45865\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n779\
        );

    \I__8180\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45859\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__45859\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n81_adj_457\
        );

    \I__8178\ : InMux
    port map (
            O => \N__45856\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17867\
        );

    \I__8177\ : InMux
    port map (
            O => \N__45853\,
            I => \N__45850\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__45850\,
            I => \N__45847\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__45847\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n130_adj_453\
        );

    \I__8174\ : InMux
    port map (
            O => \N__45844\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17868\
        );

    \I__8173\ : InMux
    port map (
            O => \N__45841\,
            I => \N__45838\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__45838\,
            I => \N__45835\
        );

    \I__8171\ : Odrv12
    port map (
            O => \N__45835\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n179_adj_452\
        );

    \I__8170\ : InMux
    port map (
            O => \N__45832\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17869\
        );

    \I__8169\ : InMux
    port map (
            O => \N__45829\,
            I => \N__45826\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__45826\,
            I => \N__45823\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__45823\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n228_adj_450\
        );

    \I__8166\ : InMux
    port map (
            O => \N__45820\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17870\
        );

    \I__8165\ : InMux
    port map (
            O => \N__45817\,
            I => \N__45814\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__45814\,
            I => \N__45811\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__45811\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n277_adj_448\
        );

    \I__8162\ : InMux
    port map (
            O => \N__45808\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17871\
        );

    \I__8161\ : InMux
    port map (
            O => \N__45805\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17885\
        );

    \I__8160\ : InMux
    port map (
            O => \N__45802\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17886\
        );

    \I__8159\ : InMux
    port map (
            O => \N__45799\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17887\
        );

    \I__8158\ : InMux
    port map (
            O => \N__45796\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17888\
        );

    \I__8157\ : InMux
    port map (
            O => \N__45793\,
            I => \bfn_18_11_0_\
        );

    \I__8156\ : InMux
    port map (
            O => \N__45790\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17890\
        );

    \I__8155\ : InMux
    port map (
            O => \N__45787\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17891\
        );

    \I__8154\ : InMux
    port map (
            O => \N__45784\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17892\
        );

    \I__8153\ : InMux
    port map (
            O => \N__45781\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17893\
        );

    \I__8152\ : InMux
    port map (
            O => \N__45778\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17952\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__45775\,
            I => \N__45771\
        );

    \I__8150\ : InMux
    port map (
            O => \N__45774\,
            I => \N__45768\
        );

    \I__8149\ : InMux
    port map (
            O => \N__45771\,
            I => \N__45765\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__45768\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n785\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__45765\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n785\
        );

    \I__8146\ : InMux
    port map (
            O => \N__45760\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17953\
        );

    \I__8145\ : CascadeMux
    port map (
            O => \N__45757\,
            I => \N__45752\
        );

    \I__8144\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45749\
        );

    \I__8143\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45746\
        );

    \I__8142\ : InMux
    port map (
            O => \N__45752\,
            I => \N__45743\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__45749\,
            I => \N__45738\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__45746\,
            I => \N__45738\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__45743\,
            I => \N__45735\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__45738\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n789\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__45735\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n789\
        );

    \I__8136\ : InMux
    port map (
            O => \N__45730\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17954\
        );

    \I__8135\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45724\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__45724\,
            I => n793
        );

    \I__8133\ : InMux
    port map (
            O => \N__45721\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17955\
        );

    \I__8132\ : InMux
    port map (
            O => \N__45718\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n795\
        );

    \I__8131\ : CascadeMux
    port map (
            O => \N__45715\,
            I => \N__45712\
        );

    \I__8130\ : InMux
    port map (
            O => \N__45712\,
            I => \N__45709\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__45709\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n84_adj_389\
        );

    \I__8128\ : InMux
    port map (
            O => \N__45706\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17882\
        );

    \I__8127\ : InMux
    port map (
            O => \N__45703\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17883\
        );

    \I__8126\ : InMux
    port map (
            O => \N__45700\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17884\
        );

    \I__8125\ : InMux
    port map (
            O => \N__45697\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17944\
        );

    \I__8124\ : InMux
    port map (
            O => \N__45694\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17945\
        );

    \I__8123\ : InMux
    port map (
            O => \N__45691\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17946\
        );

    \I__8122\ : InMux
    port map (
            O => \N__45688\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17947\
        );

    \I__8121\ : InMux
    port map (
            O => \N__45685\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17948\
        );

    \I__8120\ : InMux
    port map (
            O => \N__45682\,
            I => \bfn_18_9_0_\
        );

    \I__8119\ : InMux
    port map (
            O => \N__45679\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17950\
        );

    \I__8118\ : InMux
    port map (
            O => \N__45676\,
            I => \N__45673\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__45673\,
            I => \N__45669\
        );

    \I__8116\ : InMux
    port map (
            O => \N__45672\,
            I => \N__45666\
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__45669\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n777\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__45666\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n777\
        );

    \I__8113\ : InMux
    port map (
            O => \N__45661\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17951\
        );

    \I__8112\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45655\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__45655\,
            I => \N__45651\
        );

    \I__8110\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45648\
        );

    \I__8109\ : Odrv4
    port map (
            O => \N__45651\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n781\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__45648\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n781\
        );

    \I__8107\ : InMux
    port map (
            O => \N__45643\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17274\
        );

    \I__8106\ : CascadeMux
    port map (
            O => \N__45640\,
            I => \N__45636\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__45639\,
            I => \N__45633\
        );

    \I__8104\ : InMux
    port map (
            O => \N__45636\,
            I => \N__45629\
        );

    \I__8103\ : InMux
    port map (
            O => \N__45633\,
            I => \N__45624\
        );

    \I__8102\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45624\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__45629\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n427\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__45624\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n427\
        );

    \I__8099\ : InMux
    port map (
            O => \N__45619\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17275\
        );

    \I__8098\ : InMux
    port map (
            O => \N__45616\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352\
        );

    \I__8097\ : InMux
    port map (
            O => \N__45613\,
            I => \N__45610\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45606\
        );

    \I__8095\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45603\
        );

    \I__8094\ : Span4Mux_v
    port map (
            O => \N__45606\,
            I => \N__45598\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__45603\,
            I => \N__45598\
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__45598\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_23\
        );

    \I__8091\ : InMux
    port map (
            O => \N__45595\,
            I => \N__45589\
        );

    \I__8090\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45589\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__45589\,
            I => \N__45586\
        );

    \I__8088\ : Odrv12
    port map (
            O => \N__45586\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_19\
        );

    \I__8087\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45579\
        );

    \I__8086\ : InMux
    port map (
            O => \N__45582\,
            I => \N__45576\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__45579\,
            I => \N__45571\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__45576\,
            I => \N__45571\
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__45571\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_22\
        );

    \I__8082\ : InMux
    port map (
            O => \N__45568\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17942\
        );

    \I__8081\ : InMux
    port map (
            O => \N__45565\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17943\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__45562\,
            I => \N__45559\
        );

    \I__8079\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45556\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__45556\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n84\
        );

    \I__8077\ : InMux
    port map (
            O => \N__45553\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17266\
        );

    \I__8076\ : InMux
    port map (
            O => \N__45550\,
            I => \N__45547\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__45547\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n133\
        );

    \I__8074\ : InMux
    port map (
            O => \N__45544\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17267\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__45541\,
            I => \N__45538\
        );

    \I__8072\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45535\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__45535\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n182\
        );

    \I__8070\ : InMux
    port map (
            O => \N__45532\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17268\
        );

    \I__8069\ : InMux
    port map (
            O => \N__45529\,
            I => \N__45526\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__45526\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n231\
        );

    \I__8067\ : InMux
    port map (
            O => \N__45523\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17269\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__45520\,
            I => \N__45517\
        );

    \I__8065\ : InMux
    port map (
            O => \N__45517\,
            I => \N__45514\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__45514\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n280\
        );

    \I__8063\ : InMux
    port map (
            O => \N__45511\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17270\
        );

    \I__8062\ : InMux
    port map (
            O => \N__45508\,
            I => \N__45505\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__45505\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n329\
        );

    \I__8060\ : InMux
    port map (
            O => \N__45502\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17271\
        );

    \I__8059\ : CascadeMux
    port map (
            O => \N__45499\,
            I => \N__45496\
        );

    \I__8058\ : InMux
    port map (
            O => \N__45496\,
            I => \N__45493\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__45493\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n378\
        );

    \I__8056\ : InMux
    port map (
            O => \N__45490\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17272\
        );

    \I__8055\ : InMux
    port map (
            O => \N__45487\,
            I => \bfn_18_6_0_\
        );

    \I__8054\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45481\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__45481\,
            I => \N__45478\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__45478\,
            I => \N__45474\
        );

    \I__8051\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45471\
        );

    \I__8050\ : Span4Mux_h
    port map (
            O => \N__45474\,
            I => \N__45468\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45465\
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__45468\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n769\
        );

    \I__8047\ : Odrv4
    port map (
            O => \N__45465\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n769\
        );

    \I__8046\ : InMux
    port map (
            O => \N__45460\,
            I => \bfn_17_26_0_\
        );

    \I__8045\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45453\
        );

    \I__8044\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45450\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__45453\,
            I => \N__45447\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__45450\,
            I => \N__45444\
        );

    \I__8041\ : Span4Mux_v
    port map (
            O => \N__45447\,
            I => \N__45441\
        );

    \I__8040\ : Span4Mux_v
    port map (
            O => \N__45444\,
            I => \N__45438\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__45441\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n773\
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__45438\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n773\
        );

    \I__8037\ : InMux
    port map (
            O => \N__45433\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18377\
        );

    \I__8036\ : InMux
    port map (
            O => \N__45430\,
            I => \N__45427\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__45427\,
            I => \N__45423\
        );

    \I__8034\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45420\
        );

    \I__8033\ : Span4Mux_h
    port map (
            O => \N__45423\,
            I => \N__45417\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__45420\,
            I => \N__45414\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__45417\,
            I => \N__45409\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__45414\,
            I => \N__45409\
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__45409\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n777\
        );

    \I__8028\ : InMux
    port map (
            O => \N__45406\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18378\
        );

    \I__8027\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__45400\,
            I => \N__45396\
        );

    \I__8025\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45393\
        );

    \I__8024\ : Span4Mux_v
    port map (
            O => \N__45396\,
            I => \N__45390\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__45393\,
            I => \N__45387\
        );

    \I__8022\ : Odrv4
    port map (
            O => \N__45390\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n781\
        );

    \I__8021\ : Odrv12
    port map (
            O => \N__45387\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n781\
        );

    \I__8020\ : InMux
    port map (
            O => \N__45382\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18379\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__45379\,
            I => \N__45376\
        );

    \I__8018\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45372\
        );

    \I__8017\ : InMux
    port map (
            O => \N__45375\,
            I => \N__45369\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__45372\,
            I => \N__45366\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__45369\,
            I => \N__45363\
        );

    \I__8014\ : Odrv12
    port map (
            O => \N__45366\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n785\
        );

    \I__8013\ : Odrv4
    port map (
            O => \N__45363\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n785\
        );

    \I__8012\ : InMux
    port map (
            O => \N__45358\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18380\
        );

    \I__8011\ : CascadeMux
    port map (
            O => \N__45355\,
            I => \N__45352\
        );

    \I__8010\ : InMux
    port map (
            O => \N__45352\,
            I => \N__45349\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__45349\,
            I => \N__45346\
        );

    \I__8008\ : Odrv12
    port map (
            O => \N__45346\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n789\
        );

    \I__8007\ : InMux
    port map (
            O => \N__45343\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18381\
        );

    \I__8006\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45337\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45334\
        );

    \I__8004\ : Odrv12
    port map (
            O => \N__45334\,
            I => n793_adj_2424
        );

    \I__8003\ : InMux
    port map (
            O => \N__45331\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18382\
        );

    \I__8002\ : InMux
    port map (
            O => \N__45328\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n795\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__45325\,
            I => \N__45322\
        );

    \I__8000\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45318\
        );

    \I__7999\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45315\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__45318\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n737\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__45315\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n737\
        );

    \I__7996\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45307\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__45307\,
            I => \N__45304\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__45304\,
            I => \N__45300\
        );

    \I__7993\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45297\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__45300\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n741\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__45297\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n741\
        );

    \I__7990\ : InMux
    port map (
            O => \N__45292\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18369\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__45289\,
            I => \N__45286\
        );

    \I__7988\ : InMux
    port map (
            O => \N__45286\,
            I => \N__45283\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__45283\,
            I => \N__45279\
        );

    \I__7986\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45276\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__45279\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n745\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__45276\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n745\
        );

    \I__7983\ : InMux
    port map (
            O => \N__45271\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18370\
        );

    \I__7982\ : InMux
    port map (
            O => \N__45268\,
            I => \N__45265\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__45265\,
            I => \N__45262\
        );

    \I__7980\ : Span4Mux_v
    port map (
            O => \N__45262\,
            I => \N__45259\
        );

    \I__7979\ : Sp12to4
    port map (
            O => \N__45259\,
            I => \N__45255\
        );

    \I__7978\ : InMux
    port map (
            O => \N__45258\,
            I => \N__45252\
        );

    \I__7977\ : Span12Mux_h
    port map (
            O => \N__45255\,
            I => \N__45247\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__45252\,
            I => \N__45247\
        );

    \I__7975\ : Odrv12
    port map (
            O => \N__45247\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n749\
        );

    \I__7974\ : InMux
    port map (
            O => \N__45244\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18371\
        );

    \I__7973\ : InMux
    port map (
            O => \N__45241\,
            I => \N__45238\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__45238\,
            I => \N__45234\
        );

    \I__7971\ : InMux
    port map (
            O => \N__45237\,
            I => \N__45231\
        );

    \I__7970\ : Span4Mux_v
    port map (
            O => \N__45234\,
            I => \N__45228\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__45231\,
            I => \N__45225\
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__45228\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n753\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__45225\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n753\
        );

    \I__7966\ : InMux
    port map (
            O => \N__45220\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18372\
        );

    \I__7965\ : InMux
    port map (
            O => \N__45217\,
            I => \N__45214\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__45214\,
            I => \N__45210\
        );

    \I__7963\ : InMux
    port map (
            O => \N__45213\,
            I => \N__45207\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__45210\,
            I => \N__45204\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__45207\,
            I => \N__45201\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__45204\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n757\
        );

    \I__7959\ : Odrv12
    port map (
            O => \N__45201\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n757\
        );

    \I__7958\ : InMux
    port map (
            O => \N__45196\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18373\
        );

    \I__7957\ : InMux
    port map (
            O => \N__45193\,
            I => \N__45190\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__45190\,
            I => \N__45186\
        );

    \I__7955\ : InMux
    port map (
            O => \N__45189\,
            I => \N__45183\
        );

    \I__7954\ : Span4Mux_v
    port map (
            O => \N__45186\,
            I => \N__45180\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__45183\,
            I => \N__45177\
        );

    \I__7952\ : Odrv4
    port map (
            O => \N__45180\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n761\
        );

    \I__7951\ : Odrv4
    port map (
            O => \N__45177\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n761\
        );

    \I__7950\ : InMux
    port map (
            O => \N__45172\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18374\
        );

    \I__7949\ : InMux
    port map (
            O => \N__45169\,
            I => \N__45166\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__45166\,
            I => \N__45163\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__45163\,
            I => \N__45159\
        );

    \I__7946\ : InMux
    port map (
            O => \N__45162\,
            I => \N__45156\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__45159\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n765\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__45156\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n765\
        );

    \I__7943\ : InMux
    port map (
            O => \N__45151\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18375\
        );

    \I__7942\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45142\
        );

    \I__7941\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45142\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__45142\,
            I => \N__45139\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__45139\,
            I => \N__45136\
        );

    \I__7938\ : Odrv4
    port map (
            O => \N__45136\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_20\
        );

    \I__7937\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45130\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__45130\,
            I => \N__45116\
        );

    \I__7935\ : InMux
    port map (
            O => \N__45129\,
            I => \N__45113\
        );

    \I__7934\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45108\
        );

    \I__7933\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45108\
        );

    \I__7932\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45101\
        );

    \I__7931\ : InMux
    port map (
            O => \N__45125\,
            I => \N__45101\
        );

    \I__7930\ : InMux
    port map (
            O => \N__45124\,
            I => \N__45101\
        );

    \I__7929\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45094\
        );

    \I__7928\ : InMux
    port map (
            O => \N__45122\,
            I => \N__45094\
        );

    \I__7927\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45094\
        );

    \I__7926\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45089\
        );

    \I__7925\ : InMux
    port map (
            O => \N__45119\,
            I => \N__45089\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__45116\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__45113\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__45108\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__45101\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__45094\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__45089\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\
        );

    \I__7918\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45073\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__45073\,
            I => \N__45069\
        );

    \I__7916\ : InMux
    port map (
            O => \N__45072\,
            I => \N__45066\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__45069\,
            I => \N__45063\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__45066\,
            I => \N__45060\
        );

    \I__7913\ : Odrv4
    port map (
            O => \N__45063\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18\
        );

    \I__7912\ : Odrv4
    port map (
            O => \N__45060\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18\
        );

    \I__7911\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45052\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45044\
        );

    \I__7909\ : InMux
    port map (
            O => \N__45051\,
            I => \N__45041\
        );

    \I__7908\ : InMux
    port map (
            O => \N__45050\,
            I => \N__45036\
        );

    \I__7907\ : InMux
    port map (
            O => \N__45049\,
            I => \N__45036\
        );

    \I__7906\ : InMux
    port map (
            O => \N__45048\,
            I => \N__45031\
        );

    \I__7905\ : InMux
    port map (
            O => \N__45047\,
            I => \N__45031\
        );

    \I__7904\ : Odrv4
    port map (
            O => \N__45044\,
            I => \Error_sub_temp_30_adj_2385\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__45041\,
            I => \Error_sub_temp_30_adj_2385\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__45036\,
            I => \Error_sub_temp_30_adj_2385\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__45031\,
            I => \Error_sub_temp_30_adj_2385\
        );

    \I__7900\ : InMux
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__45019\,
            I => \N__45015\
        );

    \I__7898\ : InMux
    port map (
            O => \N__45018\,
            I => \N__45012\
        );

    \I__7897\ : Span4Mux_v
    port map (
            O => \N__45015\,
            I => \N__45007\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__45012\,
            I => \N__45007\
        );

    \I__7895\ : Odrv4
    port map (
            O => \N__45007\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_16\
        );

    \I__7894\ : InMux
    port map (
            O => \N__45004\,
            I => \N__45001\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44998\
        );

    \I__7892\ : Span4Mux_v
    port map (
            O => \N__44998\,
            I => \N__44994\
        );

    \I__7891\ : InMux
    port map (
            O => \N__44997\,
            I => \N__44991\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__44994\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__44991\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__44986\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19450_cascade_\
        );

    \I__7887\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44980\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__44980\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19743\
        );

    \I__7885\ : CascadeMux
    port map (
            O => \N__44977\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19741_cascade_\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__44974\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20180_cascade_\
        );

    \I__7883\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44968\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__44968\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n22\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__44965\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19827_cascade_\
        );

    \I__7880\ : InMux
    port map (
            O => \N__44962\,
            I => \N__44959\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__44959\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19812\
        );

    \I__7878\ : CascadeMux
    port map (
            O => \N__44956\,
            I => \N__44943\
        );

    \I__7877\ : InMux
    port map (
            O => \N__44955\,
            I => \N__44937\
        );

    \I__7876\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44937\
        );

    \I__7875\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44934\
        );

    \I__7874\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44925\
        );

    \I__7873\ : InMux
    port map (
            O => \N__44951\,
            I => \N__44925\
        );

    \I__7872\ : InMux
    port map (
            O => \N__44950\,
            I => \N__44925\
        );

    \I__7871\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44925\
        );

    \I__7870\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44918\
        );

    \I__7869\ : InMux
    port map (
            O => \N__44947\,
            I => \N__44918\
        );

    \I__7868\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44918\
        );

    \I__7867\ : InMux
    port map (
            O => \N__44943\,
            I => \N__44913\
        );

    \I__7866\ : InMux
    port map (
            O => \N__44942\,
            I => \N__44913\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44908\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__44934\,
            I => \N__44901\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__44925\,
            I => \N__44901\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__44918\,
            I => \N__44901\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__44913\,
            I => \N__44898\
        );

    \I__7860\ : InMux
    port map (
            O => \N__44912\,
            I => \N__44895\
        );

    \I__7859\ : InMux
    port map (
            O => \N__44911\,
            I => \N__44890\
        );

    \I__7858\ : Span4Mux_v
    port map (
            O => \N__44908\,
            I => \N__44885\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__44901\,
            I => \N__44885\
        );

    \I__7856\ : Span4Mux_v
    port map (
            O => \N__44898\,
            I => \N__44880\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44880\
        );

    \I__7854\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44877\
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__44893\,
            I => \N__44874\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__44890\,
            I => \N__44871\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__44885\,
            I => \N__44864\
        );

    \I__7850\ : Span4Mux_h
    port map (
            O => \N__44880\,
            I => \N__44864\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__44877\,
            I => \N__44864\
        );

    \I__7848\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44861\
        );

    \I__7847\ : Span4Mux_v
    port map (
            O => \N__44871\,
            I => \N__44857\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__44864\,
            I => \N__44852\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__44861\,
            I => \N__44852\
        );

    \I__7844\ : CascadeMux
    port map (
            O => \N__44860\,
            I => \N__44849\
        );

    \I__7843\ : Span4Mux_h
    port map (
            O => \N__44857\,
            I => \N__44846\
        );

    \I__7842\ : Span4Mux_v
    port map (
            O => \N__44852\,
            I => \N__44843\
        );

    \I__7841\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44840\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__44846\,
            I => \Amp25_out1_14\
        );

    \I__7839\ : Odrv4
    port map (
            O => \N__44843\,
            I => \Amp25_out1_14\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__44840\,
            I => \Amp25_out1_14\
        );

    \I__7837\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44829\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__44832\,
            I => \N__44824\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__44829\,
            I => \N__44818\
        );

    \I__7834\ : InMux
    port map (
            O => \N__44828\,
            I => \N__44815\
        );

    \I__7833\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44808\
        );

    \I__7832\ : InMux
    port map (
            O => \N__44824\,
            I => \N__44808\
        );

    \I__7831\ : InMux
    port map (
            O => \N__44823\,
            I => \N__44808\
        );

    \I__7830\ : InMux
    port map (
            O => \N__44822\,
            I => \N__44802\
        );

    \I__7829\ : InMux
    port map (
            O => \N__44821\,
            I => \N__44802\
        );

    \I__7828\ : Span4Mux_v
    port map (
            O => \N__44818\,
            I => \N__44795\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__44815\,
            I => \N__44795\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__44808\,
            I => \N__44795\
        );

    \I__7825\ : InMux
    port map (
            O => \N__44807\,
            I => \N__44792\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__44802\,
            I => n142_adj_2422
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__44795\,
            I => n142_adj_2422
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__44792\,
            I => n142_adj_2422
        );

    \I__7821\ : InMux
    port map (
            O => \N__44785\,
            I => \N__44782\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__44782\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n6_adj_763\
        );

    \I__7819\ : InMux
    port map (
            O => \N__44779\,
            I => \N__44776\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__44776\,
            I => \N__44773\
        );

    \I__7817\ : Odrv12
    port map (
            O => \N__44773\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n139_adj_727\
        );

    \I__7816\ : CascadeMux
    port map (
            O => \N__44770\,
            I => \n141_adj_2421_cascade_\
        );

    \I__7815\ : InMux
    port map (
            O => \N__44767\,
            I => \N__44759\
        );

    \I__7814\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44759\
        );

    \I__7813\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44754\
        );

    \I__7812\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44754\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__44759\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__44754\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761\
        );

    \I__7809\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44745\
        );

    \I__7808\ : InMux
    port map (
            O => \N__44748\,
            I => \N__44742\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__44745\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__44742\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19\
        );

    \I__7805\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44734\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__44734\,
            I => \N__44731\
        );

    \I__7803\ : Odrv12
    port map (
            O => \N__44731\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n602\
        );

    \I__7802\ : InMux
    port map (
            O => \N__44728\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17777\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__44725\,
            I => \N__44722\
        );

    \I__7800\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44719\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__44719\,
            I => \N__44716\
        );

    \I__7798\ : Odrv4
    port map (
            O => \N__44716\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n651_adj_474\
        );

    \I__7797\ : InMux
    port map (
            O => \N__44713\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17778\
        );

    \I__7796\ : CascadeMux
    port map (
            O => \N__44710\,
            I => \N__44707\
        );

    \I__7795\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44704\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__44704\,
            I => \N__44701\
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__44701\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n700_adj_455\
        );

    \I__7792\ : InMux
    port map (
            O => \N__44698\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17779\
        );

    \I__7791\ : InMux
    port map (
            O => \N__44695\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n751\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__44692\,
            I => \n142_adj_2422_cascade_\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__44689\,
            I => \N__44684\
        );

    \I__7788\ : InMux
    port map (
            O => \N__44688\,
            I => \N__44677\
        );

    \I__7787\ : InMux
    port map (
            O => \N__44687\,
            I => \N__44677\
        );

    \I__7786\ : InMux
    port map (
            O => \N__44684\,
            I => \N__44677\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__44677\,
            I => \N__44674\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__44674\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755\
        );

    \I__7783\ : CascadeMux
    port map (
            O => \N__44671\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755_cascade_\
        );

    \I__7782\ : InMux
    port map (
            O => \N__44668\,
            I => \N__44662\
        );

    \I__7781\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44662\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__44662\,
            I => \N__44659\
        );

    \I__7779\ : Odrv4
    port map (
            O => \N__44659\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n14_adj_756\
        );

    \I__7778\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44653\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__44653\,
            I => \N__44650\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__44650\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n161\
        );

    \I__7775\ : InMux
    port map (
            O => \N__44647\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17768\
        );

    \I__7774\ : InMux
    port map (
            O => \N__44644\,
            I => \N__44641\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__44641\,
            I => \N__44638\
        );

    \I__7772\ : Odrv12
    port map (
            O => \N__44638\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n210\
        );

    \I__7771\ : InMux
    port map (
            O => \N__44635\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17769\
        );

    \I__7770\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44629\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__44629\,
            I => \N__44626\
        );

    \I__7768\ : Odrv4
    port map (
            O => \N__44626\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n259\
        );

    \I__7767\ : InMux
    port map (
            O => \N__44623\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17770\
        );

    \I__7766\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44617\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__44617\,
            I => \N__44614\
        );

    \I__7764\ : Odrv4
    port map (
            O => \N__44614\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n308_adj_368\
        );

    \I__7763\ : InMux
    port map (
            O => \N__44611\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17771\
        );

    \I__7762\ : CascadeMux
    port map (
            O => \N__44608\,
            I => \N__44605\
        );

    \I__7761\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44602\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__44602\,
            I => \N__44599\
        );

    \I__7759\ : Odrv4
    port map (
            O => \N__44599\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n357_adj_366\
        );

    \I__7758\ : InMux
    port map (
            O => \N__44596\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17772\
        );

    \I__7757\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44590\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__44590\,
            I => \N__44587\
        );

    \I__7755\ : Odrv12
    port map (
            O => \N__44587\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n406_adj_363\
        );

    \I__7754\ : InMux
    port map (
            O => \N__44584\,
            I => \bfn_17_19_0_\
        );

    \I__7753\ : InMux
    port map (
            O => \N__44581\,
            I => \N__44578\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__44578\,
            I => \N__44575\
        );

    \I__7751\ : Odrv12
    port map (
            O => \N__44575\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n455_adj_350\
        );

    \I__7750\ : InMux
    port map (
            O => \N__44572\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17774\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__44569\,
            I => \N__44566\
        );

    \I__7748\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44563\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__44563\,
            I => \N__44560\
        );

    \I__7746\ : Odrv12
    port map (
            O => \N__44560\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n504\
        );

    \I__7745\ : InMux
    port map (
            O => \N__44557\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17775\
        );

    \I__7744\ : InMux
    port map (
            O => \N__44554\,
            I => \N__44551\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__44551\,
            I => \N__44548\
        );

    \I__7742\ : Odrv4
    port map (
            O => \N__44548\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n553\
        );

    \I__7741\ : InMux
    port map (
            O => \N__44545\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17776\
        );

    \I__7740\ : InMux
    port map (
            O => \N__44542\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17790\
        );

    \I__7739\ : InMux
    port map (
            O => \N__44539\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17791\
        );

    \I__7738\ : InMux
    port map (
            O => \N__44536\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17792\
        );

    \I__7737\ : InMux
    port map (
            O => \N__44533\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17793\
        );

    \I__7736\ : InMux
    port map (
            O => \N__44530\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17794\
        );

    \I__7735\ : InMux
    port map (
            O => \N__44527\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n755\
        );

    \I__7734\ : InMux
    port map (
            O => \N__44524\,
            I => \N__44521\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__44521\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n63_adj_384\
        );

    \I__7732\ : InMux
    port map (
            O => \N__44518\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17766\
        );

    \I__7731\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44512\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44509\
        );

    \I__7729\ : Odrv12
    port map (
            O => \N__44509\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n112\
        );

    \I__7728\ : InMux
    port map (
            O => \N__44506\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17767\
        );

    \I__7727\ : InMux
    port map (
            O => \N__44503\,
            I => \N__44500\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__44500\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n66_adj_433\
        );

    \I__7725\ : InMux
    port map (
            O => \N__44497\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17781\
        );

    \I__7724\ : InMux
    port map (
            O => \N__44494\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17782\
        );

    \I__7723\ : InMux
    port map (
            O => \N__44491\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17783\
        );

    \I__7722\ : InMux
    port map (
            O => \N__44488\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17784\
        );

    \I__7721\ : InMux
    port map (
            O => \N__44485\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17785\
        );

    \I__7720\ : InMux
    port map (
            O => \N__44482\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17786\
        );

    \I__7719\ : InMux
    port map (
            O => \N__44479\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17787\
        );

    \I__7718\ : InMux
    port map (
            O => \N__44476\,
            I => \bfn_17_16_0_\
        );

    \I__7717\ : InMux
    port map (
            O => \N__44473\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17789\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__44470\,
            I => \foc.u_Park_Transform.n7_cascade_\
        );

    \I__7715\ : InMux
    port map (
            O => \N__44467\,
            I => \N__44464\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__44464\,
            I => \N__44460\
        );

    \I__7713\ : InMux
    port map (
            O => \N__44463\,
            I => \N__44457\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__44460\,
            I => \N__44454\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__44457\,
            I => \N__44451\
        );

    \I__7710\ : Span4Mux_h
    port map (
            O => \N__44454\,
            I => \N__44448\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__44451\,
            I => \N__44445\
        );

    \I__7708\ : Odrv4
    port map (
            O => \N__44448\,
            I => \foc.u_Park_Transform.n791\
        );

    \I__7707\ : Odrv4
    port map (
            O => \N__44445\,
            I => \foc.u_Park_Transform.n791\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__44440\,
            I => \foc.u_Park_Transform.n4_cascade_\
        );

    \I__7705\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44431\
        );

    \I__7704\ : InMux
    port map (
            O => \N__44436\,
            I => \N__44428\
        );

    \I__7703\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44423\
        );

    \I__7702\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44423\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__44431\,
            I => \N__44419\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__44428\,
            I => \N__44414\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__44423\,
            I => \N__44414\
        );

    \I__7698\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44411\
        );

    \I__7697\ : Span4Mux_v
    port map (
            O => \N__44419\,
            I => \N__44406\
        );

    \I__7696\ : Span12Mux_v
    port map (
            O => \N__44414\,
            I => \N__44401\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__44411\,
            I => \N__44401\
        );

    \I__7694\ : InMux
    port map (
            O => \N__44410\,
            I => \N__44396\
        );

    \I__7693\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44396\
        );

    \I__7692\ : Sp12to4
    port map (
            O => \N__44406\,
            I => \N__44387\
        );

    \I__7691\ : Span12Mux_h
    port map (
            O => \N__44401\,
            I => \N__44387\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__44396\,
            I => \N__44384\
        );

    \I__7689\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44375\
        );

    \I__7688\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44375\
        );

    \I__7687\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44375\
        );

    \I__7686\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44375\
        );

    \I__7685\ : Odrv12
    port map (
            O => \N__44387\,
            I => \Look_Up_Table_out1_1_13\
        );

    \I__7684\ : Odrv4
    port map (
            O => \N__44384\,
            I => \Look_Up_Table_out1_1_13\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__44375\,
            I => \Look_Up_Table_out1_1_13\
        );

    \I__7682\ : InMux
    port map (
            O => \N__44368\,
            I => \N__44365\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__44365\,
            I => \N__44361\
        );

    \I__7680\ : InMux
    port map (
            O => \N__44364\,
            I => \N__44358\
        );

    \I__7679\ : Odrv4
    port map (
            O => \N__44361\,
            I => \foc.u_Park_Transform.n14\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__44358\,
            I => \foc.u_Park_Transform.n14\
        );

    \I__7677\ : CascadeMux
    port map (
            O => \N__44353\,
            I => \n628_cascade_\
        );

    \I__7676\ : CascadeMux
    port map (
            O => \N__44350\,
            I => \N__44346\
        );

    \I__7675\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44341\
        );

    \I__7674\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44341\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__44341\,
            I => \N__44336\
        );

    \I__7672\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44333\
        );

    \I__7671\ : InMux
    port map (
            O => \N__44339\,
            I => \N__44330\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__44336\,
            I => \foc.u_Park_Transform.n12\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__44333\,
            I => \foc.u_Park_Transform.n12\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__44330\,
            I => \foc.u_Park_Transform.n12\
        );

    \I__7667\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44320\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__44320\,
            I => \N__44310\
        );

    \I__7665\ : InMux
    port map (
            O => \N__44319\,
            I => \N__44305\
        );

    \I__7664\ : InMux
    port map (
            O => \N__44318\,
            I => \N__44305\
        );

    \I__7663\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44298\
        );

    \I__7662\ : InMux
    port map (
            O => \N__44316\,
            I => \N__44298\
        );

    \I__7661\ : InMux
    port map (
            O => \N__44315\,
            I => \N__44298\
        );

    \I__7660\ : InMux
    port map (
            O => \N__44314\,
            I => \N__44293\
        );

    \I__7659\ : InMux
    port map (
            O => \N__44313\,
            I => \N__44293\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__44310\,
            I => \N__44288\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__44305\,
            I => \N__44285\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__44298\,
            I => \N__44282\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44279\
        );

    \I__7654\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44274\
        );

    \I__7653\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44274\
        );

    \I__7652\ : Span4Mux_v
    port map (
            O => \N__44288\,
            I => \N__44271\
        );

    \I__7651\ : Span4Mux_h
    port map (
            O => \N__44285\,
            I => \N__44268\
        );

    \I__7650\ : Span4Mux_h
    port map (
            O => \N__44282\,
            I => \N__44261\
        );

    \I__7649\ : Span4Mux_h
    port map (
            O => \N__44279\,
            I => \N__44261\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__44274\,
            I => \N__44261\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__44271\,
            I => n142
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__44268\,
            I => n142
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__44261\,
            I => n142
        );

    \I__7644\ : InMux
    port map (
            O => \N__44254\,
            I => \N__44250\
        );

    \I__7643\ : InMux
    port map (
            O => \N__44253\,
            I => \N__44247\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__44250\,
            I => \N__44242\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__44247\,
            I => \N__44242\
        );

    \I__7640\ : Span4Mux_v
    port map (
            O => \N__44242\,
            I => \N__44236\
        );

    \I__7639\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44233\
        );

    \I__7638\ : InMux
    port map (
            O => \N__44240\,
            I => \N__44230\
        );

    \I__7637\ : InMux
    port map (
            O => \N__44239\,
            I => \N__44227\
        );

    \I__7636\ : Sp12to4
    port map (
            O => \N__44236\,
            I => \N__44217\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__44233\,
            I => \N__44217\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__44230\,
            I => \N__44217\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__44227\,
            I => \N__44214\
        );

    \I__7632\ : InMux
    port map (
            O => \N__44226\,
            I => \N__44209\
        );

    \I__7631\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44209\
        );

    \I__7630\ : InMux
    port map (
            O => \N__44224\,
            I => \N__44206\
        );

    \I__7629\ : Odrv12
    port map (
            O => \N__44217\,
            I => n628
        );

    \I__7628\ : Odrv12
    port map (
            O => \N__44214\,
            I => n628
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__44209\,
            I => n628
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__44206\,
            I => n628
        );

    \I__7625\ : CascadeMux
    port map (
            O => \N__44197\,
            I => \foc.u_Park_Transform.n18_cascade_\
        );

    \I__7624\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44191\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__44191\,
            I => \foc.u_Park_Transform.n19845\
        );

    \I__7622\ : InMux
    port map (
            O => \N__44188\,
            I => \N__44183\
        );

    \I__7621\ : InMux
    port map (
            O => \N__44187\,
            I => \N__44178\
        );

    \I__7620\ : InMux
    port map (
            O => \N__44186\,
            I => \N__44178\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__44183\,
            I => \N__44175\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__44178\,
            I => \N__44172\
        );

    \I__7617\ : Odrv12
    port map (
            O => \N__44175\,
            I => \foc.u_Park_Transform.n26\
        );

    \I__7616\ : Odrv12
    port map (
            O => \N__44172\,
            I => \foc.u_Park_Transform.n26\
        );

    \I__7615\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44161\
        );

    \I__7614\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44161\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__44161\,
            I => \N__44158\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__44158\,
            I => \N__44155\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__44155\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_28\
        );

    \I__7610\ : InMux
    port map (
            O => \N__44152\,
            I => \N__44146\
        );

    \I__7609\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44146\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__44146\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n4\
        );

    \I__7607\ : InMux
    port map (
            O => \N__44143\,
            I => \N__44133\
        );

    \I__7606\ : InMux
    port map (
            O => \N__44142\,
            I => \N__44133\
        );

    \I__7605\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44130\
        );

    \I__7604\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44123\
        );

    \I__7603\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44123\
        );

    \I__7602\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44123\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__44133\,
            I => \N__44116\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__44130\,
            I => \N__44116\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__44123\,
            I => \N__44116\
        );

    \I__7598\ : Span4Mux_v
    port map (
            O => \N__44116\,
            I => \N__44111\
        );

    \I__7597\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44108\
        );

    \I__7596\ : InMux
    port map (
            O => \N__44114\,
            I => \N__44105\
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__44111\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__44108\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__44105\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__44098\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n4_cascade_\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__44095\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19269_cascade_\
        );

    \I__7590\ : CascadeMux
    port map (
            O => \N__44092\,
            I => \N__44088\
        );

    \I__7589\ : CascadeMux
    port map (
            O => \N__44091\,
            I => \N__44083\
        );

    \I__7588\ : InMux
    port map (
            O => \N__44088\,
            I => \N__44078\
        );

    \I__7587\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44078\
        );

    \I__7586\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44073\
        );

    \I__7585\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44073\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__44078\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n12\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__44073\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n12\
        );

    \I__7582\ : InMux
    port map (
            O => \N__44068\,
            I => \N__44065\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__44065\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19273\
        );

    \I__7580\ : InMux
    port map (
            O => \N__44062\,
            I => \N__44047\
        );

    \I__7579\ : InMux
    port map (
            O => \N__44061\,
            I => \N__44047\
        );

    \I__7578\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44047\
        );

    \I__7577\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44047\
        );

    \I__7576\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44042\
        );

    \I__7575\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44042\
        );

    \I__7574\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44039\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__44047\,
            I => n142_adj_2419
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__44042\,
            I => n142_adj_2419
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__44039\,
            I => n142_adj_2419
        );

    \I__7570\ : CascadeMux
    port map (
            O => \N__44032\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19273_cascade_\
        );

    \I__7569\ : InMux
    port map (
            O => \N__44029\,
            I => \N__44026\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__44026\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19269\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__44023\,
            I => \N__44020\
        );

    \I__7566\ : InMux
    port map (
            O => \N__44020\,
            I => \N__44017\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__44017\,
            I => \N__44014\
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__44014\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n283\
        );

    \I__7563\ : InMux
    port map (
            O => \N__44011\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18170\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__44008\,
            I => \N__44004\
        );

    \I__7561\ : CascadeMux
    port map (
            O => \N__44007\,
            I => \N__44000\
        );

    \I__7560\ : InMux
    port map (
            O => \N__44004\,
            I => \N__43995\
        );

    \I__7559\ : InMux
    port map (
            O => \N__44003\,
            I => \N__43995\
        );

    \I__7558\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43992\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__43995\,
            I => \N__43987\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__43992\,
            I => \N__43987\
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__43987\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n332\
        );

    \I__7554\ : InMux
    port map (
            O => \N__43984\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18171\
        );

    \I__7553\ : InMux
    port map (
            O => \N__43981\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18172\
        );

    \I__7552\ : InMux
    port map (
            O => \N__43978\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n787\
        );

    \I__7551\ : InMux
    port map (
            O => \N__43975\,
            I => \N__43972\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__43972\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n188\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__43969\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n138_cascade_\
        );

    \I__7548\ : InMux
    port map (
            O => \N__43966\,
            I => \N__43963\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__43963\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n139\
        );

    \I__7546\ : CascadeMux
    port map (
            O => \N__43960\,
            I => \N__43956\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__43959\,
            I => \N__43953\
        );

    \I__7544\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43949\
        );

    \I__7543\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43944\
        );

    \I__7542\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43944\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__43949\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n237\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__43944\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n237\
        );

    \I__7539\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43933\
        );

    \I__7538\ : InMux
    port map (
            O => \N__43938\,
            I => \N__43933\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43930\
        );

    \I__7536\ : Span4Mux_v
    port map (
            O => \N__43930\,
            I => \N__43927\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__43927\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_27\
        );

    \I__7534\ : InMux
    port map (
            O => \N__43924\,
            I => \N__43918\
        );

    \I__7533\ : InMux
    port map (
            O => \N__43923\,
            I => \N__43918\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__43918\,
            I => \N__43915\
        );

    \I__7531\ : Odrv12
    port map (
            O => \N__43915\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_21\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__43912\,
            I => \N__43909\
        );

    \I__7529\ : InMux
    port map (
            O => \N__43909\,
            I => \N__43906\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__43906\,
            I => \N__43903\
        );

    \I__7527\ : Sp12to4
    port map (
            O => \N__43903\,
            I => \N__43900\
        );

    \I__7526\ : Odrv12
    port map (
            O => \N__43900\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n87_adj_400\
        );

    \I__7525\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43894\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__43894\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n90\
        );

    \I__7523\ : InMux
    port map (
            O => \N__43891\,
            I => \N__43888\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__43888\,
            I => \N__43885\
        );

    \I__7521\ : Odrv4
    port map (
            O => \N__43885\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n136_adj_399\
        );

    \I__7520\ : InMux
    port map (
            O => \N__43882\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18167\
        );

    \I__7519\ : CascadeMux
    port map (
            O => \N__43879\,
            I => \N__43876\
        );

    \I__7518\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43873\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__43873\,
            I => \N__43870\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__43870\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n185_adj_398\
        );

    \I__7515\ : InMux
    port map (
            O => \N__43867\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18168\
        );

    \I__7514\ : InMux
    port map (
            O => \N__43864\,
            I => \N__43861\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__43861\,
            I => \N__43858\
        );

    \I__7512\ : Odrv4
    port map (
            O => \N__43858\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n234_adj_397\
        );

    \I__7511\ : InMux
    port map (
            O => \N__43855\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18169\
        );

    \I__7510\ : InMux
    port map (
            O => \N__43852\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18138\
        );

    \I__7509\ : InMux
    port map (
            O => \N__43849\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18139\
        );

    \I__7508\ : InMux
    port map (
            O => \N__43846\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18140\
        );

    \I__7507\ : InMux
    port map (
            O => \N__43843\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18141\
        );

    \I__7506\ : InMux
    port map (
            O => \N__43840\,
            I => \bfn_17_6_0_\
        );

    \I__7505\ : InMux
    port map (
            O => \N__43837\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349\
        );

    \I__7504\ : InMux
    port map (
            O => \N__43834\,
            I => \N__43828\
        );

    \I__7503\ : InMux
    port map (
            O => \N__43833\,
            I => \N__43828\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__43828\,
            I => \N__43825\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__43825\,
            I => \N__43822\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__43822\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_26\
        );

    \I__7499\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43816\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__43816\,
            I => \N__43813\
        );

    \I__7497\ : Odrv12
    port map (
            O => \N__43813\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n596_adj_703\
        );

    \I__7496\ : CascadeMux
    port map (
            O => \N__43810\,
            I => \N__43807\
        );

    \I__7495\ : InMux
    port map (
            O => \N__43807\,
            I => \N__43804\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43801\
        );

    \I__7493\ : Odrv12
    port map (
            O => \N__43801\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n642\
        );

    \I__7492\ : InMux
    port map (
            O => \N__43798\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18013\
        );

    \I__7491\ : InMux
    port map (
            O => \N__43795\,
            I => \N__43792\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__43792\,
            I => \N__43789\
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__43789\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n645_adj_702\
        );

    \I__7488\ : InMux
    port map (
            O => \N__43786\,
            I => \N__43783\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__43783\,
            I => \N__43780\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__43780\,
            I => \N__43777\
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__43777\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n691_adj_717\
        );

    \I__7484\ : InMux
    port map (
            O => \N__43774\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18014\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__43771\,
            I => \N__43768\
        );

    \I__7482\ : InMux
    port map (
            O => \N__43768\,
            I => \N__43765\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__43765\,
            I => \N__43762\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__43762\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n694_adj_701\
        );

    \I__7479\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43756\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__43756\,
            I => \N__43753\
        );

    \I__7477\ : Span12Mux_h
    port map (
            O => \N__43753\,
            I => \N__43750\
        );

    \I__7476\ : Odrv12
    port map (
            O => \N__43750\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n742_adj_715\
        );

    \I__7475\ : InMux
    port map (
            O => \N__43747\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18015\
        );

    \I__7474\ : InMux
    port map (
            O => \N__43744\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__43741\,
            I => \N__43738\
        );

    \I__7472\ : InMux
    port map (
            O => \N__43738\,
            I => \N__43735\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__43735\,
            I => \N__43732\
        );

    \I__7470\ : Span12Mux_v
    port map (
            O => \N__43732\,
            I => \N__43729\
        );

    \I__7469\ : Odrv12
    port map (
            O => \N__43729\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_CO\
        );

    \I__7468\ : InMux
    port map (
            O => \N__43726\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18135\
        );

    \I__7467\ : InMux
    port map (
            O => \N__43723\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18136\
        );

    \I__7466\ : InMux
    port map (
            O => \N__43720\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18137\
        );

    \I__7465\ : InMux
    port map (
            O => \N__43717\,
            I => \N__43714\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__43714\,
            I => \N__43711\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__43711\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n204_adj_711\
        );

    \I__7462\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43705\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__43705\,
            I => \N__43702\
        );

    \I__7460\ : Odrv12
    port map (
            O => \N__43702\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n250\
        );

    \I__7459\ : InMux
    port map (
            O => \N__43699\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18005\
        );

    \I__7458\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43693\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__43693\,
            I => \N__43690\
        );

    \I__7456\ : Odrv4
    port map (
            O => \N__43690\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n253_adj_710\
        );

    \I__7455\ : CascadeMux
    port map (
            O => \N__43687\,
            I => \N__43684\
        );

    \I__7454\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43681\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__43681\,
            I => \N__43678\
        );

    \I__7452\ : Odrv12
    port map (
            O => \N__43678\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n299\
        );

    \I__7451\ : InMux
    port map (
            O => \N__43675\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18006\
        );

    \I__7450\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43669\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__43669\,
            I => \N__43666\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__43666\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n302_adj_709\
        );

    \I__7447\ : InMux
    port map (
            O => \N__43663\,
            I => \N__43660\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__43660\,
            I => \N__43657\
        );

    \I__7445\ : Odrv12
    port map (
            O => \N__43657\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n348\
        );

    \I__7444\ : InMux
    port map (
            O => \N__43654\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18007\
        );

    \I__7443\ : InMux
    port map (
            O => \N__43651\,
            I => \N__43648\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__43648\,
            I => \N__43645\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__43645\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n351_adj_708\
        );

    \I__7440\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43639\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__43639\,
            I => \N__43636\
        );

    \I__7438\ : Odrv12
    port map (
            O => \N__43636\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n397\
        );

    \I__7437\ : InMux
    port map (
            O => \N__43633\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18008\
        );

    \I__7436\ : InMux
    port map (
            O => \N__43630\,
            I => \N__43627\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__43627\,
            I => \N__43624\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__43624\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n400_adj_707\
        );

    \I__7433\ : InMux
    port map (
            O => \N__43621\,
            I => \N__43618\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__43618\,
            I => \N__43615\
        );

    \I__7431\ : Odrv12
    port map (
            O => \N__43615\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n446\
        );

    \I__7430\ : InMux
    port map (
            O => \N__43612\,
            I => \bfn_16_28_0_\
        );

    \I__7429\ : InMux
    port map (
            O => \N__43609\,
            I => \N__43606\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__43606\,
            I => \N__43603\
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__43603\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n449_adj_706\
        );

    \I__7426\ : InMux
    port map (
            O => \N__43600\,
            I => \N__43597\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43594\
        );

    \I__7424\ : Odrv12
    port map (
            O => \N__43594\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n495\
        );

    \I__7423\ : InMux
    port map (
            O => \N__43591\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18010\
        );

    \I__7422\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43585\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__43585\,
            I => \N__43582\
        );

    \I__7420\ : Odrv4
    port map (
            O => \N__43582\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n498_adj_705\
        );

    \I__7419\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43576\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__43576\,
            I => \N__43573\
        );

    \I__7417\ : Odrv12
    port map (
            O => \N__43573\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n544\
        );

    \I__7416\ : InMux
    port map (
            O => \N__43570\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18011\
        );

    \I__7415\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43564\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__43564\,
            I => \N__43561\
        );

    \I__7413\ : Odrv12
    port map (
            O => \N__43561\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n547_adj_704\
        );

    \I__7412\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43555\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__43555\,
            I => \N__43552\
        );

    \I__7410\ : Odrv12
    port map (
            O => \N__43552\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n593\
        );

    \I__7409\ : InMux
    port map (
            O => \N__43549\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18012\
        );

    \I__7408\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43543\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__43543\,
            I => \N__43540\
        );

    \I__7406\ : Odrv12
    port map (
            O => \N__43540\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n599_adj_687\
        );

    \I__7405\ : InMux
    port map (
            O => \N__43537\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18028\
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__43534\,
            I => \N__43531\
        );

    \I__7403\ : InMux
    port map (
            O => \N__43531\,
            I => \N__43528\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__43528\,
            I => \N__43525\
        );

    \I__7401\ : Odrv12
    port map (
            O => \N__43525\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n648_adj_686\
        );

    \I__7400\ : InMux
    port map (
            O => \N__43522\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18029\
        );

    \I__7399\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43516\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__43516\,
            I => \N__43513\
        );

    \I__7397\ : Odrv12
    port map (
            O => \N__43513\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n697_adj_685\
        );

    \I__7396\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43507\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__43507\,
            I => \N__43504\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__43504\,
            I => \N__43501\
        );

    \I__7393\ : Span4Mux_v
    port map (
            O => \N__43501\,
            I => \N__43498\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__43498\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n746_adj_699\
        );

    \I__7391\ : InMux
    port map (
            O => \N__43495\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18030\
        );

    \I__7390\ : InMux
    port map (
            O => \N__43492\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700\
        );

    \I__7389\ : CascadeMux
    port map (
            O => \N__43489\,
            I => \N__43486\
        );

    \I__7388\ : InMux
    port map (
            O => \N__43486\,
            I => \N__43483\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__43483\,
            I => \N__43480\
        );

    \I__7386\ : Span4Mux_h
    port map (
            O => \N__43480\,
            I => \N__43477\
        );

    \I__7385\ : Span4Mux_v
    port map (
            O => \N__43477\,
            I => \N__43474\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__43474\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_CO\
        );

    \I__7383\ : CascadeMux
    port map (
            O => \N__43471\,
            I => \N__43468\
        );

    \I__7382\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43465\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__43465\,
            I => \N__43462\
        );

    \I__7380\ : Span4Mux_v
    port map (
            O => \N__43462\,
            I => \N__43459\
        );

    \I__7379\ : Odrv4
    port map (
            O => \N__43459\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n54\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__43456\,
            I => \N__43453\
        );

    \I__7377\ : InMux
    port map (
            O => \N__43453\,
            I => \N__43450\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__43450\,
            I => \N__43447\
        );

    \I__7375\ : Odrv4
    port map (
            O => \N__43447\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n57_adj_714\
        );

    \I__7374\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43441\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__43441\,
            I => \N__43438\
        );

    \I__7372\ : Odrv12
    port map (
            O => \N__43438\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n103\
        );

    \I__7371\ : InMux
    port map (
            O => \N__43435\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18002\
        );

    \I__7370\ : InMux
    port map (
            O => \N__43432\,
            I => \N__43429\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__43429\,
            I => \N__43426\
        );

    \I__7368\ : Odrv4
    port map (
            O => \N__43426\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n106_adj_713\
        );

    \I__7367\ : CascadeMux
    port map (
            O => \N__43423\,
            I => \N__43420\
        );

    \I__7366\ : InMux
    port map (
            O => \N__43420\,
            I => \N__43417\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43414\
        );

    \I__7364\ : Odrv12
    port map (
            O => \N__43414\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n152\
        );

    \I__7363\ : InMux
    port map (
            O => \N__43411\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18003\
        );

    \I__7362\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43405\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__43405\,
            I => \N__43402\
        );

    \I__7360\ : Odrv12
    port map (
            O => \N__43402\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n155_adj_712\
        );

    \I__7359\ : InMux
    port map (
            O => \N__43399\,
            I => \N__43396\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__43396\,
            I => \N__43393\
        );

    \I__7357\ : Odrv12
    port map (
            O => \N__43393\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n201\
        );

    \I__7356\ : InMux
    port map (
            O => \N__43390\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18004\
        );

    \I__7355\ : CascadeMux
    port map (
            O => \N__43387\,
            I => \N__43384\
        );

    \I__7354\ : InMux
    port map (
            O => \N__43384\,
            I => \N__43381\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43378\
        );

    \I__7352\ : Odrv12
    port map (
            O => \N__43378\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n158_adj_696\
        );

    \I__7351\ : InMux
    port map (
            O => \N__43375\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18019\
        );

    \I__7350\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43369\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__43369\,
            I => \N__43366\
        );

    \I__7348\ : Odrv4
    port map (
            O => \N__43366\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n207_adj_695\
        );

    \I__7347\ : InMux
    port map (
            O => \N__43363\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18020\
        );

    \I__7346\ : CascadeMux
    port map (
            O => \N__43360\,
            I => \N__43357\
        );

    \I__7345\ : InMux
    port map (
            O => \N__43357\,
            I => \N__43354\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__43354\,
            I => \N__43351\
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__43351\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n256_adj_694\
        );

    \I__7342\ : InMux
    port map (
            O => \N__43348\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18021\
        );

    \I__7341\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43342\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__43342\,
            I => \N__43339\
        );

    \I__7339\ : Odrv12
    port map (
            O => \N__43339\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n305_adj_693\
        );

    \I__7338\ : InMux
    port map (
            O => \N__43336\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18022\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__43333\,
            I => \N__43330\
        );

    \I__7336\ : InMux
    port map (
            O => \N__43330\,
            I => \N__43327\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__43327\,
            I => \N__43324\
        );

    \I__7334\ : Odrv4
    port map (
            O => \N__43324\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n354_adj_692\
        );

    \I__7333\ : InMux
    port map (
            O => \N__43321\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18023\
        );

    \I__7332\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43315\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__43315\,
            I => \N__43312\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__43312\,
            I => \N__43309\
        );

    \I__7329\ : Odrv4
    port map (
            O => \N__43309\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n403_adj_691\
        );

    \I__7328\ : InMux
    port map (
            O => \N__43306\,
            I => \bfn_16_26_0_\
        );

    \I__7327\ : CascadeMux
    port map (
            O => \N__43303\,
            I => \N__43300\
        );

    \I__7326\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43297\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43294\
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__43294\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n452_adj_690\
        );

    \I__7323\ : InMux
    port map (
            O => \N__43291\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18025\
        );

    \I__7322\ : InMux
    port map (
            O => \N__43288\,
            I => \N__43285\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__43285\,
            I => \N__43282\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__43282\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n501_adj_689\
        );

    \I__7319\ : InMux
    port map (
            O => \N__43279\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18026\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__43276\,
            I => \N__43273\
        );

    \I__7317\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43270\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__43270\,
            I => \N__43267\
        );

    \I__7315\ : Odrv12
    port map (
            O => \N__43267\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n550_adj_688\
        );

    \I__7314\ : InMux
    port map (
            O => \N__43264\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18027\
        );

    \I__7313\ : InMux
    port map (
            O => \N__43261\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17996\
        );

    \I__7312\ : InMux
    port map (
            O => \N__43258\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17997\
        );

    \I__7311\ : InMux
    port map (
            O => \N__43255\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17998\
        );

    \I__7310\ : InMux
    port map (
            O => \N__43252\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17999\
        );

    \I__7309\ : CascadeMux
    port map (
            O => \N__43249\,
            I => \N__43246\
        );

    \I__7308\ : InMux
    port map (
            O => \N__43246\,
            I => \N__43242\
        );

    \I__7307\ : InMux
    port map (
            O => \N__43245\,
            I => \N__43239\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__43242\,
            I => \N__43234\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__43239\,
            I => \N__43234\
        );

    \I__7304\ : Span4Mux_v
    port map (
            O => \N__43234\,
            I => \N__43231\
        );

    \I__7303\ : Odrv4
    port map (
            O => \N__43231\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n738_adj_718\
        );

    \I__7302\ : InMux
    port map (
            O => \N__43228\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18000\
        );

    \I__7301\ : InMux
    port map (
            O => \N__43225\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n739\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__43222\,
            I => \N__43219\
        );

    \I__7299\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43216\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__43216\,
            I => \N__43213\
        );

    \I__7297\ : Span4Mux_h
    port map (
            O => \N__43213\,
            I => \N__43210\
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__43210\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_CO\
        );

    \I__7295\ : CascadeMux
    port map (
            O => \N__43207\,
            I => \N__43204\
        );

    \I__7294\ : InMux
    port map (
            O => \N__43204\,
            I => \N__43201\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__43201\,
            I => \N__43198\
        );

    \I__7292\ : Odrv12
    port map (
            O => \N__43198\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n60_adj_698\
        );

    \I__7291\ : InMux
    port map (
            O => \N__43195\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18017\
        );

    \I__7290\ : InMux
    port map (
            O => \N__43192\,
            I => \N__43189\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__43189\,
            I => \N__43186\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__43186\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n109_adj_697\
        );

    \I__7287\ : InMux
    port map (
            O => \N__43183\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18018\
        );

    \I__7286\ : InMux
    port map (
            O => \N__43180\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17987\
        );

    \I__7285\ : InMux
    port map (
            O => \N__43177\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17988\
        );

    \I__7284\ : InMux
    port map (
            O => \N__43174\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17989\
        );

    \I__7283\ : InMux
    port map (
            O => \N__43171\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17990\
        );

    \I__7282\ : InMux
    port map (
            O => \N__43168\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17991\
        );

    \I__7281\ : InMux
    port map (
            O => \N__43165\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17992\
        );

    \I__7280\ : InMux
    port map (
            O => \N__43162\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17993\
        );

    \I__7279\ : InMux
    port map (
            O => \N__43159\,
            I => \bfn_16_24_0_\
        );

    \I__7278\ : InMux
    port map (
            O => \N__43156\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17995\
        );

    \I__7277\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43147\
        );

    \I__7276\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43147\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__43147\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_27\
        );

    \I__7274\ : InMux
    port map (
            O => \N__43144\,
            I => \N__43138\
        );

    \I__7273\ : InMux
    port map (
            O => \N__43143\,
            I => \N__43138\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__43138\,
            I => \N__43135\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__43135\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_25\
        );

    \I__7270\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43126\
        );

    \I__7269\ : InMux
    port map (
            O => \N__43131\,
            I => \N__43126\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__43126\,
            I => \N__43123\
        );

    \I__7267\ : Odrv12
    port map (
            O => \N__43123\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_22\
        );

    \I__7266\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43117\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__43117\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n7\
        );

    \I__7264\ : InMux
    port map (
            O => \N__43114\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15742\
        );

    \I__7263\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43108\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__43108\,
            I => \N__43105\
        );

    \I__7261\ : Span4Mux_v
    port map (
            O => \N__43105\,
            I => \N__43102\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__43102\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n6\
        );

    \I__7259\ : InMux
    port map (
            O => \N__43099\,
            I => \bfn_16_21_0_\
        );

    \I__7258\ : InMux
    port map (
            O => \N__43096\,
            I => \N__43093\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__43093\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n5\
        );

    \I__7256\ : InMux
    port map (
            O => \N__43090\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15744\
        );

    \I__7255\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43084\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__43084\,
            I => \N__43081\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__43081\,
            I => \N__43078\
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__43078\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4\
        );

    \I__7251\ : InMux
    port map (
            O => \N__43075\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15745\
        );

    \I__7250\ : InMux
    port map (
            O => \N__43072\,
            I => \N__43069\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__43069\,
            I => \N__43066\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__43066\,
            I => \N__43063\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__43063\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n3\
        );

    \I__7246\ : InMux
    port map (
            O => \N__43060\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15746\
        );

    \I__7245\ : InMux
    port map (
            O => \N__43057\,
            I => \N__43054\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__43054\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n2\
        );

    \I__7243\ : InMux
    port map (
            O => \N__43051\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15747\
        );

    \I__7242\ : InMux
    port map (
            O => \N__43048\,
            I => \N__43045\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__43045\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n188_adj_725\
        );

    \I__7240\ : CascadeMux
    port map (
            O => \N__43042\,
            I => \N__43038\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__43041\,
            I => \N__43035\
        );

    \I__7238\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43031\
        );

    \I__7237\ : InMux
    port map (
            O => \N__43035\,
            I => \N__43026\
        );

    \I__7236\ : InMux
    port map (
            O => \N__43034\,
            I => \N__43026\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__43031\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__43026\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720\
        );

    \I__7233\ : InMux
    port map (
            O => \N__43021\,
            I => \N__43018\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__43018\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15\
        );

    \I__7231\ : InMux
    port map (
            O => \N__43015\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15734\
        );

    \I__7230\ : InMux
    port map (
            O => \N__43012\,
            I => \N__43009\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__43009\,
            I => \N__43006\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__43006\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n14\
        );

    \I__7227\ : InMux
    port map (
            O => \N__43003\,
            I => \bfn_16_20_0_\
        );

    \I__7226\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42997\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__42997\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n13\
        );

    \I__7224\ : InMux
    port map (
            O => \N__42994\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15736\
        );

    \I__7223\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42988\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__42988\,
            I => \N__42985\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__42985\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n12\
        );

    \I__7220\ : InMux
    port map (
            O => \N__42982\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15737\
        );

    \I__7219\ : InMux
    port map (
            O => \N__42979\,
            I => \N__42976\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__42976\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n11\
        );

    \I__7217\ : InMux
    port map (
            O => \N__42973\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15738\
        );

    \I__7216\ : InMux
    port map (
            O => \N__42970\,
            I => \N__42967\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__42967\,
            I => \N__42964\
        );

    \I__7214\ : Odrv12
    port map (
            O => \N__42964\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n10\
        );

    \I__7213\ : InMux
    port map (
            O => \N__42961\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15739\
        );

    \I__7212\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42955\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__42955\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n9\
        );

    \I__7210\ : InMux
    port map (
            O => \N__42952\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15740\
        );

    \I__7209\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42946\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__42946\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n8\
        );

    \I__7207\ : InMux
    port map (
            O => \N__42943\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15741\
        );

    \I__7206\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42937\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__42937\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n24\
        );

    \I__7204\ : InMux
    port map (
            O => \N__42934\,
            I => \N__42931\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__42931\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n23\
        );

    \I__7202\ : InMux
    port map (
            O => \N__42928\,
            I => \N__42925\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__42925\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n22\
        );

    \I__7200\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42919\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__42919\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_adj_752\
        );

    \I__7198\ : InMux
    port map (
            O => \N__42916\,
            I => \N__42913\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__42913\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20\
        );

    \I__7196\ : InMux
    port map (
            O => \N__42910\,
            I => \N__42907\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__42907\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19\
        );

    \I__7194\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42901\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__42901\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_751\
        );

    \I__7192\ : InMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__42895\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17\
        );

    \I__7190\ : InMux
    port map (
            O => \N__42892\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15732\
        );

    \I__7189\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42886\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__42886\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n16\
        );

    \I__7187\ : InMux
    port map (
            O => \N__42883\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15733\
        );

    \I__7186\ : InMux
    port map (
            O => \N__42880\,
            I => \N__42877\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__42877\,
            I => \N__42874\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__42874\,
            I => \foc.qCurrent_5\
        );

    \I__7183\ : InMux
    port map (
            O => \N__42871\,
            I => \N__42868\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__42868\,
            I => \N__42865\
        );

    \I__7181\ : Odrv4
    port map (
            O => \N__42865\,
            I => \foc.qCurrent_9\
        );

    \I__7180\ : InMux
    port map (
            O => \N__42862\,
            I => \N__42859\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__42859\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n30\
        );

    \I__7178\ : InMux
    port map (
            O => \N__42856\,
            I => \N__42853\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__42853\,
            I => \N__42850\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__42850\,
            I => \N__42846\
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__42849\,
            I => \N__42843\
        );

    \I__7174\ : Sp12to4
    port map (
            O => \N__42846\,
            I => \N__42840\
        );

    \I__7173\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42837\
        );

    \I__7172\ : Span12Mux_h
    port map (
            O => \N__42840\,
            I => \N__42834\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__42837\,
            I => \N__42831\
        );

    \I__7170\ : Odrv12
    port map (
            O => \N__42834\,
            I => \foc.u_DQ_Current_Control.n31\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__42831\,
            I => \foc.u_DQ_Current_Control.n31\
        );

    \I__7168\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42823\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__42823\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n29\
        );

    \I__7166\ : InMux
    port map (
            O => \N__42820\,
            I => \N__42817\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__42817\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n28\
        );

    \I__7164\ : InMux
    port map (
            O => \N__42814\,
            I => \N__42811\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__42811\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n27_adj_753\
        );

    \I__7162\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42805\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__42805\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n26\
        );

    \I__7160\ : InMux
    port map (
            O => \N__42802\,
            I => \N__42799\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__42799\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n25\
        );

    \I__7158\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42793\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__42793\,
            I => \N__42790\
        );

    \I__7156\ : Span4Mux_v
    port map (
            O => \N__42790\,
            I => \N__42786\
        );

    \I__7155\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42783\
        );

    \I__7154\ : Span4Mux_v
    port map (
            O => \N__42786\,
            I => \N__42778\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__42783\,
            I => \N__42778\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__42778\,
            I => \N__42775\
        );

    \I__7151\ : Odrv4
    port map (
            O => \N__42775\,
            I => \foc.u_Park_Transform.n745\
        );

    \I__7150\ : CascadeMux
    port map (
            O => \N__42772\,
            I => \N__42769\
        );

    \I__7149\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42766\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__42766\,
            I => \foc.u_Park_Transform.n697\
        );

    \I__7147\ : InMux
    port map (
            O => \N__42763\,
            I => \N__42760\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__42760\,
            I => \N__42757\
        );

    \I__7145\ : Span4Mux_h
    port map (
            O => \N__42757\,
            I => \N__42754\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__42754\,
            I => \foc.u_Park_Transform.n746_adj_2011\
        );

    \I__7143\ : InMux
    port map (
            O => \N__42751\,
            I => \foc.u_Park_Transform.n17051\
        );

    \I__7142\ : InMux
    port map (
            O => \N__42748\,
            I => \foc.u_Park_Transform.n747_adj_2012\
        );

    \I__7141\ : CascadeMux
    port map (
            O => \N__42745\,
            I => \N__42742\
        );

    \I__7140\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42739\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__42739\,
            I => \N__42736\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__42736\,
            I => \N__42733\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__42733\,
            I => \N__42730\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__42730\,
            I => \foc.u_Park_Transform.n747_adj_2012_THRU_CO\
        );

    \I__7135\ : CascadeMux
    port map (
            O => \N__42727\,
            I => \foc.u_Park_Transform.n6_cascade_\
        );

    \I__7134\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42721\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__42721\,
            I => \N__42718\
        );

    \I__7132\ : Span4Mux_v
    port map (
            O => \N__42718\,
            I => \N__42715\
        );

    \I__7131\ : Sp12to4
    port map (
            O => \N__42715\,
            I => \N__42711\
        );

    \I__7130\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42708\
        );

    \I__7129\ : Odrv12
    port map (
            O => \N__42711\,
            I => \foc.Look_Up_Table_out1_1_2\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__42708\,
            I => \foc.Look_Up_Table_out1_1_2\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__42703\,
            I => \N__42693\
        );

    \I__7126\ : CascadeMux
    port map (
            O => \N__42702\,
            I => \N__42689\
        );

    \I__7125\ : CascadeMux
    port map (
            O => \N__42701\,
            I => \N__42685\
        );

    \I__7124\ : CascadeMux
    port map (
            O => \N__42700\,
            I => \N__42680\
        );

    \I__7123\ : CascadeMux
    port map (
            O => \N__42699\,
            I => \N__42677\
        );

    \I__7122\ : CascadeMux
    port map (
            O => \N__42698\,
            I => \N__42674\
        );

    \I__7121\ : CascadeMux
    port map (
            O => \N__42697\,
            I => \N__42671\
        );

    \I__7120\ : CascadeMux
    port map (
            O => \N__42696\,
            I => \N__42667\
        );

    \I__7119\ : InMux
    port map (
            O => \N__42693\,
            I => \N__42653\
        );

    \I__7118\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42653\
        );

    \I__7117\ : InMux
    port map (
            O => \N__42689\,
            I => \N__42653\
        );

    \I__7116\ : InMux
    port map (
            O => \N__42688\,
            I => \N__42653\
        );

    \I__7115\ : InMux
    port map (
            O => \N__42685\,
            I => \N__42653\
        );

    \I__7114\ : InMux
    port map (
            O => \N__42684\,
            I => \N__42653\
        );

    \I__7113\ : InMux
    port map (
            O => \N__42683\,
            I => \N__42648\
        );

    \I__7112\ : InMux
    port map (
            O => \N__42680\,
            I => \N__42648\
        );

    \I__7111\ : InMux
    port map (
            O => \N__42677\,
            I => \N__42645\
        );

    \I__7110\ : InMux
    port map (
            O => \N__42674\,
            I => \N__42634\
        );

    \I__7109\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42634\
        );

    \I__7108\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42634\
        );

    \I__7107\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42634\
        );

    \I__7106\ : InMux
    port map (
            O => \N__42666\,
            I => \N__42634\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__42653\,
            I => \N__42623\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__42648\,
            I => \N__42623\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__42645\,
            I => \N__42618\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__42634\,
            I => \N__42618\
        );

    \I__7101\ : InMux
    port map (
            O => \N__42633\,
            I => \N__42615\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__42632\,
            I => \N__42612\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__42631\,
            I => \N__42608\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__42630\,
            I => \N__42604\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__42629\,
            I => \N__42600\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__42628\,
            I => \N__42597\
        );

    \I__7095\ : Span4Mux_h
    port map (
            O => \N__42623\,
            I => \N__42590\
        );

    \I__7094\ : Span4Mux_h
    port map (
            O => \N__42618\,
            I => \N__42585\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__42615\,
            I => \N__42585\
        );

    \I__7092\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42570\
        );

    \I__7091\ : InMux
    port map (
            O => \N__42611\,
            I => \N__42570\
        );

    \I__7090\ : InMux
    port map (
            O => \N__42608\,
            I => \N__42570\
        );

    \I__7089\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42570\
        );

    \I__7088\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42570\
        );

    \I__7087\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42570\
        );

    \I__7086\ : InMux
    port map (
            O => \N__42600\,
            I => \N__42570\
        );

    \I__7085\ : InMux
    port map (
            O => \N__42597\,
            I => \N__42567\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__42596\,
            I => \N__42564\
        );

    \I__7083\ : CascadeMux
    port map (
            O => \N__42595\,
            I => \N__42560\
        );

    \I__7082\ : CascadeMux
    port map (
            O => \N__42594\,
            I => \N__42556\
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__42593\,
            I => \N__42552\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__42590\,
            I => \N__42549\
        );

    \I__7079\ : Span4Mux_v
    port map (
            O => \N__42585\,
            I => \N__42542\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__42570\,
            I => \N__42542\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__42567\,
            I => \N__42542\
        );

    \I__7076\ : InMux
    port map (
            O => \N__42564\,
            I => \N__42529\
        );

    \I__7075\ : InMux
    port map (
            O => \N__42563\,
            I => \N__42529\
        );

    \I__7074\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42529\
        );

    \I__7073\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42529\
        );

    \I__7072\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42529\
        );

    \I__7071\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42529\
        );

    \I__7070\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42526\
        );

    \I__7069\ : Odrv4
    port map (
            O => \N__42549\,
            I => \foc.u_Park_Transform.n595\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__42542\,
            I => \foc.u_Park_Transform.n595\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__42529\,
            I => \foc.u_Park_Transform.n595\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__42526\,
            I => \foc.u_Park_Transform.n595\
        );

    \I__7065\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42511\
        );

    \I__7064\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42511\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__42511\,
            I => \N__42508\
        );

    \I__7062\ : Span4Mux_h
    port map (
            O => \N__42508\,
            I => \N__42504\
        );

    \I__7061\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42501\
        );

    \I__7060\ : Odrv4
    port map (
            O => \N__42504\,
            I => n4
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__42501\,
            I => n4
        );

    \I__7058\ : InMux
    port map (
            O => \N__42496\,
            I => \N__42493\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__42493\,
            I => \N__42490\
        );

    \I__7056\ : Odrv12
    port map (
            O => \N__42490\,
            I => \foc.qCurrent_10\
        );

    \I__7055\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42484\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42481\
        );

    \I__7053\ : Odrv12
    port map (
            O => \N__42481\,
            I => \foc.qCurrent_7\
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__42478\,
            I => \N__42475\
        );

    \I__7051\ : InMux
    port map (
            O => \N__42475\,
            I => \N__42472\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__42472\,
            I => \foc.u_Park_Transform.n305\
        );

    \I__7049\ : CascadeMux
    port map (
            O => \N__42469\,
            I => \N__42466\
        );

    \I__7048\ : InMux
    port map (
            O => \N__42466\,
            I => \N__42463\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__42463\,
            I => \N__42460\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__42460\,
            I => \foc.u_Park_Transform.n351\
        );

    \I__7045\ : InMux
    port map (
            O => \N__42457\,
            I => \foc.u_Park_Transform.n17043\
        );

    \I__7044\ : InMux
    port map (
            O => \N__42454\,
            I => \N__42451\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__42451\,
            I => \foc.u_Park_Transform.n354\
        );

    \I__7042\ : CascadeMux
    port map (
            O => \N__42448\,
            I => \N__42445\
        );

    \I__7041\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42442\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__42442\,
            I => \N__42439\
        );

    \I__7039\ : Span4Mux_v
    port map (
            O => \N__42439\,
            I => \N__42436\
        );

    \I__7038\ : Odrv4
    port map (
            O => \N__42436\,
            I => \foc.u_Park_Transform.n400\
        );

    \I__7037\ : InMux
    port map (
            O => \N__42433\,
            I => \foc.u_Park_Transform.n17044\
        );

    \I__7036\ : CascadeMux
    port map (
            O => \N__42430\,
            I => \N__42427\
        );

    \I__7035\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42424\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__42424\,
            I => \foc.u_Park_Transform.n403\
        );

    \I__7033\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42418\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__42418\,
            I => \N__42415\
        );

    \I__7031\ : Odrv4
    port map (
            O => \N__42415\,
            I => \foc.u_Park_Transform.n449\
        );

    \I__7030\ : InMux
    port map (
            O => \N__42412\,
            I => \bfn_16_14_0_\
        );

    \I__7029\ : InMux
    port map (
            O => \N__42409\,
            I => \N__42406\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__42406\,
            I => \foc.u_Park_Transform.n452\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__42403\,
            I => \N__42400\
        );

    \I__7026\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42397\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__42397\,
            I => \N__42394\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__42394\,
            I => \N__42391\
        );

    \I__7023\ : Odrv4
    port map (
            O => \N__42391\,
            I => \foc.u_Park_Transform.n498\
        );

    \I__7022\ : InMux
    port map (
            O => \N__42388\,
            I => \foc.u_Park_Transform.n17046\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__42385\,
            I => \N__42382\
        );

    \I__7020\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42379\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__42379\,
            I => \foc.u_Park_Transform.n501\
        );

    \I__7018\ : InMux
    port map (
            O => \N__42376\,
            I => \N__42373\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__42373\,
            I => \N__42370\
        );

    \I__7016\ : Odrv4
    port map (
            O => \N__42370\,
            I => \foc.u_Park_Transform.n547\
        );

    \I__7015\ : InMux
    port map (
            O => \N__42367\,
            I => \foc.u_Park_Transform.n17047\
        );

    \I__7014\ : InMux
    port map (
            O => \N__42364\,
            I => \N__42361\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__42361\,
            I => \foc.u_Park_Transform.n550\
        );

    \I__7012\ : CascadeMux
    port map (
            O => \N__42358\,
            I => \N__42355\
        );

    \I__7011\ : InMux
    port map (
            O => \N__42355\,
            I => \N__42352\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__42352\,
            I => \N__42349\
        );

    \I__7009\ : Odrv4
    port map (
            O => \N__42349\,
            I => \foc.u_Park_Transform.n596\
        );

    \I__7008\ : InMux
    port map (
            O => \N__42346\,
            I => \foc.u_Park_Transform.n17048\
        );

    \I__7007\ : CascadeMux
    port map (
            O => \N__42343\,
            I => \N__42340\
        );

    \I__7006\ : InMux
    port map (
            O => \N__42340\,
            I => \N__42337\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__42337\,
            I => \foc.u_Park_Transform.n599\
        );

    \I__7004\ : CascadeMux
    port map (
            O => \N__42334\,
            I => \N__42331\
        );

    \I__7003\ : InMux
    port map (
            O => \N__42331\,
            I => \N__42328\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__42328\,
            I => \N__42325\
        );

    \I__7001\ : Odrv4
    port map (
            O => \N__42325\,
            I => \foc.u_Park_Transform.n645\
        );

    \I__7000\ : InMux
    port map (
            O => \N__42322\,
            I => \foc.u_Park_Transform.n17049\
        );

    \I__6999\ : InMux
    port map (
            O => \N__42319\,
            I => \N__42316\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__42316\,
            I => \foc.u_Park_Transform.n648\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__42313\,
            I => \N__42310\
        );

    \I__6996\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42307\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__42307\,
            I => \N__42304\
        );

    \I__6994\ : Span4Mux_h
    port map (
            O => \N__42304\,
            I => \N__42301\
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__42301\,
            I => \foc.u_Park_Transform.n694\
        );

    \I__6992\ : InMux
    port map (
            O => \N__42298\,
            I => \foc.u_Park_Transform.n17050\
        );

    \I__6991\ : InMux
    port map (
            O => \N__42295\,
            I => \N__42292\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__42292\,
            I => \N__42288\
        );

    \I__6989\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42285\
        );

    \I__6988\ : Span4Mux_v
    port map (
            O => \N__42288\,
            I => \N__42282\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__42285\,
            I => \N__42279\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__42282\,
            I => \N__42276\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__42279\,
            I => \N__42273\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__42276\,
            I => \foc.u_Park_Transform.n749\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__42273\,
            I => \foc.u_Park_Transform.n749\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__42268\,
            I => \N__42265\
        );

    \I__6981\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42262\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__42262\,
            I => \N__42259\
        );

    \I__6979\ : Odrv12
    port map (
            O => \N__42259\,
            I => \foc.u_Park_Transform.n700_adj_2141\
        );

    \I__6978\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42253\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__42253\,
            I => \N__42250\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__42250\,
            I => \N__42247\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__42247\,
            I => \foc.u_Park_Transform.n750\
        );

    \I__6974\ : InMux
    port map (
            O => \N__42244\,
            I => \foc.u_Park_Transform.n17219\
        );

    \I__6973\ : InMux
    port map (
            O => \N__42241\,
            I => \foc.u_Park_Transform.n751_adj_2142\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__42238\,
            I => \N__42235\
        );

    \I__6971\ : InMux
    port map (
            O => \N__42235\,
            I => \N__42232\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__42232\,
            I => \N__42229\
        );

    \I__6969\ : Span4Mux_h
    port map (
            O => \N__42229\,
            I => \N__42226\
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__42226\,
            I => \foc.u_Park_Transform.n751_adj_2142_THRU_CO\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__42223\,
            I => \N__42212\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__42222\,
            I => \N__42208\
        );

    \I__6965\ : CascadeMux
    port map (
            O => \N__42221\,
            I => \N__42204\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__42220\,
            I => \N__42200\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__42219\,
            I => \N__42197\
        );

    \I__6962\ : CascadeMux
    port map (
            O => \N__42218\,
            I => \N__42194\
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__42217\,
            I => \N__42191\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__42216\,
            I => \N__42187\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__42215\,
            I => \N__42179\
        );

    \I__6958\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42164\
        );

    \I__6957\ : InMux
    port map (
            O => \N__42211\,
            I => \N__42164\
        );

    \I__6956\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42164\
        );

    \I__6955\ : InMux
    port map (
            O => \N__42207\,
            I => \N__42164\
        );

    \I__6954\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42164\
        );

    \I__6953\ : InMux
    port map (
            O => \N__42203\,
            I => \N__42164\
        );

    \I__6952\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42164\
        );

    \I__6951\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42161\
        );

    \I__6950\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42150\
        );

    \I__6949\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42150\
        );

    \I__6948\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42150\
        );

    \I__6947\ : InMux
    port map (
            O => \N__42187\,
            I => \N__42150\
        );

    \I__6946\ : InMux
    port map (
            O => \N__42186\,
            I => \N__42150\
        );

    \I__6945\ : CascadeMux
    port map (
            O => \N__42185\,
            I => \N__42147\
        );

    \I__6944\ : CascadeMux
    port map (
            O => \N__42184\,
            I => \N__42143\
        );

    \I__6943\ : CascadeMux
    port map (
            O => \N__42183\,
            I => \N__42139\
        );

    \I__6942\ : InMux
    port map (
            O => \N__42182\,
            I => \N__42131\
        );

    \I__6941\ : InMux
    port map (
            O => \N__42179\,
            I => \N__42127\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__42164\,
            I => \N__42120\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__42161\,
            I => \N__42120\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__42150\,
            I => \N__42120\
        );

    \I__6937\ : InMux
    port map (
            O => \N__42147\,
            I => \N__42107\
        );

    \I__6936\ : InMux
    port map (
            O => \N__42146\,
            I => \N__42107\
        );

    \I__6935\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42107\
        );

    \I__6934\ : InMux
    port map (
            O => \N__42142\,
            I => \N__42107\
        );

    \I__6933\ : InMux
    port map (
            O => \N__42139\,
            I => \N__42107\
        );

    \I__6932\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42107\
        );

    \I__6931\ : CascadeMux
    port map (
            O => \N__42137\,
            I => \N__42104\
        );

    \I__6930\ : CascadeMux
    port map (
            O => \N__42136\,
            I => \N__42100\
        );

    \I__6929\ : CascadeMux
    port map (
            O => \N__42135\,
            I => \N__42096\
        );

    \I__6928\ : CascadeMux
    port map (
            O => \N__42134\,
            I => \N__42092\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__42131\,
            I => \N__42088\
        );

    \I__6926\ : InMux
    port map (
            O => \N__42130\,
            I => \N__42085\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__42127\,
            I => \N__42082\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__42120\,
            I => \N__42077\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__42107\,
            I => \N__42077\
        );

    \I__6922\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42060\
        );

    \I__6921\ : InMux
    port map (
            O => \N__42103\,
            I => \N__42060\
        );

    \I__6920\ : InMux
    port map (
            O => \N__42100\,
            I => \N__42060\
        );

    \I__6919\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42060\
        );

    \I__6918\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42060\
        );

    \I__6917\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42060\
        );

    \I__6916\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42060\
        );

    \I__6915\ : InMux
    port map (
            O => \N__42091\,
            I => \N__42060\
        );

    \I__6914\ : Span4Mux_v
    port map (
            O => \N__42088\,
            I => \N__42057\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__42085\,
            I => \N__42054\
        );

    \I__6912\ : Span4Mux_v
    port map (
            O => \N__42082\,
            I => \N__42047\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__42077\,
            I => \N__42047\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__42060\,
            I => \N__42047\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__42057\,
            I => \foc.u_Park_Transform.n598\
        );

    \I__6908\ : Odrv12
    port map (
            O => \N__42054\,
            I => \foc.u_Park_Transform.n598\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__42047\,
            I => \foc.u_Park_Transform.n598\
        );

    \I__6906\ : InMux
    port map (
            O => \N__42040\,
            I => \N__42037\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__42037\,
            I => \N__42034\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__42034\,
            I => \foc.u_Park_Transform.n57\
        );

    \I__6903\ : InMux
    port map (
            O => \N__42031\,
            I => \N__42028\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__42028\,
            I => \foc.u_Park_Transform.n60\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__42025\,
            I => \N__42022\
        );

    \I__6900\ : InMux
    port map (
            O => \N__42022\,
            I => \N__42019\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__42019\,
            I => \N__42016\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__42016\,
            I => \N__42013\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__42013\,
            I => \foc.u_Park_Transform.n106\
        );

    \I__6896\ : InMux
    port map (
            O => \N__42010\,
            I => \foc.u_Park_Transform.n17038\
        );

    \I__6895\ : CascadeMux
    port map (
            O => \N__42007\,
            I => \N__42004\
        );

    \I__6894\ : InMux
    port map (
            O => \N__42004\,
            I => \N__42001\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__42001\,
            I => \foc.u_Park_Transform.n109\
        );

    \I__6892\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41995\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__41995\,
            I => \N__41992\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__41992\,
            I => \foc.u_Park_Transform.n155\
        );

    \I__6889\ : InMux
    port map (
            O => \N__41989\,
            I => \foc.u_Park_Transform.n17039\
        );

    \I__6888\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41983\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__41983\,
            I => \foc.u_Park_Transform.n158\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__41980\,
            I => \N__41977\
        );

    \I__6885\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41974\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__41974\,
            I => \N__41971\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__41971\,
            I => \foc.u_Park_Transform.n204\
        );

    \I__6882\ : InMux
    port map (
            O => \N__41968\,
            I => \foc.u_Park_Transform.n17040\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__41965\,
            I => \N__41962\
        );

    \I__6880\ : InMux
    port map (
            O => \N__41962\,
            I => \N__41959\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__41959\,
            I => \foc.u_Park_Transform.n207\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__41956\,
            I => \N__41953\
        );

    \I__6877\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41950\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__41950\,
            I => \N__41947\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__41947\,
            I => \foc.u_Park_Transform.n253\
        );

    \I__6874\ : InMux
    port map (
            O => \N__41944\,
            I => \foc.u_Park_Transform.n17041\
        );

    \I__6873\ : InMux
    port map (
            O => \N__41941\,
            I => \N__41938\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__41938\,
            I => \foc.u_Park_Transform.n256\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__41935\,
            I => \N__41932\
        );

    \I__6870\ : InMux
    port map (
            O => \N__41932\,
            I => \N__41929\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__41929\,
            I => \N__41926\
        );

    \I__6868\ : Span4Mux_h
    port map (
            O => \N__41926\,
            I => \N__41923\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__41923\,
            I => \foc.u_Park_Transform.n302\
        );

    \I__6866\ : InMux
    port map (
            O => \N__41920\,
            I => \foc.u_Park_Transform.n17042\
        );

    \I__6865\ : InMux
    port map (
            O => \N__41917\,
            I => \N__41914\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__41914\,
            I => \N__41911\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__41911\,
            I => \foc.u_Park_Transform.n354_adj_2133\
        );

    \I__6862\ : InMux
    port map (
            O => \N__41908\,
            I => \foc.u_Park_Transform.n17211\
        );

    \I__6861\ : InMux
    port map (
            O => \N__41905\,
            I => \N__41902\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__41902\,
            I => \N__41899\
        );

    \I__6859\ : Odrv12
    port map (
            O => \N__41899\,
            I => \foc.u_Park_Transform.n357_adj_2151\
        );

    \I__6858\ : CascadeMux
    port map (
            O => \N__41896\,
            I => \N__41893\
        );

    \I__6857\ : InMux
    port map (
            O => \N__41893\,
            I => \N__41890\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__41890\,
            I => \N__41887\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__41887\,
            I => \N__41884\
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__41884\,
            I => \foc.u_Park_Transform.n403_adj_2132\
        );

    \I__6853\ : InMux
    port map (
            O => \N__41881\,
            I => \foc.u_Park_Transform.n17212\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__41878\,
            I => \N__41875\
        );

    \I__6851\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41872\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__41872\,
            I => \N__41869\
        );

    \I__6849\ : Span4Mux_h
    port map (
            O => \N__41869\,
            I => \N__41866\
        );

    \I__6848\ : Odrv4
    port map (
            O => \N__41866\,
            I => \foc.u_Park_Transform.n406_adj_2150\
        );

    \I__6847\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41860\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__41860\,
            I => \N__41857\
        );

    \I__6845\ : Odrv4
    port map (
            O => \N__41857\,
            I => \foc.u_Park_Transform.n452_adj_2131\
        );

    \I__6844\ : InMux
    port map (
            O => \N__41854\,
            I => \bfn_16_12_0_\
        );

    \I__6843\ : InMux
    port map (
            O => \N__41851\,
            I => \N__41848\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__41848\,
            I => \N__41845\
        );

    \I__6841\ : Odrv12
    port map (
            O => \N__41845\,
            I => \foc.u_Park_Transform.n455_adj_2148\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__41842\,
            I => \N__41839\
        );

    \I__6839\ : InMux
    port map (
            O => \N__41839\,
            I => \N__41836\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__41836\,
            I => \N__41833\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__41833\,
            I => \foc.u_Park_Transform.n501_adj_2130\
        );

    \I__6836\ : InMux
    port map (
            O => \N__41830\,
            I => \foc.u_Park_Transform.n17214\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__41827\,
            I => \N__41824\
        );

    \I__6834\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41821\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__41821\,
            I => \N__41818\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__41818\,
            I => \foc.u_Park_Transform.n504_adj_2147\
        );

    \I__6831\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41812\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__41812\,
            I => \N__41809\
        );

    \I__6829\ : Span4Mux_h
    port map (
            O => \N__41809\,
            I => \N__41806\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__41806\,
            I => \foc.u_Park_Transform.n550_adj_2129\
        );

    \I__6827\ : InMux
    port map (
            O => \N__41803\,
            I => \foc.u_Park_Transform.n17215\
        );

    \I__6826\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41797\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__41797\,
            I => \N__41794\
        );

    \I__6824\ : Odrv12
    port map (
            O => \N__41794\,
            I => \foc.u_Park_Transform.n553_adj_2146\
        );

    \I__6823\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41788\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__41788\,
            I => \N__41785\
        );

    \I__6821\ : Odrv12
    port map (
            O => \N__41785\,
            I => \foc.u_Park_Transform.n599_adj_2128\
        );

    \I__6820\ : InMux
    port map (
            O => \N__41782\,
            I => \foc.u_Park_Transform.n17216\
        );

    \I__6819\ : InMux
    port map (
            O => \N__41779\,
            I => \N__41776\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__41776\,
            I => \N__41773\
        );

    \I__6817\ : Odrv12
    port map (
            O => \N__41773\,
            I => \foc.u_Park_Transform.n602_adj_2144\
        );

    \I__6816\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41767\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__41767\,
            I => \N__41764\
        );

    \I__6814\ : Odrv12
    port map (
            O => \N__41764\,
            I => \foc.u_Park_Transform.n648_adj_2124\
        );

    \I__6813\ : InMux
    port map (
            O => \N__41761\,
            I => \foc.u_Park_Transform.n17217\
        );

    \I__6812\ : InMux
    port map (
            O => \N__41758\,
            I => \N__41755\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__41755\,
            I => \N__41752\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__41752\,
            I => \foc.u_Park_Transform.n651_adj_2143\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__41749\,
            I => \N__41746\
        );

    \I__6808\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41743\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__41743\,
            I => \N__41740\
        );

    \I__6806\ : Odrv12
    port map (
            O => \N__41740\,
            I => \foc.u_Park_Transform.n697_adj_2121\
        );

    \I__6805\ : InMux
    port map (
            O => \N__41737\,
            I => \foc.u_Park_Transform.n17218\
        );

    \I__6804\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41731\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__41731\,
            I => \N__41728\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__41728\,
            I => \N__41725\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__41725\,
            I => \foc.dCurrent_27\
        );

    \I__6800\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41719\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__41719\,
            I => \N__41716\
        );

    \I__6798\ : Sp12to4
    port map (
            O => \N__41716\,
            I => \N__41713\
        );

    \I__6797\ : Odrv12
    port map (
            O => \N__41713\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n6\
        );

    \I__6796\ : InMux
    port map (
            O => \N__41710\,
            I => \N__41704\
        );

    \I__6795\ : CascadeMux
    port map (
            O => \N__41709\,
            I => \N__41701\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__41708\,
            I => \N__41697\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__41707\,
            I => \N__41693\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__41704\,
            I => \N__41682\
        );

    \I__6791\ : InMux
    port map (
            O => \N__41701\,
            I => \N__41669\
        );

    \I__6790\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41669\
        );

    \I__6789\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41669\
        );

    \I__6788\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41669\
        );

    \I__6787\ : InMux
    port map (
            O => \N__41693\,
            I => \N__41669\
        );

    \I__6786\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41669\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__41691\,
            I => \N__41663\
        );

    \I__6784\ : CascadeMux
    port map (
            O => \N__41690\,
            I => \N__41657\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__41689\,
            I => \N__41654\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__41688\,
            I => \N__41648\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__41687\,
            I => \N__41644\
        );

    \I__6780\ : CascadeMux
    port map (
            O => \N__41686\,
            I => \N__41640\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__41685\,
            I => \N__41635\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__41682\,
            I => \N__41630\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__41669\,
            I => \N__41630\
        );

    \I__6776\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41621\
        );

    \I__6775\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41621\
        );

    \I__6774\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41621\
        );

    \I__6773\ : InMux
    port map (
            O => \N__41663\,
            I => \N__41621\
        );

    \I__6772\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41612\
        );

    \I__6771\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41612\
        );

    \I__6770\ : InMux
    port map (
            O => \N__41660\,
            I => \N__41612\
        );

    \I__6769\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41612\
        );

    \I__6768\ : InMux
    port map (
            O => \N__41654\,
            I => \N__41609\
        );

    \I__6767\ : CascadeMux
    port map (
            O => \N__41653\,
            I => \N__41605\
        );

    \I__6766\ : CascadeMux
    port map (
            O => \N__41652\,
            I => \N__41601\
        );

    \I__6765\ : CascadeMux
    port map (
            O => \N__41651\,
            I => \N__41597\
        );

    \I__6764\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41584\
        );

    \I__6763\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41584\
        );

    \I__6762\ : InMux
    port map (
            O => \N__41644\,
            I => \N__41584\
        );

    \I__6761\ : InMux
    port map (
            O => \N__41643\,
            I => \N__41584\
        );

    \I__6760\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41584\
        );

    \I__6759\ : InMux
    port map (
            O => \N__41639\,
            I => \N__41584\
        );

    \I__6758\ : InMux
    port map (
            O => \N__41638\,
            I => \N__41579\
        );

    \I__6757\ : InMux
    port map (
            O => \N__41635\,
            I => \N__41579\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__41630\,
            I => \N__41572\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__41621\,
            I => \N__41572\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__41612\,
            I => \N__41572\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__41609\,
            I => \N__41569\
        );

    \I__6752\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41556\
        );

    \I__6751\ : InMux
    port map (
            O => \N__41605\,
            I => \N__41556\
        );

    \I__6750\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41556\
        );

    \I__6749\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41556\
        );

    \I__6748\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41556\
        );

    \I__6747\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41556\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__41584\,
            I => \N__41551\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41551\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__41572\,
            I => \foc.u_Park_Transform.n601\
        );

    \I__6743\ : Odrv12
    port map (
            O => \N__41569\,
            I => \foc.u_Park_Transform.n601\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__41556\,
            I => \foc.u_Park_Transform.n601\
        );

    \I__6741\ : Odrv4
    port map (
            O => \N__41551\,
            I => \foc.u_Park_Transform.n601\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__41542\,
            I => \N__41539\
        );

    \I__6739\ : InMux
    port map (
            O => \N__41539\,
            I => \N__41536\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__41536\,
            I => \N__41533\
        );

    \I__6737\ : Odrv4
    port map (
            O => \N__41533\,
            I => \foc.u_Park_Transform.n60_adj_2140\
        );

    \I__6736\ : InMux
    port map (
            O => \N__41530\,
            I => \N__41527\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__41527\,
            I => \N__41524\
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__41524\,
            I => \foc.u_Park_Transform.n63_adj_2158\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__41521\,
            I => \N__41518\
        );

    \I__6732\ : InMux
    port map (
            O => \N__41518\,
            I => \N__41515\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__41515\,
            I => \N__41512\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__41512\,
            I => \foc.u_Park_Transform.n109_adj_2139\
        );

    \I__6729\ : InMux
    port map (
            O => \N__41509\,
            I => \foc.u_Park_Transform.n17206\
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__41506\,
            I => \N__41503\
        );

    \I__6727\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41500\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41497\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__41497\,
            I => \foc.u_Park_Transform.n112_adj_2157\
        );

    \I__6724\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41491\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__41491\,
            I => \N__41488\
        );

    \I__6722\ : Odrv12
    port map (
            O => \N__41488\,
            I => \foc.u_Park_Transform.n158_adj_2137\
        );

    \I__6721\ : InMux
    port map (
            O => \N__41485\,
            I => \foc.u_Park_Transform.n17207\
        );

    \I__6720\ : InMux
    port map (
            O => \N__41482\,
            I => \N__41479\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__41479\,
            I => \N__41476\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__41476\,
            I => \foc.u_Park_Transform.n161_adj_2156\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__41473\,
            I => \N__41470\
        );

    \I__6716\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41467\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__41467\,
            I => \N__41464\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__41464\,
            I => \foc.u_Park_Transform.n207_adj_2136\
        );

    \I__6713\ : InMux
    port map (
            O => \N__41461\,
            I => \foc.u_Park_Transform.n17208\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__41458\,
            I => \N__41455\
        );

    \I__6711\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41452\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__41452\,
            I => \N__41449\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__41449\,
            I => \foc.u_Park_Transform.n210_adj_2155\
        );

    \I__6708\ : InMux
    port map (
            O => \N__41446\,
            I => \N__41443\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__41443\,
            I => \N__41440\
        );

    \I__6706\ : Span4Mux_h
    port map (
            O => \N__41440\,
            I => \N__41437\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__41437\,
            I => \foc.u_Park_Transform.n256_adj_2135\
        );

    \I__6704\ : InMux
    port map (
            O => \N__41434\,
            I => \foc.u_Park_Transform.n17209\
        );

    \I__6703\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41428\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__41428\,
            I => \N__41425\
        );

    \I__6701\ : Odrv12
    port map (
            O => \N__41425\,
            I => \foc.u_Park_Transform.n259_adj_2154\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__41422\,
            I => \N__41419\
        );

    \I__6699\ : InMux
    port map (
            O => \N__41419\,
            I => \N__41416\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__41416\,
            I => \N__41413\
        );

    \I__6697\ : Span4Mux_v
    port map (
            O => \N__41413\,
            I => \N__41410\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__41410\,
            I => \foc.u_Park_Transform.n305_adj_2134\
        );

    \I__6695\ : InMux
    port map (
            O => \N__41407\,
            I => \foc.u_Park_Transform.n17210\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__41404\,
            I => \N__41401\
        );

    \I__6693\ : InMux
    port map (
            O => \N__41401\,
            I => \N__41398\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__41398\,
            I => \N__41395\
        );

    \I__6691\ : Odrv12
    port map (
            O => \N__41395\,
            I => \foc.u_Park_Transform.n308_adj_2153\
        );

    \I__6690\ : InMux
    port map (
            O => \N__41392\,
            I => \N__41388\
        );

    \I__6689\ : InMux
    port map (
            O => \N__41391\,
            I => \N__41385\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__41388\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__41385\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18\
        );

    \I__6686\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41374\
        );

    \I__6685\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41374\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__41374\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_25\
        );

    \I__6683\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41368\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__41368\,
            I => \N__41364\
        );

    \I__6681\ : InMux
    port map (
            O => \N__41367\,
            I => \N__41361\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__41364\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__41361\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17\
        );

    \I__6678\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41350\
        );

    \I__6677\ : InMux
    port map (
            O => \N__41355\,
            I => \N__41350\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__41350\,
            I => \N__41347\
        );

    \I__6675\ : Odrv4
    port map (
            O => \N__41347\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_24\
        );

    \I__6674\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41341\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41338\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__41338\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n611_adj_623\
        );

    \I__6671\ : InMux
    port map (
            O => \N__41335\,
            I => \N__41332\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__41332\,
            I => \N__41329\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__41329\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n657_adj_638\
        );

    \I__6668\ : InMux
    port map (
            O => \N__41326\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18088\
        );

    \I__6667\ : CascadeMux
    port map (
            O => \N__41323\,
            I => \N__41320\
        );

    \I__6666\ : InMux
    port map (
            O => \N__41320\,
            I => \N__41317\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__41317\,
            I => \N__41314\
        );

    \I__6664\ : Odrv12
    port map (
            O => \N__41314\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n660_adj_622\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__41311\,
            I => \N__41308\
        );

    \I__6662\ : InMux
    port map (
            O => \N__41308\,
            I => \N__41305\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__41305\,
            I => \N__41302\
        );

    \I__6660\ : Odrv4
    port map (
            O => \N__41302\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n706_adj_637\
        );

    \I__6659\ : InMux
    port map (
            O => \N__41299\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18089\
        );

    \I__6658\ : CascadeMux
    port map (
            O => \N__41296\,
            I => \N__41293\
        );

    \I__6657\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41290\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__41290\,
            I => \N__41287\
        );

    \I__6655\ : Odrv12
    port map (
            O => \N__41287\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n709_adj_621\
        );

    \I__6654\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41281\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41278\
        );

    \I__6652\ : Span12Mux_v
    port map (
            O => \N__41278\,
            I => \N__41275\
        );

    \I__6651\ : Odrv12
    port map (
            O => \N__41275\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n762_adj_635\
        );

    \I__6650\ : InMux
    port map (
            O => \N__41272\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18090\
        );

    \I__6649\ : InMux
    port map (
            O => \N__41269\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636\
        );

    \I__6648\ : CascadeMux
    port map (
            O => \N__41266\,
            I => \N__41263\
        );

    \I__6647\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41260\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__41260\,
            I => \N__41257\
        );

    \I__6645\ : Span4Mux_h
    port map (
            O => \N__41257\,
            I => \N__41254\
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__41254\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_CO\
        );

    \I__6643\ : InMux
    port map (
            O => \N__41251\,
            I => \N__41245\
        );

    \I__6642\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41245\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__41245\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_16\
        );

    \I__6640\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41238\
        );

    \I__6639\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41235\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__41238\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__41235\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20\
        );

    \I__6636\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41227\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__6634\ : Odrv12
    port map (
            O => \N__41224\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n219_adj_631\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__41221\,
            I => \N__41218\
        );

    \I__6632\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41215\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__41215\,
            I => \N__41212\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__41212\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n265_adj_646\
        );

    \I__6629\ : InMux
    port map (
            O => \N__41209\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18080\
        );

    \I__6628\ : CascadeMux
    port map (
            O => \N__41206\,
            I => \N__41203\
        );

    \I__6627\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41200\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__41200\,
            I => \N__41197\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__41197\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n268_adj_630\
        );

    \I__6624\ : InMux
    port map (
            O => \N__41194\,
            I => \N__41191\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__41191\,
            I => \N__41188\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__41188\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n314_adj_645\
        );

    \I__6621\ : InMux
    port map (
            O => \N__41185\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18081\
        );

    \I__6620\ : CascadeMux
    port map (
            O => \N__41182\,
            I => \N__41179\
        );

    \I__6619\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41176\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__41176\,
            I => \N__41173\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__41173\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n317_adj_629\
        );

    \I__6616\ : CascadeMux
    port map (
            O => \N__41170\,
            I => \N__41167\
        );

    \I__6615\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41164\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__41164\,
            I => \N__41161\
        );

    \I__6613\ : Odrv4
    port map (
            O => \N__41161\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n363_adj_644\
        );

    \I__6612\ : InMux
    port map (
            O => \N__41158\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18082\
        );

    \I__6611\ : InMux
    port map (
            O => \N__41155\,
            I => \N__41152\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__41152\,
            I => \N__41149\
        );

    \I__6609\ : Odrv12
    port map (
            O => \N__41149\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n366_adj_628\
        );

    \I__6608\ : InMux
    port map (
            O => \N__41146\,
            I => \N__41143\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__41143\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n412_adj_643\
        );

    \I__6606\ : InMux
    port map (
            O => \N__41140\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18083\
        );

    \I__6605\ : InMux
    port map (
            O => \N__41137\,
            I => \N__41134\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__41134\,
            I => \N__41131\
        );

    \I__6603\ : Span4Mux_v
    port map (
            O => \N__41131\,
            I => \N__41128\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__41128\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n415_adj_627\
        );

    \I__6601\ : CascadeMux
    port map (
            O => \N__41125\,
            I => \N__41122\
        );

    \I__6600\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41119\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__41119\,
            I => \N__41116\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__41116\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n461_adj_642\
        );

    \I__6597\ : InMux
    port map (
            O => \N__41113\,
            I => \bfn_15_26_0_\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__41110\,
            I => \N__41107\
        );

    \I__6595\ : InMux
    port map (
            O => \N__41107\,
            I => \N__41104\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__41101\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n464_adj_626\
        );

    \I__6592\ : InMux
    port map (
            O => \N__41098\,
            I => \N__41095\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__41095\,
            I => \N__41092\
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__41092\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n510_adj_641\
        );

    \I__6589\ : InMux
    port map (
            O => \N__41089\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18085\
        );

    \I__6588\ : InMux
    port map (
            O => \N__41086\,
            I => \N__41083\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__41083\,
            I => \N__41080\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__41080\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n513_adj_625\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__41077\,
            I => \N__41074\
        );

    \I__6584\ : InMux
    port map (
            O => \N__41074\,
            I => \N__41071\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__41071\,
            I => \N__41068\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__41068\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n559_adj_640\
        );

    \I__6581\ : InMux
    port map (
            O => \N__41065\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18086\
        );

    \I__6580\ : CascadeMux
    port map (
            O => \N__41062\,
            I => \N__41059\
        );

    \I__6579\ : InMux
    port map (
            O => \N__41059\,
            I => \N__41056\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41053\
        );

    \I__6577\ : Odrv12
    port map (
            O => \N__41053\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n562_adj_624\
        );

    \I__6576\ : InMux
    port map (
            O => \N__41050\,
            I => \N__41047\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__41047\,
            I => \N__41044\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__41044\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n608_adj_639\
        );

    \I__6573\ : InMux
    port map (
            O => \N__41041\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18087\
        );

    \I__6572\ : InMux
    port map (
            O => \N__41038\,
            I => \N__41035\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__41035\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n654_adj_654\
        );

    \I__6570\ : InMux
    port map (
            O => \N__41032\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18073\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__41029\,
            I => \N__41026\
        );

    \I__6568\ : InMux
    port map (
            O => \N__41026\,
            I => \N__41023\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__41023\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n703_adj_653\
        );

    \I__6566\ : InMux
    port map (
            O => \N__41020\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18074\
        );

    \I__6565\ : InMux
    port map (
            O => \N__41017\,
            I => \N__41014\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__41014\,
            I => \N__41011\
        );

    \I__6563\ : Span4Mux_v
    port map (
            O => \N__41011\,
            I => \N__41008\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__41008\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n758_adj_651\
        );

    \I__6561\ : InMux
    port map (
            O => \N__41005\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18075\
        );

    \I__6560\ : InMux
    port map (
            O => \N__41002\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__40999\,
            I => \N__40996\
        );

    \I__6558\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40993\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__40993\,
            I => \N__40990\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__40990\,
            I => \N__40987\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__40987\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_CO\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__40984\,
            I => \N__40981\
        );

    \I__6553\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40978\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__40978\,
            I => \N__40975\
        );

    \I__6551\ : Odrv12
    port map (
            O => \N__40975\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n69_adj_650\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__40972\,
            I => \N__40969\
        );

    \I__6549\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40966\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__40966\,
            I => \N__40963\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__40963\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n72_adj_634\
        );

    \I__6546\ : InMux
    port map (
            O => \N__40960\,
            I => \N__40957\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__40957\,
            I => \N__40954\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__40954\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n118_adj_649\
        );

    \I__6543\ : InMux
    port map (
            O => \N__40951\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18077\
        );

    \I__6542\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40945\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__40945\,
            I => \N__40942\
        );

    \I__6540\ : Odrv12
    port map (
            O => \N__40942\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n121_adj_633\
        );

    \I__6539\ : CascadeMux
    port map (
            O => \N__40939\,
            I => \N__40936\
        );

    \I__6538\ : InMux
    port map (
            O => \N__40936\,
            I => \N__40933\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__40933\,
            I => \N__40930\
        );

    \I__6536\ : Odrv12
    port map (
            O => \N__40930\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n167_adj_648\
        );

    \I__6535\ : InMux
    port map (
            O => \N__40927\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18078\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__40924\,
            I => \N__40921\
        );

    \I__6533\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40918\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40915\
        );

    \I__6531\ : Odrv12
    port map (
            O => \N__40915\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n170_adj_632\
        );

    \I__6530\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40909\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__40909\,
            I => \N__40906\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__40906\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n216_adj_647\
        );

    \I__6527\ : InMux
    port map (
            O => \N__40903\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18079\
        );

    \I__6526\ : InMux
    port map (
            O => \N__40900\,
            I => \N__40897\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__40897\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n262_adj_662\
        );

    \I__6524\ : InMux
    port map (
            O => \N__40894\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18065\
        );

    \I__6523\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40888\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__40888\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n311_adj_661\
        );

    \I__6521\ : InMux
    port map (
            O => \N__40885\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18066\
        );

    \I__6520\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40879\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__40879\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n360_adj_660\
        );

    \I__6518\ : InMux
    port map (
            O => \N__40876\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18067\
        );

    \I__6517\ : InMux
    port map (
            O => \N__40873\,
            I => \N__40870\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__40870\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n409_adj_659\
        );

    \I__6515\ : InMux
    port map (
            O => \N__40867\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18068\
        );

    \I__6514\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40861\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__40861\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n458_adj_658\
        );

    \I__6512\ : InMux
    port map (
            O => \N__40858\,
            I => \bfn_15_24_0_\
        );

    \I__6511\ : InMux
    port map (
            O => \N__40855\,
            I => \N__40852\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__40852\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n507_adj_657\
        );

    \I__6509\ : InMux
    port map (
            O => \N__40849\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18070\
        );

    \I__6508\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40843\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__40843\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n556_adj_656\
        );

    \I__6506\ : InMux
    port map (
            O => \N__40840\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18071\
        );

    \I__6505\ : InMux
    port map (
            O => \N__40837\,
            I => \N__40834\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__40834\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n605_adj_655\
        );

    \I__6503\ : InMux
    port map (
            O => \N__40831\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18072\
        );

    \I__6502\ : InMux
    port map (
            O => \N__40828\,
            I => \N__40825\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__40825\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n90_adj_729\
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__40822\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n7_adj_760_cascade_\
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__40819\,
            I => \N__40816\
        );

    \I__6498\ : InMux
    port map (
            O => \N__40816\,
            I => \N__40813\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__40813\,
            I => \N__40810\
        );

    \I__6496\ : Span4Mux_v
    port map (
            O => \N__40810\,
            I => \N__40807\
        );

    \I__6495\ : Odrv4
    port map (
            O => \N__40807\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_adj_732\
        );

    \I__6494\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40795\
        );

    \I__6493\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40795\
        );

    \I__6492\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40795\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__40795\,
            I => \N__40792\
        );

    \I__6490\ : Odrv4
    port map (
            O => \N__40792\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n26_adj_759\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__40789\,
            I => \N__40786\
        );

    \I__6488\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40783\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__40783\,
            I => \N__40780\
        );

    \I__6486\ : Span4Mux_v
    port map (
            O => \N__40780\,
            I => \N__40777\
        );

    \I__6485\ : Odrv4
    port map (
            O => \N__40777\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n790_adj_733\
        );

    \I__6484\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40771\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__40771\,
            I => \N__40768\
        );

    \I__6482\ : Span4Mux_h
    port map (
            O => \N__40768\,
            I => \N__40765\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__40765\,
            I => n794_adj_2425
        );

    \I__6480\ : InMux
    port map (
            O => \N__40762\,
            I => \N__40759\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__40759\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n66_adj_666\
        );

    \I__6478\ : InMux
    port map (
            O => \N__40756\,
            I => \N__40753\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__40753\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n115_adj_665\
        );

    \I__6476\ : InMux
    port map (
            O => \N__40750\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18062\
        );

    \I__6475\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40744\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__40744\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n164_adj_664\
        );

    \I__6473\ : InMux
    port map (
            O => \N__40741\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18063\
        );

    \I__6472\ : InMux
    port map (
            O => \N__40738\,
            I => \N__40735\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__40735\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n213_adj_663\
        );

    \I__6470\ : InMux
    port map (
            O => \N__40732\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18064\
        );

    \I__6469\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40726\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__40726\,
            I => \foc.qCurrent_25\
        );

    \I__6467\ : InMux
    port map (
            O => \N__40723\,
            I => \N__40720\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__40720\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n87_adj_730\
        );

    \I__6465\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40714\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__40714\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n136_adj_728\
        );

    \I__6463\ : InMux
    port map (
            O => \N__40711\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17973\
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__40708\,
            I => \N__40705\
        );

    \I__6461\ : InMux
    port map (
            O => \N__40705\,
            I => \N__40702\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__40702\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n185_adj_726\
        );

    \I__6459\ : InMux
    port map (
            O => \N__40699\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17974\
        );

    \I__6458\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40693\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__40693\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n234_adj_724\
        );

    \I__6456\ : InMux
    port map (
            O => \N__40690\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17975\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__40687\,
            I => \N__40684\
        );

    \I__6454\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40681\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__40681\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n283_adj_723\
        );

    \I__6452\ : InMux
    port map (
            O => \N__40678\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17976\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__40675\,
            I => \N__40671\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__40674\,
            I => \N__40667\
        );

    \I__6449\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40664\
        );

    \I__6448\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40659\
        );

    \I__6447\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40659\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__40664\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__40659\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722\
        );

    \I__6444\ : InMux
    port map (
            O => \N__40654\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17977\
        );

    \I__6443\ : InMux
    port map (
            O => \N__40651\,
            I => \N__40648\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__40648\,
            I => \N__40645\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__40645\,
            I => \N__40642\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__40642\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n786_adj_719\
        );

    \I__6439\ : InMux
    port map (
            O => \N__40639\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17978\
        );

    \I__6438\ : InMux
    port map (
            O => \N__40636\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721\
        );

    \I__6437\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40630\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__40630\,
            I => \N__40627\
        );

    \I__6435\ : Span4Mux_h
    port map (
            O => \N__40627\,
            I => \N__40624\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__40624\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_CO\
        );

    \I__6433\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40618\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__40618\,
            I => \foc.qCurrent_26\
        );

    \I__6431\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40612\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__40612\,
            I => \foc.qCurrent_12\
        );

    \I__6429\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40606\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__40606\,
            I => \foc.qCurrent_28\
        );

    \I__6427\ : InMux
    port map (
            O => \N__40603\,
            I => \N__40600\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__40600\,
            I => \foc.qCurrent_20\
        );

    \I__6425\ : CascadeMux
    port map (
            O => \N__40597\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_757_cascade_\
        );

    \I__6424\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40591\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__40591\,
            I => \N__40588\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__40588\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_758\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__40585\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19841_cascade_\
        );

    \I__6420\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40579\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__40579\,
            I => \foc.qCurrent_31\
        );

    \I__6418\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__40573\,
            I => \foc.qCurrent_16\
        );

    \I__6416\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40567\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__40567\,
            I => \foc.qCurrent_14\
        );

    \I__6414\ : InMux
    port map (
            O => \N__40564\,
            I => \N__40561\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__40561\,
            I => \foc.qCurrent_4\
        );

    \I__6412\ : InMux
    port map (
            O => \N__40558\,
            I => \N__40555\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__40555\,
            I => \foc.qCurrent_11\
        );

    \I__6410\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40549\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__40549\,
            I => \foc.qCurrent_15\
        );

    \I__6408\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40543\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__40543\,
            I => \foc.qCurrent_22\
        );

    \I__6406\ : InMux
    port map (
            O => \N__40540\,
            I => \N__40537\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__40537\,
            I => \foc.qCurrent_17\
        );

    \I__6404\ : InMux
    port map (
            O => \N__40534\,
            I => \N__40531\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__40531\,
            I => \foc.qCurrent_24\
        );

    \I__6402\ : InMux
    port map (
            O => \N__40528\,
            I => \N__40525\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__40525\,
            I => \foc.qCurrent_27\
        );

    \I__6400\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40519\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__40519\,
            I => \foc.qCurrent_6\
        );

    \I__6398\ : InMux
    port map (
            O => \N__40516\,
            I => \N__40513\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__40513\,
            I => \N__40509\
        );

    \I__6396\ : InMux
    port map (
            O => \N__40512\,
            I => \N__40506\
        );

    \I__6395\ : Odrv12
    port map (
            O => \N__40509\,
            I => \foc.u_Park_Transform.n741\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__40506\,
            I => \foc.u_Park_Transform.n741\
        );

    \I__6393\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40498\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__40498\,
            I => \N__40494\
        );

    \I__6391\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40491\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__40494\,
            I => \N__40486\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__40491\,
            I => \N__40486\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__40486\,
            I => \N__40481\
        );

    \I__6387\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40476\
        );

    \I__6386\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40476\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__40481\,
            I => \N__40470\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__40476\,
            I => \N__40470\
        );

    \I__6383\ : InMux
    port map (
            O => \N__40475\,
            I => \N__40467\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__40470\,
            I => \Look_Up_Table_out1_1_14\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__40467\,
            I => \Look_Up_Table_out1_1_14\
        );

    \I__6380\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40459\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__40459\,
            I => \N__40454\
        );

    \I__6378\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40451\
        );

    \I__6377\ : InMux
    port map (
            O => \N__40457\,
            I => \N__40448\
        );

    \I__6376\ : Span4Mux_v
    port map (
            O => \N__40454\,
            I => \N__40443\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__40451\,
            I => \N__40440\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__40448\,
            I => \N__40437\
        );

    \I__6373\ : InMux
    port map (
            O => \N__40447\,
            I => \N__40434\
        );

    \I__6372\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40431\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__40443\,
            I => \N__40426\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__40440\,
            I => \N__40426\
        );

    \I__6369\ : Span4Mux_h
    port map (
            O => \N__40437\,
            I => \N__40421\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__40434\,
            I => \N__40421\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__40431\,
            I => \N__40418\
        );

    \I__6366\ : Odrv4
    port map (
            O => \N__40426\,
            I => \Look_Up_Table_out1_1_15\
        );

    \I__6365\ : Odrv4
    port map (
            O => \N__40421\,
            I => \Look_Up_Table_out1_1_15\
        );

    \I__6364\ : Odrv12
    port map (
            O => \N__40418\,
            I => \Look_Up_Table_out1_1_15\
        );

    \I__6363\ : InMux
    port map (
            O => \N__40411\,
            I => \N__40408\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__40408\,
            I => \foc.qCurrent_8\
        );

    \I__6361\ : InMux
    port map (
            O => \N__40405\,
            I => \N__40399\
        );

    \I__6360\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40399\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__40399\,
            I => \N__40396\
        );

    \I__6358\ : Span4Mux_v
    port map (
            O => \N__40396\,
            I => \N__40393\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__40393\,
            I => \foc.Look_Up_Table_out1_1_1\
        );

    \I__6356\ : InMux
    port map (
            O => \N__40390\,
            I => \N__40380\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__40389\,
            I => \N__40377\
        );

    \I__6354\ : CascadeMux
    port map (
            O => \N__40388\,
            I => \N__40373\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__40387\,
            I => \N__40369\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__40386\,
            I => \N__40364\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__40385\,
            I => \N__40361\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__40384\,
            I => \N__40357\
        );

    \I__6349\ : CascadeMux
    port map (
            O => \N__40383\,
            I => \N__40353\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__40380\,
            I => \N__40345\
        );

    \I__6347\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40332\
        );

    \I__6346\ : InMux
    port map (
            O => \N__40376\,
            I => \N__40332\
        );

    \I__6345\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40332\
        );

    \I__6344\ : InMux
    port map (
            O => \N__40372\,
            I => \N__40332\
        );

    \I__6343\ : InMux
    port map (
            O => \N__40369\,
            I => \N__40332\
        );

    \I__6342\ : InMux
    port map (
            O => \N__40368\,
            I => \N__40332\
        );

    \I__6341\ : InMux
    port map (
            O => \N__40367\,
            I => \N__40327\
        );

    \I__6340\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40327\
        );

    \I__6339\ : InMux
    port map (
            O => \N__40361\,
            I => \N__40314\
        );

    \I__6338\ : InMux
    port map (
            O => \N__40360\,
            I => \N__40314\
        );

    \I__6337\ : InMux
    port map (
            O => \N__40357\,
            I => \N__40314\
        );

    \I__6336\ : InMux
    port map (
            O => \N__40356\,
            I => \N__40314\
        );

    \I__6335\ : InMux
    port map (
            O => \N__40353\,
            I => \N__40314\
        );

    \I__6334\ : InMux
    port map (
            O => \N__40352\,
            I => \N__40314\
        );

    \I__6333\ : CascadeMux
    port map (
            O => \N__40351\,
            I => \N__40308\
        );

    \I__6332\ : CascadeMux
    port map (
            O => \N__40350\,
            I => \N__40304\
        );

    \I__6331\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40296\
        );

    \I__6330\ : InMux
    port map (
            O => \N__40348\,
            I => \N__40296\
        );

    \I__6329\ : Span4Mux_v
    port map (
            O => \N__40345\,
            I => \N__40287\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40287\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__40327\,
            I => \N__40287\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__40314\,
            I => \N__40287\
        );

    \I__6325\ : InMux
    port map (
            O => \N__40313\,
            I => \N__40284\
        );

    \I__6324\ : InMux
    port map (
            O => \N__40312\,
            I => \N__40271\
        );

    \I__6323\ : InMux
    port map (
            O => \N__40311\,
            I => \N__40271\
        );

    \I__6322\ : InMux
    port map (
            O => \N__40308\,
            I => \N__40271\
        );

    \I__6321\ : InMux
    port map (
            O => \N__40307\,
            I => \N__40271\
        );

    \I__6320\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40271\
        );

    \I__6319\ : InMux
    port map (
            O => \N__40303\,
            I => \N__40271\
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__40302\,
            I => \N__40266\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__40301\,
            I => \N__40262\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__40296\,
            I => \N__40258\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__40287\,
            I => \N__40251\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__40284\,
            I => \N__40251\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__40271\,
            I => \N__40251\
        );

    \I__6312\ : InMux
    port map (
            O => \N__40270\,
            I => \N__40248\
        );

    \I__6311\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40237\
        );

    \I__6310\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40237\
        );

    \I__6309\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40237\
        );

    \I__6308\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40237\
        );

    \I__6307\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40237\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__40258\,
            I => \foc.u_Park_Transform.n592\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__40251\,
            I => \foc.u_Park_Transform.n592\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__40248\,
            I => \foc.u_Park_Transform.n592\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__40237\,
            I => \foc.u_Park_Transform.n592\
        );

    \I__6302\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40225\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__40225\,
            I => \N__40222\
        );

    \I__6300\ : Odrv4
    port map (
            O => \N__40222\,
            I => \foc.qCurrent_3\
        );

    \I__6299\ : InMux
    port map (
            O => \N__40219\,
            I => \N__40216\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__40216\,
            I => \foc.qCurrent_18\
        );

    \I__6297\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__40210\,
            I => \foc.qCurrent_19\
        );

    \I__6295\ : InMux
    port map (
            O => \N__40207\,
            I => \N__40204\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__40204\,
            I => \foc.qCurrent_13\
        );

    \I__6293\ : InMux
    port map (
            O => \N__40201\,
            I => \foc.u_Park_Transform.n17059\
        );

    \I__6292\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40195\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__40195\,
            I => \foc.u_Park_Transform.n446\
        );

    \I__6290\ : InMux
    port map (
            O => \N__40192\,
            I => \bfn_15_16_0_\
        );

    \I__6289\ : InMux
    port map (
            O => \N__40189\,
            I => \N__40186\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__40186\,
            I => \foc.u_Park_Transform.n495\
        );

    \I__6287\ : InMux
    port map (
            O => \N__40183\,
            I => \foc.u_Park_Transform.n17061\
        );

    \I__6286\ : InMux
    port map (
            O => \N__40180\,
            I => \N__40177\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__40177\,
            I => \foc.u_Park_Transform.n544\
        );

    \I__6284\ : InMux
    port map (
            O => \N__40174\,
            I => \foc.u_Park_Transform.n17062\
        );

    \I__6283\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40168\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__40168\,
            I => \foc.u_Park_Transform.n593\
        );

    \I__6281\ : InMux
    port map (
            O => \N__40165\,
            I => \foc.u_Park_Transform.n17063\
        );

    \I__6280\ : InMux
    port map (
            O => \N__40162\,
            I => \N__40159\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__40159\,
            I => \foc.u_Park_Transform.n642\
        );

    \I__6278\ : InMux
    port map (
            O => \N__40156\,
            I => \foc.u_Park_Transform.n17064\
        );

    \I__6277\ : CascadeMux
    port map (
            O => \N__40153\,
            I => \N__40150\
        );

    \I__6276\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40147\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__40147\,
            I => \foc.u_Park_Transform.n691\
        );

    \I__6274\ : InMux
    port map (
            O => \N__40144\,
            I => \foc.u_Park_Transform.n17065\
        );

    \I__6273\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40138\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__40138\,
            I => \N__40135\
        );

    \I__6271\ : Span4Mux_v
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__6270\ : Odrv4
    port map (
            O => \N__40132\,
            I => \foc.u_Park_Transform.n742_adj_2086\
        );

    \I__6269\ : InMux
    port map (
            O => \N__40129\,
            I => \foc.u_Park_Transform.n17066\
        );

    \I__6268\ : InMux
    port map (
            O => \N__40126\,
            I => \foc.u_Park_Transform.n743_adj_2096\
        );

    \I__6267\ : CascadeMux
    port map (
            O => \N__40123\,
            I => \N__40120\
        );

    \I__6266\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40117\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__40117\,
            I => \N__40114\
        );

    \I__6264\ : Span4Mux_v
    port map (
            O => \N__40114\,
            I => \N__40111\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__40111\,
            I => \foc.u_Park_Transform.n743_adj_2096_THRU_CO\
        );

    \I__6262\ : InMux
    port map (
            O => \N__40108\,
            I => \foc.u_Park_Transform.n751\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__40105\,
            I => \N__40102\
        );

    \I__6260\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40099\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__40099\,
            I => \N__40096\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__40096\,
            I => \N__40093\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__40093\,
            I => \foc.u_Park_Transform.n751_THRU_CO\
        );

    \I__6256\ : CascadeMux
    port map (
            O => \N__40090\,
            I => \N__40087\
        );

    \I__6255\ : InMux
    port map (
            O => \N__40087\,
            I => \N__40084\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__40084\,
            I => \foc.u_Park_Transform.n54\
        );

    \I__6253\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40078\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__40078\,
            I => \foc.u_Park_Transform.n103\
        );

    \I__6251\ : InMux
    port map (
            O => \N__40075\,
            I => \foc.u_Park_Transform.n17053\
        );

    \I__6250\ : CascadeMux
    port map (
            O => \N__40072\,
            I => \N__40069\
        );

    \I__6249\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40066\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__40066\,
            I => \foc.u_Park_Transform.n152\
        );

    \I__6247\ : InMux
    port map (
            O => \N__40063\,
            I => \foc.u_Park_Transform.n17054\
        );

    \I__6246\ : InMux
    port map (
            O => \N__40060\,
            I => \N__40057\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__40057\,
            I => \foc.u_Park_Transform.n201\
        );

    \I__6244\ : InMux
    port map (
            O => \N__40054\,
            I => \foc.u_Park_Transform.n17055\
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__40051\,
            I => \N__40048\
        );

    \I__6242\ : InMux
    port map (
            O => \N__40048\,
            I => \N__40045\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__40045\,
            I => \foc.u_Park_Transform.n250\
        );

    \I__6240\ : InMux
    port map (
            O => \N__40042\,
            I => \foc.u_Park_Transform.n17056\
        );

    \I__6239\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40036\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__40036\,
            I => \foc.u_Park_Transform.n299\
        );

    \I__6237\ : InMux
    port map (
            O => \N__40033\,
            I => \foc.u_Park_Transform.n17057\
        );

    \I__6236\ : CascadeMux
    port map (
            O => \N__40030\,
            I => \N__40027\
        );

    \I__6235\ : InMux
    port map (
            O => \N__40027\,
            I => \N__40024\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__40024\,
            I => \foc.u_Park_Transform.n348\
        );

    \I__6233\ : InMux
    port map (
            O => \N__40021\,
            I => \foc.u_Park_Transform.n17058\
        );

    \I__6232\ : InMux
    port map (
            O => \N__40018\,
            I => \N__40015\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__40015\,
            I => \foc.u_Park_Transform.n397\
        );

    \I__6230\ : InMux
    port map (
            O => \N__40012\,
            I => \N__40009\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__40009\,
            I => \foc.u_Park_Transform.n357\
        );

    \I__6228\ : InMux
    port map (
            O => \N__40006\,
            I => \foc.u_Park_Transform.n17029\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__40003\,
            I => \N__40000\
        );

    \I__6226\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39997\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__39997\,
            I => \foc.u_Park_Transform.n406\
        );

    \I__6224\ : InMux
    port map (
            O => \N__39994\,
            I => \bfn_15_14_0_\
        );

    \I__6223\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39988\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__39988\,
            I => \foc.u_Park_Transform.n455\
        );

    \I__6221\ : InMux
    port map (
            O => \N__39985\,
            I => \foc.u_Park_Transform.n17031\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__39982\,
            I => \N__39979\
        );

    \I__6219\ : InMux
    port map (
            O => \N__39979\,
            I => \N__39976\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__39976\,
            I => \foc.u_Park_Transform.n504\
        );

    \I__6217\ : InMux
    port map (
            O => \N__39973\,
            I => \foc.u_Park_Transform.n17032\
        );

    \I__6216\ : InMux
    port map (
            O => \N__39970\,
            I => \N__39967\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__39967\,
            I => \foc.u_Park_Transform.n553\
        );

    \I__6214\ : InMux
    port map (
            O => \N__39964\,
            I => \foc.u_Park_Transform.n17033\
        );

    \I__6213\ : CascadeMux
    port map (
            O => \N__39961\,
            I => \N__39958\
        );

    \I__6212\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39955\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__39955\,
            I => \foc.u_Park_Transform.n602\
        );

    \I__6210\ : InMux
    port map (
            O => \N__39952\,
            I => \foc.u_Park_Transform.n17034\
        );

    \I__6209\ : InMux
    port map (
            O => \N__39949\,
            I => \N__39946\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__39946\,
            I => \foc.u_Park_Transform.n651\
        );

    \I__6207\ : InMux
    port map (
            O => \N__39943\,
            I => \foc.u_Park_Transform.n17035\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__39940\,
            I => \N__39937\
        );

    \I__6205\ : InMux
    port map (
            O => \N__39937\,
            I => \N__39934\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__39934\,
            I => \foc.u_Park_Transform.n700\
        );

    \I__6203\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39928\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__39928\,
            I => \N__39925\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__39925\,
            I => \N__39922\
        );

    \I__6200\ : Odrv4
    port map (
            O => \N__39922\,
            I => \foc.u_Park_Transform.n750_adj_2117\
        );

    \I__6199\ : InMux
    port map (
            O => \N__39919\,
            I => \foc.u_Park_Transform.n17036\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__39916\,
            I => \N__39913\
        );

    \I__6197\ : InMux
    port map (
            O => \N__39913\,
            I => \N__39910\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__39910\,
            I => \foc.u_Park_Transform.n694_adj_2097\
        );

    \I__6195\ : InMux
    port map (
            O => \N__39907\,
            I => \N__39904\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__39904\,
            I => \N__39901\
        );

    \I__6193\ : Span4Mux_h
    port map (
            O => \N__39901\,
            I => \N__39898\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__39898\,
            I => \foc.u_Park_Transform.n742\
        );

    \I__6191\ : InMux
    port map (
            O => \N__39895\,
            I => \foc.u_Park_Transform.n17249\
        );

    \I__6190\ : InMux
    port map (
            O => \N__39892\,
            I => \foc.u_Park_Transform.n743\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__39889\,
            I => \N__39886\
        );

    \I__6188\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39883\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__39883\,
            I => \N__39880\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__39880\,
            I => \N__39877\
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__39877\,
            I => \foc.u_Park_Transform.n743_THRU_CO\
        );

    \I__6184\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39871\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__39871\,
            I => \foc.u_Park_Transform.n63\
        );

    \I__6182\ : InMux
    port map (
            O => \N__39868\,
            I => \foc.u_Park_Transform.n17023\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__39865\,
            I => \N__39862\
        );

    \I__6180\ : InMux
    port map (
            O => \N__39862\,
            I => \N__39859\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__39859\,
            I => \foc.u_Park_Transform.n112\
        );

    \I__6178\ : InMux
    port map (
            O => \N__39856\,
            I => \foc.u_Park_Transform.n17024\
        );

    \I__6177\ : InMux
    port map (
            O => \N__39853\,
            I => \N__39850\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__39850\,
            I => \foc.u_Park_Transform.n161\
        );

    \I__6175\ : InMux
    port map (
            O => \N__39847\,
            I => \foc.u_Park_Transform.n17025\
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__39844\,
            I => \N__39841\
        );

    \I__6173\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39838\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__39838\,
            I => \foc.u_Park_Transform.n210\
        );

    \I__6171\ : InMux
    port map (
            O => \N__39835\,
            I => \foc.u_Park_Transform.n17026\
        );

    \I__6170\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39829\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__39829\,
            I => \foc.u_Park_Transform.n259\
        );

    \I__6168\ : InMux
    port map (
            O => \N__39826\,
            I => \foc.u_Park_Transform.n17027\
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__39823\,
            I => \N__39820\
        );

    \I__6166\ : InMux
    port map (
            O => \N__39820\,
            I => \N__39817\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__39817\,
            I => \N__39814\
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__39814\,
            I => \foc.u_Park_Transform.n308\
        );

    \I__6163\ : InMux
    port map (
            O => \N__39811\,
            I => \foc.u_Park_Transform.n17028\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__39808\,
            I => \N__39805\
        );

    \I__6161\ : InMux
    port map (
            O => \N__39805\,
            I => \N__39802\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__39802\,
            I => \N__39799\
        );

    \I__6159\ : Odrv4
    port map (
            O => \N__39799\,
            I => \foc.u_Park_Transform.n348_adj_2082\
        );

    \I__6158\ : InMux
    port map (
            O => \N__39796\,
            I => \foc.u_Park_Transform.n17241\
        );

    \I__6157\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39790\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__39790\,
            I => \foc.u_Park_Transform.n351_adj_2108\
        );

    \I__6155\ : InMux
    port map (
            O => \N__39787\,
            I => \N__39784\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__39784\,
            I => \foc.u_Park_Transform.n397_adj_2081\
        );

    \I__6153\ : InMux
    port map (
            O => \N__39781\,
            I => \foc.u_Park_Transform.n17242\
        );

    \I__6152\ : CascadeMux
    port map (
            O => \N__39778\,
            I => \N__39775\
        );

    \I__6151\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39772\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__39772\,
            I => \foc.u_Park_Transform.n400_adj_2106\
        );

    \I__6149\ : CascadeMux
    port map (
            O => \N__39769\,
            I => \N__39766\
        );

    \I__6148\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39763\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__39763\,
            I => \N__39760\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__39760\,
            I => \foc.u_Park_Transform.n446_adj_2079\
        );

    \I__6145\ : InMux
    port map (
            O => \N__39757\,
            I => \bfn_15_12_0_\
        );

    \I__6144\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39751\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__39751\,
            I => \foc.u_Park_Transform.n449_adj_2103\
        );

    \I__6142\ : InMux
    port map (
            O => \N__39748\,
            I => \N__39745\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__39745\,
            I => \N__39742\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__39742\,
            I => \foc.u_Park_Transform.n495_adj_2077\
        );

    \I__6139\ : InMux
    port map (
            O => \N__39739\,
            I => \foc.u_Park_Transform.n17244\
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__39736\,
            I => \N__39733\
        );

    \I__6137\ : InMux
    port map (
            O => \N__39733\,
            I => \N__39730\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__39730\,
            I => \foc.u_Park_Transform.n498_adj_2102\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__39727\,
            I => \N__39724\
        );

    \I__6134\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39721\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__39721\,
            I => \N__39718\
        );

    \I__6132\ : Odrv4
    port map (
            O => \N__39718\,
            I => \foc.u_Park_Transform.n544_adj_2074\
        );

    \I__6131\ : InMux
    port map (
            O => \N__39715\,
            I => \foc.u_Park_Transform.n17245\
        );

    \I__6130\ : InMux
    port map (
            O => \N__39712\,
            I => \N__39709\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__39709\,
            I => \foc.u_Park_Transform.n547_adj_2100\
        );

    \I__6128\ : InMux
    port map (
            O => \N__39706\,
            I => \N__39703\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__39703\,
            I => \N__39700\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__39700\,
            I => \foc.u_Park_Transform.n593_adj_2073\
        );

    \I__6125\ : InMux
    port map (
            O => \N__39697\,
            I => \foc.u_Park_Transform.n17246\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__39694\,
            I => \N__39691\
        );

    \I__6123\ : InMux
    port map (
            O => \N__39691\,
            I => \N__39688\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__39688\,
            I => \foc.u_Park_Transform.n596_adj_2099\
        );

    \I__6121\ : CascadeMux
    port map (
            O => \N__39685\,
            I => \N__39682\
        );

    \I__6120\ : InMux
    port map (
            O => \N__39682\,
            I => \N__39679\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__39679\,
            I => \N__39676\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__39676\,
            I => \foc.u_Park_Transform.n642_adj_2072\
        );

    \I__6117\ : InMux
    port map (
            O => \N__39673\,
            I => \foc.u_Park_Transform.n17247\
        );

    \I__6116\ : InMux
    port map (
            O => \N__39670\,
            I => \N__39667\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__39667\,
            I => \foc.u_Park_Transform.n645_adj_2098\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__39664\,
            I => \N__39661\
        );

    \I__6113\ : InMux
    port map (
            O => \N__39661\,
            I => \N__39658\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__39658\,
            I => \N__39655\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__39655\,
            I => \foc.u_Park_Transform.n691_adj_2071\
        );

    \I__6110\ : InMux
    port map (
            O => \N__39652\,
            I => \foc.u_Park_Transform.n17248\
        );

    \I__6109\ : CascadeMux
    port map (
            O => \N__39649\,
            I => \N__39646\
        );

    \I__6108\ : InMux
    port map (
            O => \N__39646\,
            I => \N__39642\
        );

    \I__6107\ : InMux
    port map (
            O => \N__39645\,
            I => \N__39639\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39634\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39634\
        );

    \I__6104\ : Span4Mux_v
    port map (
            O => \N__39634\,
            I => \N__39631\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__39631\,
            I => \foc.u_Park_Transform.n738\
        );

    \I__6102\ : InMux
    port map (
            O => \N__39628\,
            I => \foc.u_Park_Transform.n17264\
        );

    \I__6101\ : InMux
    port map (
            O => \N__39625\,
            I => \foc.u_Park_Transform.n739\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__39622\,
            I => \N__39619\
        );

    \I__6099\ : InMux
    port map (
            O => \N__39619\,
            I => \N__39616\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__39616\,
            I => \N__39613\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__39613\,
            I => \N__39610\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__39610\,
            I => \foc.u_Park_Transform.n739_THRU_CO\
        );

    \I__6095\ : InMux
    port map (
            O => \N__39607\,
            I => \N__39604\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__39604\,
            I => \N__39601\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__39601\,
            I => \foc.u_Park_Transform.n54_adj_2095\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__39598\,
            I => \N__39595\
        );

    \I__6091\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39592\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__39592\,
            I => \foc.u_Park_Transform.n57_adj_2116\
        );

    \I__6089\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39586\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__39586\,
            I => \N__39583\
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__39583\,
            I => \foc.u_Park_Transform.n103_adj_2092\
        );

    \I__6086\ : InMux
    port map (
            O => \N__39580\,
            I => \foc.u_Park_Transform.n17236\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__39577\,
            I => \N__39574\
        );

    \I__6084\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39571\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__39571\,
            I => \foc.u_Park_Transform.n106_adj_2115\
        );

    \I__6082\ : CascadeMux
    port map (
            O => \N__39568\,
            I => \N__39565\
        );

    \I__6081\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39562\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__39562\,
            I => \N__39559\
        );

    \I__6079\ : Odrv12
    port map (
            O => \N__39559\,
            I => \foc.u_Park_Transform.n152_adj_2088\
        );

    \I__6078\ : InMux
    port map (
            O => \N__39556\,
            I => \foc.u_Park_Transform.n17237\
        );

    \I__6077\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39550\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__39550\,
            I => \foc.u_Park_Transform.n155_adj_2114\
        );

    \I__6075\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39544\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__39544\,
            I => \N__39541\
        );

    \I__6073\ : Odrv12
    port map (
            O => \N__39541\,
            I => \foc.u_Park_Transform.n201_adj_2085\
        );

    \I__6072\ : InMux
    port map (
            O => \N__39538\,
            I => \foc.u_Park_Transform.n17238\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__39535\,
            I => \N__39532\
        );

    \I__6070\ : InMux
    port map (
            O => \N__39532\,
            I => \N__39529\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__39529\,
            I => \foc.u_Park_Transform.n204_adj_2113\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__39526\,
            I => \N__39523\
        );

    \I__6067\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39520\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__39520\,
            I => \N__39517\
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__39517\,
            I => \foc.u_Park_Transform.n250_adj_2084\
        );

    \I__6064\ : InMux
    port map (
            O => \N__39514\,
            I => \foc.u_Park_Transform.n17239\
        );

    \I__6063\ : InMux
    port map (
            O => \N__39511\,
            I => \N__39508\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__39508\,
            I => \foc.u_Park_Transform.n253_adj_2112\
        );

    \I__6061\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39502\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__39502\,
            I => \N__39499\
        );

    \I__6059\ : Odrv4
    port map (
            O => \N__39499\,
            I => \foc.u_Park_Transform.n299_adj_2083\
        );

    \I__6058\ : InMux
    port map (
            O => \N__39496\,
            I => \foc.u_Park_Transform.n17240\
        );

    \I__6057\ : CascadeMux
    port map (
            O => \N__39493\,
            I => \N__39490\
        );

    \I__6056\ : InMux
    port map (
            O => \N__39490\,
            I => \N__39487\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__39487\,
            I => \foc.u_Park_Transform.n302_adj_2111\
        );

    \I__6054\ : InMux
    port map (
            O => \N__39484\,
            I => \N__39481\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__39481\,
            I => \N__39478\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__39478\,
            I => \foc.u_Park_Transform.Product1_mul_temp_7\
        );

    \I__6051\ : InMux
    port map (
            O => \N__39475\,
            I => \foc.u_Park_Transform.n17256\
        );

    \I__6050\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39469\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__39469\,
            I => \N__39466\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__39466\,
            I => \N__39463\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__39463\,
            I => \foc.u_Park_Transform.Product1_mul_temp_8\
        );

    \I__6046\ : InMux
    port map (
            O => \N__39460\,
            I => \foc.u_Park_Transform.n17257\
        );

    \I__6045\ : InMux
    port map (
            O => \N__39457\,
            I => \N__39454\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__39454\,
            I => \N__39451\
        );

    \I__6043\ : Sp12to4
    port map (
            O => \N__39451\,
            I => \N__39448\
        );

    \I__6042\ : Odrv12
    port map (
            O => \N__39448\,
            I => \foc.u_Park_Transform.Product1_mul_temp_9\
        );

    \I__6041\ : InMux
    port map (
            O => \N__39445\,
            I => \bfn_15_10_0_\
        );

    \I__6040\ : InMux
    port map (
            O => \N__39442\,
            I => \N__39439\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__39439\,
            I => \N__39436\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__39436\,
            I => \N__39433\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__39433\,
            I => \foc.u_Park_Transform.Product1_mul_temp_10\
        );

    \I__6036\ : InMux
    port map (
            O => \N__39430\,
            I => \foc.u_Park_Transform.n17259\
        );

    \I__6035\ : InMux
    port map (
            O => \N__39427\,
            I => \N__39424\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__39424\,
            I => \N__39421\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__39421\,
            I => \foc.u_Park_Transform.Product1_mul_temp_11\
        );

    \I__6032\ : InMux
    port map (
            O => \N__39418\,
            I => \foc.u_Park_Transform.n17260\
        );

    \I__6031\ : InMux
    port map (
            O => \N__39415\,
            I => \N__39412\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__39412\,
            I => \N__39409\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__39409\,
            I => \foc.u_Park_Transform.Product1_mul_temp_12\
        );

    \I__6028\ : InMux
    port map (
            O => \N__39406\,
            I => \foc.u_Park_Transform.n17261\
        );

    \I__6027\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39400\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__39400\,
            I => \N__39397\
        );

    \I__6025\ : Odrv4
    port map (
            O => \N__39397\,
            I => \foc.u_Park_Transform.Product1_mul_temp_13\
        );

    \I__6024\ : InMux
    port map (
            O => \N__39394\,
            I => \foc.u_Park_Transform.n17262\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__39391\,
            I => \N__39381\
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__39390\,
            I => \N__39377\
        );

    \I__6021\ : CascadeMux
    port map (
            O => \N__39389\,
            I => \N__39373\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__39388\,
            I => \N__39369\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__39387\,
            I => \N__39366\
        );

    \I__6018\ : CascadeMux
    port map (
            O => \N__39386\,
            I => \N__39362\
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__39385\,
            I => \N__39358\
        );

    \I__6016\ : CascadeMux
    port map (
            O => \N__39384\,
            I => \N__39354\
        );

    \I__6015\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39345\
        );

    \I__6014\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39330\
        );

    \I__6013\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39330\
        );

    \I__6012\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39330\
        );

    \I__6011\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39330\
        );

    \I__6010\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39330\
        );

    \I__6009\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39330\
        );

    \I__6008\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39330\
        );

    \I__6007\ : InMux
    port map (
            O => \N__39365\,
            I => \N__39317\
        );

    \I__6006\ : InMux
    port map (
            O => \N__39362\,
            I => \N__39317\
        );

    \I__6005\ : InMux
    port map (
            O => \N__39361\,
            I => \N__39317\
        );

    \I__6004\ : InMux
    port map (
            O => \N__39358\,
            I => \N__39317\
        );

    \I__6003\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39317\
        );

    \I__6002\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39317\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__39353\,
            I => \N__39310\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__39352\,
            I => \N__39307\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__39351\,
            I => \N__39304\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__39350\,
            I => \N__39301\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__39349\,
            I => \N__39298\
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__39348\,
            I => \N__39295\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__39345\,
            I => \N__39292\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__39330\,
            I => \N__39287\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__39317\,
            I => \N__39287\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__39316\,
            I => \N__39283\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__39315\,
            I => \N__39279\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__39314\,
            I => \N__39275\
        );

    \I__5989\ : CascadeMux
    port map (
            O => \N__39313\,
            I => \N__39271\
        );

    \I__5988\ : InMux
    port map (
            O => \N__39310\,
            I => \N__39264\
        );

    \I__5987\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39264\
        );

    \I__5986\ : InMux
    port map (
            O => \N__39304\,
            I => \N__39264\
        );

    \I__5985\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39257\
        );

    \I__5984\ : InMux
    port map (
            O => \N__39298\,
            I => \N__39257\
        );

    \I__5983\ : InMux
    port map (
            O => \N__39295\,
            I => \N__39257\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__39292\,
            I => \N__39252\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__39287\,
            I => \N__39252\
        );

    \I__5980\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39235\
        );

    \I__5979\ : InMux
    port map (
            O => \N__39283\,
            I => \N__39235\
        );

    \I__5978\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39235\
        );

    \I__5977\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39235\
        );

    \I__5976\ : InMux
    port map (
            O => \N__39278\,
            I => \N__39235\
        );

    \I__5975\ : InMux
    port map (
            O => \N__39275\,
            I => \N__39235\
        );

    \I__5974\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39235\
        );

    \I__5973\ : InMux
    port map (
            O => \N__39271\,
            I => \N__39235\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__39264\,
            I => \N__39232\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__39257\,
            I => \N__39229\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__39252\,
            I => \N__39224\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__39235\,
            I => \N__39224\
        );

    \I__5968\ : Span4Mux_v
    port map (
            O => \N__39232\,
            I => \N__39219\
        );

    \I__5967\ : Span4Mux_v
    port map (
            O => \N__39229\,
            I => \N__39219\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__39224\,
            I => \N__39216\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__39219\,
            I => \foc.u_Park_Transform.dCurrent_2\
        );

    \I__5964\ : Odrv4
    port map (
            O => \N__39216\,
            I => \foc.u_Park_Transform.dCurrent_2\
        );

    \I__5963\ : InMux
    port map (
            O => \N__39211\,
            I => \N__39208\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__39208\,
            I => \N__39205\
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__39205\,
            I => \foc.u_Park_Transform.Product1_mul_temp_14\
        );

    \I__5960\ : InMux
    port map (
            O => \N__39202\,
            I => \foc.u_Park_Transform.n17263\
        );

    \I__5959\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39196\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__39196\,
            I => \N__39192\
        );

    \I__5957\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39189\
        );

    \I__5956\ : Span4Mux_v
    port map (
            O => \N__39192\,
            I => \N__39186\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39183\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__39186\,
            I => \N__39178\
        );

    \I__5953\ : Span4Mux_h
    port map (
            O => \N__39183\,
            I => \N__39178\
        );

    \I__5952\ : Odrv4
    port map (
            O => \N__39178\,
            I => \foc.u_Park_Transform.n737\
        );

    \I__5951\ : InMux
    port map (
            O => \N__39175\,
            I => \N__39172\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__39172\,
            I => \N__39169\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__39169\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n2\
        );

    \I__5948\ : InMux
    port map (
            O => \N__39166\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15804\
        );

    \I__5947\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__39160\,
            I => \foc.dCurrent_26\
        );

    \I__5945\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39154\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__39154\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n7\
        );

    \I__5943\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39148\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__39148\,
            I => \N__39145\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__39145\,
            I => \N__39142\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__39142\,
            I => \foc.dCurrent_3\
        );

    \I__5939\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39136\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__39136\,
            I => \N__39133\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__39133\,
            I => \foc.u_Park_Transform.Product1_mul_temp_2\
        );

    \I__5936\ : InMux
    port map (
            O => \N__39130\,
            I => \foc.u_Park_Transform.n17251\
        );

    \I__5935\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39124\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39121\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__39121\,
            I => \foc.u_Park_Transform.Product1_mul_temp_3\
        );

    \I__5932\ : InMux
    port map (
            O => \N__39118\,
            I => \foc.u_Park_Transform.n17252\
        );

    \I__5931\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39112\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__39112\,
            I => \N__39109\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__39109\,
            I => \foc.u_Park_Transform.Product1_mul_temp_4\
        );

    \I__5928\ : InMux
    port map (
            O => \N__39106\,
            I => \foc.u_Park_Transform.n17253\
        );

    \I__5927\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39100\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__39100\,
            I => \N__39097\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__39097\,
            I => \foc.u_Park_Transform.Product1_mul_temp_5\
        );

    \I__5924\ : InMux
    port map (
            O => \N__39094\,
            I => \foc.u_Park_Transform.n17254\
        );

    \I__5923\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39088\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__39088\,
            I => \N__39085\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__39085\,
            I => \foc.u_Park_Transform.Product1_mul_temp_6\
        );

    \I__5920\ : InMux
    port map (
            O => \N__39082\,
            I => \foc.u_Park_Transform.n17255\
        );

    \I__5919\ : InMux
    port map (
            O => \N__39079\,
            I => \N__39076\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__39076\,
            I => \N__39073\
        );

    \I__5917\ : Span4Mux_v
    port map (
            O => \N__39073\,
            I => \N__39070\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__39070\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n11\
        );

    \I__5915\ : InMux
    port map (
            O => \N__39067\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15795\
        );

    \I__5914\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39061\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__39058\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__39058\,
            I => \N__39055\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__39055\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n10\
        );

    \I__5910\ : InMux
    port map (
            O => \N__39052\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15796\
        );

    \I__5909\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39046\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__39046\,
            I => \N__39043\
        );

    \I__5907\ : Span4Mux_h
    port map (
            O => \N__39043\,
            I => \N__39040\
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__39040\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n9\
        );

    \I__5905\ : InMux
    port map (
            O => \N__39037\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15797\
        );

    \I__5904\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39031\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__39031\,
            I => \N__39028\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__39028\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n8\
        );

    \I__5901\ : InMux
    port map (
            O => \N__39025\,
            I => \bfn_15_8_0_\
        );

    \I__5900\ : InMux
    port map (
            O => \N__39022\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15799\
        );

    \I__5899\ : InMux
    port map (
            O => \N__39019\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15800\
        );

    \I__5898\ : InMux
    port map (
            O => \N__39016\,
            I => \N__39013\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__39013\,
            I => \N__39010\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__39010\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n5\
        );

    \I__5895\ : InMux
    port map (
            O => \N__39007\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15801\
        );

    \I__5894\ : InMux
    port map (
            O => \N__39004\,
            I => \N__39001\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__39001\,
            I => \N__38998\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__38998\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n4_adj_515\
        );

    \I__5891\ : InMux
    port map (
            O => \N__38995\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15802\
        );

    \I__5890\ : InMux
    port map (
            O => \N__38992\,
            I => \N__38989\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__38986\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n3\
        );

    \I__5887\ : InMux
    port map (
            O => \N__38983\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15803\
        );

    \I__5886\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38977\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__38977\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n19\
        );

    \I__5884\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38971\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__38971\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n18\
        );

    \I__5882\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38965\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__38965\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n17\
        );

    \I__5880\ : InMux
    port map (
            O => \N__38962\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15789\
        );

    \I__5879\ : InMux
    port map (
            O => \N__38959\,
            I => \N__38956\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__38956\,
            I => \N__38953\
        );

    \I__5877\ : Span4Mux_h
    port map (
            O => \N__38953\,
            I => \N__38950\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__38950\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n16\
        );

    \I__5875\ : InMux
    port map (
            O => \N__38947\,
            I => \bfn_15_7_0_\
        );

    \I__5874\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38941\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__38941\,
            I => \N__38938\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__38938\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15_adj_518\
        );

    \I__5871\ : InMux
    port map (
            O => \N__38935\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15791\
        );

    \I__5870\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38929\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__38929\,
            I => \N__38926\
        );

    \I__5868\ : Span4Mux_h
    port map (
            O => \N__38926\,
            I => \N__38923\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__38923\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n14_adj_517\
        );

    \I__5866\ : InMux
    port map (
            O => \N__38920\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15792\
        );

    \I__5865\ : InMux
    port map (
            O => \N__38917\,
            I => \N__38914\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38911\
        );

    \I__5863\ : Span4Mux_h
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__38908\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n13\
        );

    \I__5861\ : InMux
    port map (
            O => \N__38905\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15793\
        );

    \I__5860\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38899\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__38899\,
            I => \N__38896\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__38896\,
            I => \N__38893\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__38893\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n12_adj_516\
        );

    \I__5856\ : InMux
    port map (
            O => \N__38890\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n15794\
        );

    \I__5855\ : InMux
    port map (
            O => \N__38887\,
            I => \N__38884\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__38884\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n28\
        );

    \I__5853\ : InMux
    port map (
            O => \N__38881\,
            I => \N__38878\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__38878\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n27\
        );

    \I__5851\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38872\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__38872\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n26\
        );

    \I__5849\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38866\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__38866\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n25\
        );

    \I__5847\ : InMux
    port map (
            O => \N__38863\,
            I => \N__38860\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__38860\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n24\
        );

    \I__5845\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38854\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__38854\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n23\
        );

    \I__5843\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38848\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__38848\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n22\
        );

    \I__5841\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38842\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__38842\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n21\
        );

    \I__5839\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38836\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__38836\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n20\
        );

    \I__5837\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38830\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__38830\,
            I => \N__38827\
        );

    \I__5835\ : Odrv4
    port map (
            O => \N__38827\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n602_adj_671\
        );

    \I__5834\ : InMux
    port map (
            O => \N__38824\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18043\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__38821\,
            I => \N__38818\
        );

    \I__5832\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38815\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__38815\,
            I => \N__38812\
        );

    \I__5830\ : Odrv12
    port map (
            O => \N__38812\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n651_adj_670\
        );

    \I__5829\ : InMux
    port map (
            O => \N__38809\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18044\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__38806\,
            I => \N__38803\
        );

    \I__5827\ : InMux
    port map (
            O => \N__38803\,
            I => \N__38800\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__38800\,
            I => \N__38797\
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__38797\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n700_adj_669\
        );

    \I__5824\ : InMux
    port map (
            O => \N__38794\,
            I => \N__38791\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__38791\,
            I => \N__38788\
        );

    \I__5822\ : Span4Mux_v
    port map (
            O => \N__38788\,
            I => \N__38785\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__38785\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n750_adj_683\
        );

    \I__5820\ : InMux
    port map (
            O => \N__38782\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18045\
        );

    \I__5819\ : InMux
    port map (
            O => \N__38779\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__38776\,
            I => \N__38773\
        );

    \I__5817\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38770\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__38770\,
            I => \N__38767\
        );

    \I__5815\ : Span4Mux_v
    port map (
            O => \N__38767\,
            I => \N__38764\
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__38764\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_CO\
        );

    \I__5813\ : InMux
    port map (
            O => \N__38761\,
            I => \N__38758\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__38758\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n30\
        );

    \I__5811\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38752\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__38752\,
            I => \foc.u_DQ_Current_Control.u_D_Current_Control.n29\
        );

    \I__5809\ : InMux
    port map (
            O => \N__38749\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18034\
        );

    \I__5808\ : InMux
    port map (
            O => \N__38746\,
            I => \N__38743\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__38743\,
            I => \N__38740\
        );

    \I__5806\ : Odrv12
    port map (
            O => \N__38740\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n210_adj_679\
        );

    \I__5805\ : InMux
    port map (
            O => \N__38737\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18035\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__38734\,
            I => \N__38731\
        );

    \I__5803\ : InMux
    port map (
            O => \N__38731\,
            I => \N__38728\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__38728\,
            I => \N__38725\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__38725\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n259_adj_678\
        );

    \I__5800\ : InMux
    port map (
            O => \N__38722\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18036\
        );

    \I__5799\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38716\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__38716\,
            I => \N__38713\
        );

    \I__5797\ : Odrv12
    port map (
            O => \N__38713\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n308_adj_677\
        );

    \I__5796\ : InMux
    port map (
            O => \N__38710\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18037\
        );

    \I__5795\ : CascadeMux
    port map (
            O => \N__38707\,
            I => \N__38704\
        );

    \I__5794\ : InMux
    port map (
            O => \N__38704\,
            I => \N__38701\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__38701\,
            I => \N__38698\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__38698\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n357_adj_676\
        );

    \I__5791\ : InMux
    port map (
            O => \N__38695\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18038\
        );

    \I__5790\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38689\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__38689\,
            I => \N__38686\
        );

    \I__5788\ : Odrv12
    port map (
            O => \N__38686\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n406_adj_675\
        );

    \I__5787\ : InMux
    port map (
            O => \N__38683\,
            I => \bfn_14_26_0_\
        );

    \I__5786\ : CascadeMux
    port map (
            O => \N__38680\,
            I => \N__38677\
        );

    \I__5785\ : InMux
    port map (
            O => \N__38677\,
            I => \N__38674\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__38674\,
            I => \N__38671\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__38671\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n455_adj_674\
        );

    \I__5782\ : InMux
    port map (
            O => \N__38668\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18040\
        );

    \I__5781\ : InMux
    port map (
            O => \N__38665\,
            I => \N__38662\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__38662\,
            I => \N__38659\
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__38659\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n504_adj_673\
        );

    \I__5778\ : InMux
    port map (
            O => \N__38656\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18041\
        );

    \I__5777\ : CascadeMux
    port map (
            O => \N__38653\,
            I => \N__38650\
        );

    \I__5776\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38647\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__38647\,
            I => \N__38644\
        );

    \I__5774\ : Odrv12
    port map (
            O => \N__38644\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n553_adj_672\
        );

    \I__5773\ : InMux
    port map (
            O => \N__38641\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18042\
        );

    \I__5772\ : InMux
    port map (
            O => \N__38638\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18057\
        );

    \I__5771\ : InMux
    port map (
            O => \N__38635\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18058\
        );

    \I__5770\ : InMux
    port map (
            O => \N__38632\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18059\
        );

    \I__5769\ : InMux
    port map (
            O => \N__38629\,
            I => \N__38626\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__38626\,
            I => \N__38623\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__38623\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n754_adj_667\
        );

    \I__5766\ : InMux
    port map (
            O => \N__38620\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18060\
        );

    \I__5765\ : InMux
    port map (
            O => \N__38617\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__38614\,
            I => \N__38611\
        );

    \I__5763\ : InMux
    port map (
            O => \N__38611\,
            I => \N__38608\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__38608\,
            I => \N__38605\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__38605\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_CO\
        );

    \I__5760\ : CascadeMux
    port map (
            O => \N__38602\,
            I => \N__38599\
        );

    \I__5759\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38596\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__38596\,
            I => \N__38593\
        );

    \I__5757\ : Odrv4
    port map (
            O => \N__38593\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n63_adj_682\
        );

    \I__5756\ : InMux
    port map (
            O => \N__38590\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18032\
        );

    \I__5755\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38584\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__38584\,
            I => \N__38581\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__38581\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n112_adj_681\
        );

    \I__5752\ : InMux
    port map (
            O => \N__38578\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18033\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__38575\,
            I => \N__38572\
        );

    \I__5750\ : InMux
    port map (
            O => \N__38572\,
            I => \N__38569\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__38569\,
            I => \N__38566\
        );

    \I__5748\ : Odrv12
    port map (
            O => \N__38566\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n161_adj_680\
        );

    \I__5747\ : InMux
    port map (
            O => \N__38563\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18048\
        );

    \I__5746\ : InMux
    port map (
            O => \N__38560\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18049\
        );

    \I__5745\ : InMux
    port map (
            O => \N__38557\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18050\
        );

    \I__5744\ : InMux
    port map (
            O => \N__38554\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18051\
        );

    \I__5743\ : InMux
    port map (
            O => \N__38551\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18052\
        );

    \I__5742\ : InMux
    port map (
            O => \N__38548\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18053\
        );

    \I__5741\ : InMux
    port map (
            O => \N__38545\,
            I => \bfn_14_24_0_\
        );

    \I__5740\ : InMux
    port map (
            O => \N__38542\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18055\
        );

    \I__5739\ : InMux
    port map (
            O => \N__38539\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18056\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__38536\,
            I => \N__38533\
        );

    \I__5737\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38530\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__38530\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n280_adj_743\
        );

    \I__5735\ : InMux
    port map (
            O => \N__38527\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17730\
        );

    \I__5734\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38521\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__38521\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n329_adj_740\
        );

    \I__5732\ : InMux
    port map (
            O => \N__38518\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17731\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__38515\,
            I => \N__38512\
        );

    \I__5730\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38509\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__38509\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n378_adj_739\
        );

    \I__5728\ : InMux
    port map (
            O => \N__38506\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17732\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__38503\,
            I => \N__38499\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__38502\,
            I => \N__38496\
        );

    \I__5725\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38492\
        );

    \I__5724\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38487\
        );

    \I__5723\ : InMux
    port map (
            O => \N__38495\,
            I => \N__38487\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__38492\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__38487\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738\
        );

    \I__5720\ : InMux
    port map (
            O => \N__38482\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17733\
        );

    \I__5719\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38476\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__38476\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n782_adj_735\
        );

    \I__5717\ : InMux
    port map (
            O => \N__38473\,
            I => \bfn_14_22_0_\
        );

    \I__5716\ : InMux
    port map (
            O => \N__38470\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__38467\,
            I => \N__38464\
        );

    \I__5714\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38461\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__38461\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_CO\
        );

    \I__5712\ : InMux
    port map (
            O => \N__38458\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18047\
        );

    \I__5711\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38452\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__38452\,
            I => \N__38449\
        );

    \I__5709\ : Span4Mux_v
    port map (
            O => \N__38449\,
            I => \N__38446\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__38446\,
            I => \foc.u_Park_Transform.Product4_mul_temp_29\
        );

    \I__5707\ : InMux
    port map (
            O => \N__38443\,
            I => \foc.u_Park_Transform.n15774\
        );

    \I__5706\ : InMux
    port map (
            O => \N__38440\,
            I => \N__38437\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__38437\,
            I => \foc.qCurrent_21\
        );

    \I__5704\ : InMux
    port map (
            O => \N__38434\,
            I => \N__38431\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__38431\,
            I => \foc.qCurrent_29\
        );

    \I__5702\ : InMux
    port map (
            O => \N__38428\,
            I => \N__38425\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__38425\,
            I => \foc.qCurrent_23\
        );

    \I__5700\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38419\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__38419\,
            I => \foc.qCurrent_30\
        );

    \I__5698\ : CascadeMux
    port map (
            O => \N__38416\,
            I => \N__38413\
        );

    \I__5697\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38410\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__38410\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n84_adj_749\
        );

    \I__5695\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38404\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__38404\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n133_adj_747\
        );

    \I__5693\ : InMux
    port map (
            O => \N__38401\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17727\
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__38398\,
            I => \N__38395\
        );

    \I__5691\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38392\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__38392\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n182_adj_745\
        );

    \I__5689\ : InMux
    port map (
            O => \N__38389\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17728\
        );

    \I__5688\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38383\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__38383\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n231_adj_744\
        );

    \I__5686\ : InMux
    port map (
            O => \N__38380\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17729\
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__38377\,
            I => \N__38374\
        );

    \I__5684\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38371\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38368\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__38368\,
            I => \N__38365\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__38365\,
            I => \foc.u_Park_Transform.Product4_mul_temp_21\
        );

    \I__5680\ : InMux
    port map (
            O => \N__38362\,
            I => \foc.u_Park_Transform.n15766\
        );

    \I__5679\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38356\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__38356\,
            I => \N__38353\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__38353\,
            I => \N__38350\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__38350\,
            I => \foc.u_Park_Transform.Product4_mul_temp_22\
        );

    \I__5675\ : InMux
    port map (
            O => \N__38347\,
            I => \foc.u_Park_Transform.n15767\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__38344\,
            I => \N__38341\
        );

    \I__5673\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38338\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__38338\,
            I => \N__38335\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__38335\,
            I => \N__38332\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__38332\,
            I => \foc.u_Park_Transform.Product4_mul_temp_23\
        );

    \I__5669\ : InMux
    port map (
            O => \N__38329\,
            I => \foc.u_Park_Transform.n15768\
        );

    \I__5668\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38323\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__38323\,
            I => \N__38320\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__38320\,
            I => \N__38317\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__38317\,
            I => \foc.u_Park_Transform.Product4_mul_temp_24\
        );

    \I__5664\ : InMux
    port map (
            O => \N__38314\,
            I => \foc.u_Park_Transform.n15769\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__38311\,
            I => \N__38308\
        );

    \I__5662\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__38305\,
            I => \N__38302\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__38302\,
            I => \N__38299\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__38299\,
            I => \foc.u_Park_Transform.Product4_mul_temp_25\
        );

    \I__5658\ : InMux
    port map (
            O => \N__38296\,
            I => \foc.u_Park_Transform.n15770\
        );

    \I__5657\ : InMux
    port map (
            O => \N__38293\,
            I => \N__38290\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__38290\,
            I => \N__38287\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__38287\,
            I => \N__38284\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__38284\,
            I => \foc.u_Park_Transform.Product4_mul_temp_26\
        );

    \I__5653\ : InMux
    port map (
            O => \N__38281\,
            I => \bfn_14_20_0_\
        );

    \I__5652\ : CascadeMux
    port map (
            O => \N__38278\,
            I => \N__38275\
        );

    \I__5651\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__38272\,
            I => \N__38269\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__38269\,
            I => \N__38266\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__38266\,
            I => \foc.u_Park_Transform.Product4_mul_temp_27\
        );

    \I__5647\ : InMux
    port map (
            O => \N__38263\,
            I => \foc.u_Park_Transform.n15772\
        );

    \I__5646\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38257\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38254\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__38254\,
            I => \N__38251\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__38251\,
            I => \foc.u_Park_Transform.Product4_mul_temp_28\
        );

    \I__5642\ : InMux
    port map (
            O => \N__38248\,
            I => \foc.u_Park_Transform.n15773\
        );

    \I__5641\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38242\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38239\
        );

    \I__5639\ : Odrv12
    port map (
            O => \N__38239\,
            I => \foc.u_Park_Transform.Product4_mul_temp_12\
        );

    \I__5638\ : InMux
    port map (
            O => \N__38236\,
            I => \foc.u_Park_Transform.n15757\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__38233\,
            I => \N__38230\
        );

    \I__5636\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38224\
        );

    \I__5634\ : Odrv4
    port map (
            O => \N__38224\,
            I => \foc.u_Park_Transform.Product4_mul_temp_13\
        );

    \I__5633\ : InMux
    port map (
            O => \N__38221\,
            I => \foc.u_Park_Transform.n15758\
        );

    \I__5632\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38215\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__38215\,
            I => \N__38212\
        );

    \I__5630\ : Odrv4
    port map (
            O => \N__38212\,
            I => \foc.u_Park_Transform.Product4_mul_temp_14\
        );

    \I__5629\ : InMux
    port map (
            O => \N__38209\,
            I => \foc.u_Park_Transform.n15759\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__38206\,
            I => \N__38203\
        );

    \I__5627\ : InMux
    port map (
            O => \N__38203\,
            I => \N__38200\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__38200\,
            I => \N__38197\
        );

    \I__5625\ : Span4Mux_v
    port map (
            O => \N__38197\,
            I => \N__38194\
        );

    \I__5624\ : Odrv4
    port map (
            O => \N__38194\,
            I => \foc.u_Park_Transform.Product4_mul_temp_15\
        );

    \I__5623\ : InMux
    port map (
            O => \N__38191\,
            I => \foc.u_Park_Transform.n15760\
        );

    \I__5622\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__38185\,
            I => \N__38182\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__38182\,
            I => \N__38179\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__38179\,
            I => \foc.u_Park_Transform.Product4_mul_temp_16\
        );

    \I__5618\ : InMux
    port map (
            O => \N__38176\,
            I => \foc.u_Park_Transform.n15761\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__38173\,
            I => \N__38170\
        );

    \I__5616\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38167\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__5614\ : Span4Mux_h
    port map (
            O => \N__38164\,
            I => \N__38161\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__38161\,
            I => \foc.u_Park_Transform.Product4_mul_temp_17\
        );

    \I__5612\ : InMux
    port map (
            O => \N__38158\,
            I => \foc.u_Park_Transform.n15762\
        );

    \I__5611\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38152\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__38152\,
            I => \N__38149\
        );

    \I__5609\ : Span4Mux_h
    port map (
            O => \N__38149\,
            I => \N__38146\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__38146\,
            I => \foc.u_Park_Transform.Product4_mul_temp_18\
        );

    \I__5607\ : InMux
    port map (
            O => \N__38143\,
            I => \bfn_14_19_0_\
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__38140\,
            I => \N__38137\
        );

    \I__5605\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38134\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__38134\,
            I => \N__38131\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__38131\,
            I => \N__38128\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__38128\,
            I => \foc.u_Park_Transform.Product4_mul_temp_19\
        );

    \I__5601\ : InMux
    port map (
            O => \N__38125\,
            I => \foc.u_Park_Transform.n15764\
        );

    \I__5600\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38119\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__38116\,
            I => \N__38113\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__38113\,
            I => \foc.u_Park_Transform.Product4_mul_temp_20\
        );

    \I__5596\ : InMux
    port map (
            O => \N__38110\,
            I => \foc.u_Park_Transform.n15765\
        );

    \I__5595\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38101\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__38101\,
            I => \foc.u_Park_Transform.Product4_mul_temp_4\
        );

    \I__5592\ : InMux
    port map (
            O => \N__38098\,
            I => \foc.u_Park_Transform.n15749\
        );

    \I__5591\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38092\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__38092\,
            I => \N__38089\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__38089\,
            I => \foc.u_Park_Transform.Product4_mul_temp_5\
        );

    \I__5588\ : InMux
    port map (
            O => \N__38086\,
            I => \foc.u_Park_Transform.n15750\
        );

    \I__5587\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38080\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__38077\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__38077\,
            I => \foc.u_Park_Transform.Product4_mul_temp_6\
        );

    \I__5584\ : InMux
    port map (
            O => \N__38074\,
            I => \foc.u_Park_Transform.n15751\
        );

    \I__5583\ : InMux
    port map (
            O => \N__38071\,
            I => \N__38068\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__38068\,
            I => \N__38065\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__38065\,
            I => \foc.u_Park_Transform.Product4_mul_temp_7\
        );

    \I__5580\ : InMux
    port map (
            O => \N__38062\,
            I => \foc.u_Park_Transform.n15752\
        );

    \I__5579\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38056\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__38056\,
            I => \N__38053\
        );

    \I__5577\ : Odrv12
    port map (
            O => \N__38053\,
            I => \foc.u_Park_Transform.Product4_mul_temp_8\
        );

    \I__5576\ : InMux
    port map (
            O => \N__38050\,
            I => \foc.u_Park_Transform.n15753\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__38047\,
            I => \N__38044\
        );

    \I__5574\ : InMux
    port map (
            O => \N__38044\,
            I => \N__38041\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__38041\,
            I => \foc.u_Park_Transform.Product4_mul_temp_9\
        );

    \I__5572\ : InMux
    port map (
            O => \N__38038\,
            I => \foc.u_Park_Transform.n15754\
        );

    \I__5571\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38032\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__38032\,
            I => \N__38029\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__38029\,
            I => \foc.u_Park_Transform.Product4_mul_temp_10\
        );

    \I__5568\ : InMux
    port map (
            O => \N__38026\,
            I => \bfn_14_18_0_\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__38023\,
            I => \N__38020\
        );

    \I__5566\ : InMux
    port map (
            O => \N__38020\,
            I => \N__38017\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__38017\,
            I => \N__38014\
        );

    \I__5564\ : Odrv12
    port map (
            O => \N__38014\,
            I => \foc.u_Park_Transform.Product4_mul_temp_11\
        );

    \I__5563\ : InMux
    port map (
            O => \N__38011\,
            I => \foc.u_Park_Transform.n15756\
        );

    \I__5562\ : InMux
    port map (
            O => \N__38008\,
            I => \foc.u_Park_Transform.n17076\
        );

    \I__5561\ : InMux
    port map (
            O => \N__38005\,
            I => \foc.u_Park_Transform.n17077\
        );

    \I__5560\ : InMux
    port map (
            O => \N__38002\,
            I => \foc.u_Park_Transform.n17078\
        );

    \I__5559\ : InMux
    port map (
            O => \N__37999\,
            I => \foc.u_Park_Transform.n17079\
        );

    \I__5558\ : InMux
    port map (
            O => \N__37996\,
            I => \foc.u_Park_Transform.n17080\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__37993\,
            I => \N__37990\
        );

    \I__5556\ : InMux
    port map (
            O => \N__37990\,
            I => \N__37986\
        );

    \I__5555\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37983\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37978\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37978\
        );

    \I__5552\ : Span4Mux_v
    port map (
            O => \N__37978\,
            I => \N__37975\
        );

    \I__5551\ : Odrv4
    port map (
            O => \N__37975\,
            I => \foc.u_Park_Transform.n738_adj_2003\
        );

    \I__5550\ : InMux
    port map (
            O => \N__37972\,
            I => \foc.u_Park_Transform.n17081\
        );

    \I__5549\ : InMux
    port map (
            O => \N__37969\,
            I => \foc.u_Park_Transform.n739_adj_2006\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__5547\ : InMux
    port map (
            O => \N__37963\,
            I => \N__37960\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__37960\,
            I => \N__37957\
        );

    \I__5545\ : Span4Mux_v
    port map (
            O => \N__37957\,
            I => \N__37954\
        );

    \I__5544\ : Odrv4
    port map (
            O => \N__37954\,
            I => \foc.u_Park_Transform.n739_adj_2006_THRU_CO\
        );

    \I__5543\ : InMux
    port map (
            O => \N__37951\,
            I => \N__37948\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__37948\,
            I => \N__37945\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__37945\,
            I => \foc.u_Park_Transform.Product4_mul_temp_2\
        );

    \I__5540\ : InMux
    port map (
            O => \N__37942\,
            I => \bfn_14_17_0_\
        );

    \I__5539\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37936\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__37936\,
            I => \N__37933\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__37933\,
            I => \foc.u_Park_Transform.Product4_mul_temp_3\
        );

    \I__5536\ : InMux
    port map (
            O => \N__37930\,
            I => \foc.u_Park_Transform.n15748\
        );

    \I__5535\ : InMux
    port map (
            O => \N__37927\,
            I => \foc.u_Park_Transform.n17068\
        );

    \I__5534\ : InMux
    port map (
            O => \N__37924\,
            I => \foc.u_Park_Transform.n17069\
        );

    \I__5533\ : InMux
    port map (
            O => \N__37921\,
            I => \foc.u_Park_Transform.n17070\
        );

    \I__5532\ : InMux
    port map (
            O => \N__37918\,
            I => \foc.u_Park_Transform.n17071\
        );

    \I__5531\ : InMux
    port map (
            O => \N__37915\,
            I => \foc.u_Park_Transform.n17072\
        );

    \I__5530\ : InMux
    port map (
            O => \N__37912\,
            I => \foc.u_Park_Transform.n17073\
        );

    \I__5529\ : InMux
    port map (
            O => \N__37909\,
            I => \foc.u_Park_Transform.n17074\
        );

    \I__5528\ : InMux
    port map (
            O => \N__37906\,
            I => \bfn_14_16_0_\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__37903\,
            I => \N__37900\
        );

    \I__5526\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37897\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__37897\,
            I => \foc.u_Park_Transform.n409_adj_1997\
        );

    \I__5524\ : InMux
    port map (
            O => \N__37894\,
            I => \bfn_14_14_0_\
        );

    \I__5523\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37888\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__37888\,
            I => \foc.u_Park_Transform.n458_adj_2093\
        );

    \I__5521\ : InMux
    port map (
            O => \N__37885\,
            I => \foc.u_Park_Transform.n17016\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__5519\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37876\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__37876\,
            I => \foc.u_Park_Transform.n507\
        );

    \I__5517\ : InMux
    port map (
            O => \N__37873\,
            I => \foc.u_Park_Transform.n17017\
        );

    \I__5516\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37867\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__37867\,
            I => \foc.u_Park_Transform.n556\
        );

    \I__5514\ : InMux
    port map (
            O => \N__37864\,
            I => \foc.u_Park_Transform.n17018\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__37861\,
            I => \N__37858\
        );

    \I__5512\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37855\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__37855\,
            I => \foc.u_Park_Transform.n605\
        );

    \I__5510\ : InMux
    port map (
            O => \N__37852\,
            I => \foc.u_Park_Transform.n17019\
        );

    \I__5509\ : InMux
    port map (
            O => \N__37849\,
            I => \N__37846\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__37846\,
            I => \foc.u_Park_Transform.n654\
        );

    \I__5507\ : InMux
    port map (
            O => \N__37843\,
            I => \foc.u_Park_Transform.n17020\
        );

    \I__5506\ : InMux
    port map (
            O => \N__37840\,
            I => \N__37837\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__37837\,
            I => \N__37834\
        );

    \I__5504\ : Span4Mux_v
    port map (
            O => \N__37834\,
            I => \N__37830\
        );

    \I__5503\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37827\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__37830\,
            I => \foc.u_Park_Transform.n753\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__37827\,
            I => \foc.u_Park_Transform.n753\
        );

    \I__5500\ : CascadeMux
    port map (
            O => \N__37822\,
            I => \N__37819\
        );

    \I__5499\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37816\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__37816\,
            I => \foc.u_Park_Transform.n703\
        );

    \I__5497\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37810\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__37810\,
            I => \N__37807\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__37807\,
            I => \N__37804\
        );

    \I__5494\ : Odrv4
    port map (
            O => \N__37804\,
            I => \foc.u_Park_Transform.n754\
        );

    \I__5493\ : InMux
    port map (
            O => \N__37801\,
            I => \foc.u_Park_Transform.n17021\
        );

    \I__5492\ : InMux
    port map (
            O => \N__37798\,
            I => \foc.u_Park_Transform.n755\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__5490\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37789\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__37789\,
            I => \N__37786\
        );

    \I__5488\ : Span4Mux_h
    port map (
            O => \N__37786\,
            I => \N__37783\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__37783\,
            I => \foc.u_Park_Transform.n755_THRU_CO\
        );

    \I__5486\ : InMux
    port map (
            O => \N__37780\,
            I => \foc.u_Park_Transform.n747\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__37777\,
            I => \N__37774\
        );

    \I__5484\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37771\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__37771\,
            I => \N__37768\
        );

    \I__5482\ : Span4Mux_v
    port map (
            O => \N__37768\,
            I => \N__37765\
        );

    \I__5481\ : Odrv4
    port map (
            O => \N__37765\,
            I => \foc.u_Park_Transform.n747_THRU_CO\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__37762\,
            I => \N__37746\
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__37761\,
            I => \N__37742\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__37760\,
            I => \N__37738\
        );

    \I__5477\ : CascadeMux
    port map (
            O => \N__37759\,
            I => \N__37733\
        );

    \I__5476\ : CascadeMux
    port map (
            O => \N__37758\,
            I => \N__37730\
        );

    \I__5475\ : CascadeMux
    port map (
            O => \N__37757\,
            I => \N__37726\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__37756\,
            I => \N__37722\
        );

    \I__5473\ : CascadeMux
    port map (
            O => \N__37755\,
            I => \N__37717\
        );

    \I__5472\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37710\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__37753\,
            I => \N__37707\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__37752\,
            I => \N__37704\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__37751\,
            I => \N__37701\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__37750\,
            I => \N__37697\
        );

    \I__5467\ : InMux
    port map (
            O => \N__37749\,
            I => \N__37693\
        );

    \I__5466\ : InMux
    port map (
            O => \N__37746\,
            I => \N__37680\
        );

    \I__5465\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37680\
        );

    \I__5464\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37680\
        );

    \I__5463\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37680\
        );

    \I__5462\ : InMux
    port map (
            O => \N__37738\,
            I => \N__37680\
        );

    \I__5461\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37680\
        );

    \I__5460\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37675\
        );

    \I__5459\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37675\
        );

    \I__5458\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37662\
        );

    \I__5457\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37662\
        );

    \I__5456\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37662\
        );

    \I__5455\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37662\
        );

    \I__5454\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37662\
        );

    \I__5453\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37662\
        );

    \I__5452\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37657\
        );

    \I__5451\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37657\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__37716\,
            I => \N__37654\
        );

    \I__5449\ : CascadeMux
    port map (
            O => \N__37715\,
            I => \N__37651\
        );

    \I__5448\ : CascadeMux
    port map (
            O => \N__37714\,
            I => \N__37648\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__37713\,
            I => \N__37644\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__37710\,
            I => \N__37640\
        );

    \I__5445\ : InMux
    port map (
            O => \N__37707\,
            I => \N__37637\
        );

    \I__5444\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37626\
        );

    \I__5443\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37626\
        );

    \I__5442\ : InMux
    port map (
            O => \N__37700\,
            I => \N__37626\
        );

    \I__5441\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37626\
        );

    \I__5440\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37626\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__37693\,
            I => \N__37623\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__37680\,
            I => \N__37618\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__37675\,
            I => \N__37618\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__37662\,
            I => \N__37613\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__37657\,
            I => \N__37613\
        );

    \I__5434\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37610\
        );

    \I__5433\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37599\
        );

    \I__5432\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37599\
        );

    \I__5431\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37599\
        );

    \I__5430\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37599\
        );

    \I__5429\ : InMux
    port map (
            O => \N__37643\,
            I => \N__37599\
        );

    \I__5428\ : Odrv4
    port map (
            O => \N__37640\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__37637\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__37626\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__37623\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5424\ : Odrv12
    port map (
            O => \N__37618\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__37613\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__37610\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__37599\,
            I => \foc.u_Park_Transform.n604\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__37582\,
            I => \N__37579\
        );

    \I__5419\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37576\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__37576\,
            I => \foc.u_Park_Transform.n66_adj_2033\
        );

    \I__5417\ : InMux
    port map (
            O => \N__37573\,
            I => \foc.u_Park_Transform.n17008\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__37570\,
            I => \N__37567\
        );

    \I__5415\ : InMux
    port map (
            O => \N__37567\,
            I => \N__37564\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__37564\,
            I => \foc.u_Park_Transform.n115_adj_2028\
        );

    \I__5413\ : InMux
    port map (
            O => \N__37561\,
            I => \foc.u_Park_Transform.n17009\
        );

    \I__5412\ : InMux
    port map (
            O => \N__37558\,
            I => \N__37555\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__37555\,
            I => \foc.u_Park_Transform.n164_adj_2014\
        );

    \I__5410\ : InMux
    port map (
            O => \N__37552\,
            I => \foc.u_Park_Transform.n17010\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__37549\,
            I => \N__37546\
        );

    \I__5408\ : InMux
    port map (
            O => \N__37546\,
            I => \N__37543\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__37543\,
            I => \foc.u_Park_Transform.n213_adj_1999\
        );

    \I__5406\ : InMux
    port map (
            O => \N__37540\,
            I => \foc.u_Park_Transform.n17011\
        );

    \I__5405\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37534\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__37534\,
            I => \foc.u_Park_Transform.n262\
        );

    \I__5403\ : InMux
    port map (
            O => \N__37531\,
            I => \foc.u_Park_Transform.n17012\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__37528\,
            I => \N__37525\
        );

    \I__5401\ : InMux
    port map (
            O => \N__37525\,
            I => \N__37522\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__37522\,
            I => \foc.u_Park_Transform.n311_adj_2022\
        );

    \I__5399\ : InMux
    port map (
            O => \N__37519\,
            I => \foc.u_Park_Transform.n17013\
        );

    \I__5398\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37513\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__37513\,
            I => \foc.u_Park_Transform.n360_adj_2009\
        );

    \I__5396\ : InMux
    port map (
            O => \N__37510\,
            I => \foc.u_Park_Transform.n17014\
        );

    \I__5395\ : InMux
    port map (
            O => \N__37507\,
            I => \foc.u_Park_Transform.n17226\
        );

    \I__5394\ : InMux
    port map (
            O => \N__37504\,
            I => \foc.u_Park_Transform.n17227\
        );

    \I__5393\ : InMux
    port map (
            O => \N__37501\,
            I => \bfn_14_12_0_\
        );

    \I__5392\ : InMux
    port map (
            O => \N__37498\,
            I => \foc.u_Park_Transform.n17229\
        );

    \I__5391\ : InMux
    port map (
            O => \N__37495\,
            I => \foc.u_Park_Transform.n17230\
        );

    \I__5390\ : InMux
    port map (
            O => \N__37492\,
            I => \foc.u_Park_Transform.n17231\
        );

    \I__5389\ : InMux
    port map (
            O => \N__37489\,
            I => \foc.u_Park_Transform.n17232\
        );

    \I__5388\ : InMux
    port map (
            O => \N__37486\,
            I => \foc.u_Park_Transform.n17233\
        );

    \I__5387\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37480\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__37480\,
            I => \N__37477\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__37477\,
            I => \N__37474\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__37474\,
            I => \foc.u_Park_Transform.n746\
        );

    \I__5383\ : InMux
    port map (
            O => \N__37471\,
            I => \foc.u_Park_Transform.n17234\
        );

    \I__5382\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37465\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__37465\,
            I => \foc.dCurrent_29\
        );

    \I__5380\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37459\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__37459\,
            I => \foc.dCurrent_28\
        );

    \I__5378\ : InMux
    port map (
            O => \N__37456\,
            I => \N__37453\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__37453\,
            I => \foc.dCurrent_30\
        );

    \I__5376\ : InMux
    port map (
            O => \N__37450\,
            I => \foc.u_Park_Transform.n17221\
        );

    \I__5375\ : InMux
    port map (
            O => \N__37447\,
            I => \foc.u_Park_Transform.n17222\
        );

    \I__5374\ : InMux
    port map (
            O => \N__37444\,
            I => \foc.u_Park_Transform.n17223\
        );

    \I__5373\ : InMux
    port map (
            O => \N__37441\,
            I => \foc.u_Park_Transform.n17224\
        );

    \I__5372\ : InMux
    port map (
            O => \N__37438\,
            I => \foc.u_Park_Transform.n17225\
        );

    \I__5371\ : InMux
    port map (
            O => \N__37435\,
            I => \N__37432\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__37432\,
            I => \foc.u_Park_Transform.Product1_mul_temp_23\
        );

    \I__5369\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37426\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__37426\,
            I => \N__37423\
        );

    \I__5367\ : Odrv12
    port map (
            O => \N__37423\,
            I => \foc.dCurrent_25\
        );

    \I__5366\ : InMux
    port map (
            O => \N__37420\,
            I => \foc.u_Park_Transform.n17297\
        );

    \I__5365\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37414\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__37414\,
            I => \foc.u_Park_Transform.Product1_mul_temp_24\
        );

    \I__5363\ : InMux
    port map (
            O => \N__37411\,
            I => \foc.u_Park_Transform.n17298\
        );

    \I__5362\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37405\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__37405\,
            I => \foc.u_Park_Transform.Product1_mul_temp_25\
        );

    \I__5360\ : InMux
    port map (
            O => \N__37402\,
            I => \foc.u_Park_Transform.n17299\
        );

    \I__5359\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37396\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__37396\,
            I => \foc.u_Park_Transform.Product1_mul_temp_26\
        );

    \I__5357\ : InMux
    port map (
            O => \N__37393\,
            I => \bfn_14_10_0_\
        );

    \I__5356\ : InMux
    port map (
            O => \N__37390\,
            I => \N__37387\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__37387\,
            I => \foc.u_Park_Transform.Product1_mul_temp_27\
        );

    \I__5354\ : InMux
    port map (
            O => \N__37384\,
            I => \foc.u_Park_Transform.n17301\
        );

    \I__5353\ : InMux
    port map (
            O => \N__37381\,
            I => \N__37378\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__37378\,
            I => \foc.u_Park_Transform.Product1_mul_temp_28\
        );

    \I__5351\ : InMux
    port map (
            O => \N__37375\,
            I => \foc.u_Park_Transform.n17302\
        );

    \I__5350\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37369\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__37369\,
            I => \foc.u_Park_Transform.Product1_mul_temp_29\
        );

    \I__5348\ : InMux
    port map (
            O => \N__37366\,
            I => \foc.u_Park_Transform.n17303\
        );

    \I__5347\ : CascadeMux
    port map (
            O => \N__37363\,
            I => \foc.dCurrent_31_cascade_\
        );

    \I__5346\ : InMux
    port map (
            O => \N__37360\,
            I => \N__37357\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__37357\,
            I => \foc.u_Park_Transform.Product1_mul_temp_15\
        );

    \I__5344\ : InMux
    port map (
            O => \N__37354\,
            I => \N__37351\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__37351\,
            I => \N__37348\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__37348\,
            I => \foc.dCurrent_17\
        );

    \I__5341\ : InMux
    port map (
            O => \N__37345\,
            I => \foc.u_Park_Transform.n17289\
        );

    \I__5340\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37339\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__37339\,
            I => \foc.u_Park_Transform.Product1_mul_temp_16\
        );

    \I__5338\ : InMux
    port map (
            O => \N__37336\,
            I => \N__37333\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__37333\,
            I => \N__37330\
        );

    \I__5336\ : Odrv12
    port map (
            O => \N__37330\,
            I => \foc.dCurrent_18\
        );

    \I__5335\ : InMux
    port map (
            O => \N__37327\,
            I => \foc.u_Park_Transform.n17290\
        );

    \I__5334\ : InMux
    port map (
            O => \N__37324\,
            I => \N__37321\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__37321\,
            I => \foc.u_Park_Transform.Product1_mul_temp_17\
        );

    \I__5332\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37315\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__37315\,
            I => \N__37312\
        );

    \I__5330\ : Odrv4
    port map (
            O => \N__37312\,
            I => \foc.dCurrent_19\
        );

    \I__5329\ : InMux
    port map (
            O => \N__37309\,
            I => \foc.u_Park_Transform.n17291\
        );

    \I__5328\ : InMux
    port map (
            O => \N__37306\,
            I => \N__37303\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__37303\,
            I => \foc.u_Park_Transform.Product1_mul_temp_18\
        );

    \I__5326\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37297\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__37297\,
            I => \N__37294\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__37294\,
            I => \foc.dCurrent_20\
        );

    \I__5323\ : InMux
    port map (
            O => \N__37291\,
            I => \bfn_14_9_0_\
        );

    \I__5322\ : InMux
    port map (
            O => \N__37288\,
            I => \N__37285\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__37285\,
            I => \foc.u_Park_Transform.Product1_mul_temp_19\
        );

    \I__5320\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37279\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__37279\,
            I => \N__37276\
        );

    \I__5318\ : Odrv4
    port map (
            O => \N__37276\,
            I => \foc.dCurrent_21\
        );

    \I__5317\ : InMux
    port map (
            O => \N__37273\,
            I => \foc.u_Park_Transform.n17293\
        );

    \I__5316\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37267\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__37267\,
            I => \foc.u_Park_Transform.Product1_mul_temp_20\
        );

    \I__5314\ : InMux
    port map (
            O => \N__37264\,
            I => \N__37261\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__37261\,
            I => \N__37258\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__37258\,
            I => \foc.dCurrent_22\
        );

    \I__5311\ : InMux
    port map (
            O => \N__37255\,
            I => \foc.u_Park_Transform.n17294\
        );

    \I__5310\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37249\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__37249\,
            I => \foc.u_Park_Transform.Product1_mul_temp_21\
        );

    \I__5308\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37243\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37240\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__37240\,
            I => \foc.dCurrent_23\
        );

    \I__5305\ : InMux
    port map (
            O => \N__37237\,
            I => \foc.u_Park_Transform.n17295\
        );

    \I__5304\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37231\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__37231\,
            I => \foc.u_Park_Transform.Product1_mul_temp_22\
        );

    \I__5302\ : InMux
    port map (
            O => \N__37228\,
            I => \N__37225\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__37225\,
            I => \N__37222\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__37222\,
            I => \foc.dCurrent_24\
        );

    \I__5299\ : InMux
    port map (
            O => \N__37219\,
            I => \foc.u_Park_Transform.n17296\
        );

    \I__5298\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37213\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__37213\,
            I => \foc.dCurrent_9\
        );

    \I__5296\ : InMux
    port map (
            O => \N__37210\,
            I => \foc.u_Park_Transform.n17281\
        );

    \I__5295\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37204\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__37204\,
            I => \foc.dCurrent_10\
        );

    \I__5293\ : InMux
    port map (
            O => \N__37201\,
            I => \foc.u_Park_Transform.n17282\
        );

    \I__5292\ : InMux
    port map (
            O => \N__37198\,
            I => \N__37195\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__37195\,
            I => \foc.dCurrent_11\
        );

    \I__5290\ : InMux
    port map (
            O => \N__37192\,
            I => \foc.u_Park_Transform.n17283\
        );

    \I__5289\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37186\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__37186\,
            I => \N__37183\
        );

    \I__5287\ : Odrv12
    port map (
            O => \N__37183\,
            I => \foc.dCurrent_12\
        );

    \I__5286\ : InMux
    port map (
            O => \N__37180\,
            I => \bfn_14_8_0_\
        );

    \I__5285\ : InMux
    port map (
            O => \N__37177\,
            I => \N__37174\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__37174\,
            I => \N__37171\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__37171\,
            I => \foc.dCurrent_13\
        );

    \I__5282\ : InMux
    port map (
            O => \N__37168\,
            I => \foc.u_Park_Transform.n17285\
        );

    \I__5281\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37162\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__37162\,
            I => \N__37159\
        );

    \I__5279\ : Odrv12
    port map (
            O => \N__37159\,
            I => \foc.dCurrent_14\
        );

    \I__5278\ : InMux
    port map (
            O => \N__37156\,
            I => \foc.u_Park_Transform.n17286\
        );

    \I__5277\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37150\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__37150\,
            I => \N__37147\
        );

    \I__5275\ : Odrv12
    port map (
            O => \N__37147\,
            I => \foc.dCurrent_15\
        );

    \I__5274\ : InMux
    port map (
            O => \N__37144\,
            I => \foc.u_Park_Transform.n17287\
        );

    \I__5273\ : InMux
    port map (
            O => \N__37141\,
            I => \N__37138\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__37138\,
            I => \N__37135\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__37135\,
            I => \foc.dCurrent_16\
        );

    \I__5270\ : InMux
    port map (
            O => \N__37132\,
            I => \foc.u_Park_Transform.n17288\
        );

    \I__5269\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37126\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__37126\,
            I => \N__37123\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__37123\,
            I => \foc.dCurrent_4\
        );

    \I__5266\ : InMux
    port map (
            O => \N__37120\,
            I => \N__37117\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__37117\,
            I => \N__37114\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__37114\,
            I => \foc.dCurrent_5\
        );

    \I__5263\ : InMux
    port map (
            O => \N__37111\,
            I => \foc.u_Park_Transform.n17277\
        );

    \I__5262\ : InMux
    port map (
            O => \N__37108\,
            I => \N__37105\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__37105\,
            I => \N__37102\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__37102\,
            I => \foc.dCurrent_6\
        );

    \I__5259\ : InMux
    port map (
            O => \N__37099\,
            I => \foc.u_Park_Transform.n17278\
        );

    \I__5258\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37093\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__37093\,
            I => \N__37090\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__37090\,
            I => \foc.dCurrent_7\
        );

    \I__5255\ : InMux
    port map (
            O => \N__37087\,
            I => \foc.u_Park_Transform.n17279\
        );

    \I__5254\ : InMux
    port map (
            O => \N__37084\,
            I => \N__37081\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__37081\,
            I => \N__37078\
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__37078\,
            I => \foc.dCurrent_8\
        );

    \I__5251\ : InMux
    port map (
            O => \N__37075\,
            I => \foc.u_Park_Transform.n17280\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__37072\,
            I => \N__37069\
        );

    \I__5249\ : InMux
    port map (
            O => \N__37069\,
            I => \N__37066\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__37066\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n467_adj_604\
        );

    \I__5247\ : InMux
    port map (
            O => \N__37063\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18100\
        );

    \I__5246\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37057\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__37057\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n516_adj_603\
        );

    \I__5244\ : InMux
    port map (
            O => \N__37054\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18101\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__37051\,
            I => \N__37048\
        );

    \I__5242\ : InMux
    port map (
            O => \N__37048\,
            I => \N__37045\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__37045\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n565_adj_602\
        );

    \I__5240\ : InMux
    port map (
            O => \N__37042\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18102\
        );

    \I__5239\ : InMux
    port map (
            O => \N__37039\,
            I => \N__37036\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__37036\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n614_adj_601\
        );

    \I__5237\ : InMux
    port map (
            O => \N__37033\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18103\
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__37030\,
            I => \N__37027\
        );

    \I__5235\ : InMux
    port map (
            O => \N__37027\,
            I => \N__37024\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__37024\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n663_adj_600\
        );

    \I__5233\ : InMux
    port map (
            O => \N__37021\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18104\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__5231\ : InMux
    port map (
            O => \N__37015\,
            I => \N__37012\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__37012\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n712_adj_599\
        );

    \I__5229\ : InMux
    port map (
            O => \N__37009\,
            I => \N__37006\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__37006\,
            I => \N__37003\
        );

    \I__5227\ : Odrv12
    port map (
            O => \N__37003\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n766_adj_619\
        );

    \I__5226\ : InMux
    port map (
            O => \N__37000\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18105\
        );

    \I__5225\ : InMux
    port map (
            O => \N__36997\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620\
        );

    \I__5224\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36991\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__36991\,
            I => \N__36988\
        );

    \I__5222\ : Odrv12
    port map (
            O => \N__36988\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_CO\
        );

    \I__5221\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36982\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__36982\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n75_adj_618\
        );

    \I__5219\ : InMux
    port map (
            O => \N__36979\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18092\
        );

    \I__5218\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36973\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__36973\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n124_adj_616\
        );

    \I__5216\ : InMux
    port map (
            O => \N__36970\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18093\
        );

    \I__5215\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36964\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__36964\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n173_adj_614\
        );

    \I__5213\ : InMux
    port map (
            O => \N__36961\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18094\
        );

    \I__5212\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36955\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__36955\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n222_adj_612\
        );

    \I__5210\ : InMux
    port map (
            O => \N__36952\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18095\
        );

    \I__5209\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36946\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__36946\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n271_adj_610\
        );

    \I__5207\ : InMux
    port map (
            O => \N__36943\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18096\
        );

    \I__5206\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36937\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__36937\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n320_adj_608\
        );

    \I__5204\ : InMux
    port map (
            O => \N__36934\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18097\
        );

    \I__5203\ : InMux
    port map (
            O => \N__36931\,
            I => \N__36928\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__36928\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n369_adj_606\
        );

    \I__5201\ : InMux
    port map (
            O => \N__36925\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18098\
        );

    \I__5200\ : InMux
    port map (
            O => \N__36922\,
            I => \N__36919\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__36919\,
            I => \N__36916\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__36916\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n418_adj_605\
        );

    \I__5197\ : InMux
    port map (
            O => \N__36913\,
            I => \bfn_13_26_0_\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__36910\,
            I => \N__36907\
        );

    \I__5195\ : InMux
    port map (
            O => \N__36907\,
            I => \N__36904\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__36904\,
            I => \N__36901\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__36901\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n770_adj_597\
        );

    \I__5192\ : InMux
    port map (
            O => \N__36898\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17965\
        );

    \I__5191\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36892\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__36892\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n774\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__36889\,
            I => \N__36886\
        );

    \I__5188\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36883\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__36883\,
            I => \N__36880\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__36880\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_CO\
        );

    \I__5185\ : InMux
    port map (
            O => \N__36877\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17966\
        );

    \I__5184\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36871\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36868\
        );

    \I__5182\ : Odrv12
    port map (
            O => \N__36868\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n778_adj_737\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__36865\,
            I => \N__36862\
        );

    \I__5180\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36859\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__36859\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_CO\
        );

    \I__5178\ : InMux
    port map (
            O => \N__36856\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17967\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__36853\,
            I => \N__36850\
        );

    \I__5176\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36847\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__36847\,
            I => \N__36844\
        );

    \I__5174\ : Odrv12
    port map (
            O => \N__36844\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_CO\
        );

    \I__5173\ : InMux
    port map (
            O => \N__36841\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17968\
        );

    \I__5172\ : InMux
    port map (
            O => \N__36838\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17969\
        );

    \I__5171\ : InMux
    port map (
            O => \N__36835\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17970\
        );

    \I__5170\ : InMux
    port map (
            O => \N__36832\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17971\
        );

    \I__5169\ : InMux
    port map (
            O => \N__36829\,
            I => \bfn_13_24_0_\
        );

    \I__5168\ : InMux
    port map (
            O => \N__36826\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17957\
        );

    \I__5167\ : InMux
    port map (
            O => \N__36823\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17958\
        );

    \I__5166\ : InMux
    port map (
            O => \N__36820\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17959\
        );

    \I__5165\ : InMux
    port map (
            O => \N__36817\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17960\
        );

    \I__5164\ : InMux
    port map (
            O => \N__36814\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17961\
        );

    \I__5163\ : InMux
    port map (
            O => \N__36811\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17962\
        );

    \I__5162\ : InMux
    port map (
            O => \N__36808\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17963\
        );

    \I__5161\ : InMux
    port map (
            O => \N__36805\,
            I => \bfn_13_23_0_\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__36802\,
            I => \N__36799\
        );

    \I__5159\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36796\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__36796\,
            I => \N__36793\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__36793\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n228_adj_742\
        );

    \I__5156\ : InMux
    port map (
            O => \N__36790\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17858\
        );

    \I__5155\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36784\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36781\
        );

    \I__5153\ : Span4Mux_h
    port map (
            O => \N__36781\,
            I => \N__36778\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__36778\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n277_adj_741\
        );

    \I__5151\ : InMux
    port map (
            O => \N__36775\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17859\
        );

    \I__5150\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36769\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__36769\,
            I => \N__36766\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__36766\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n326\
        );

    \I__5147\ : InMux
    port map (
            O => \N__36763\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17860\
        );

    \I__5146\ : InMux
    port map (
            O => \N__36760\,
            I => \N__36757\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__36757\,
            I => \N__36754\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__36754\,
            I => \N__36751\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__36751\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n375\
        );

    \I__5142\ : InMux
    port map (
            O => \N__36748\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17861\
        );

    \I__5141\ : InMux
    port map (
            O => \N__36745\,
            I => \N__36742\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__36742\,
            I => \N__36739\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__36739\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n424\
        );

    \I__5138\ : InMux
    port map (
            O => \N__36736\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17862\
        );

    \I__5137\ : InMux
    port map (
            O => \N__36733\,
            I => \N__36730\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__36730\,
            I => \N__36727\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__36727\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n473\
        );

    \I__5134\ : InMux
    port map (
            O => \N__36724\,
            I => \bfn_13_21_0_\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__36721\,
            I => \N__36717\
        );

    \I__5132\ : CascadeMux
    port map (
            O => \N__36720\,
            I => \N__36713\
        );

    \I__5131\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36706\
        );

    \I__5130\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36706\
        );

    \I__5129\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36706\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__36706\,
            I => \N__36703\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__36703\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n522\
        );

    \I__5126\ : InMux
    port map (
            O => \N__36700\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17864\
        );

    \I__5125\ : InMux
    port map (
            O => \N__36697\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17865\
        );

    \I__5124\ : InMux
    port map (
            O => \N__36694\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736\
        );

    \I__5123\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36688\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__36688\,
            I => \N__36685\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__36685\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3014\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__36682\,
            I => \N__36675\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__36681\,
            I => \N__36672\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__36680\,
            I => \N__36669\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__36679\,
            I => \N__36666\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__36678\,
            I => \N__36662\
        );

    \I__5115\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36655\
        );

    \I__5114\ : InMux
    port map (
            O => \N__36672\,
            I => \N__36655\
        );

    \I__5113\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36644\
        );

    \I__5112\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36644\
        );

    \I__5111\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36644\
        );

    \I__5110\ : InMux
    port map (
            O => \N__36662\,
            I => \N__36644\
        );

    \I__5109\ : InMux
    port map (
            O => \N__36661\,
            I => \N__36644\
        );

    \I__5108\ : InMux
    port map (
            O => \N__36660\,
            I => \N__36641\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__36655\,
            I => \N__36636\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__36644\,
            I => \N__36636\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__36641\,
            I => \N__36633\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__36636\,
            I => \N__36630\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__36633\,
            I => \N__36627\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__36630\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__36627\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810\
        );

    \I__5100\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36619\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__36619\,
            I => \N__36616\
        );

    \I__5098\ : Span4Mux_h
    port map (
            O => \N__36616\,
            I => \N__36613\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__36613\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3111\
        );

    \I__5096\ : InMux
    port map (
            O => \N__36610\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373\
        );

    \I__5095\ : InMux
    port map (
            O => \N__36607\,
            I => \N__36604\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__36604\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3114\
        );

    \I__5093\ : InMux
    port map (
            O => \N__36601\,
            I => \N__36598\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__36598\,
            I => \N__36595\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__36595\,
            I => \N__36592\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__36592\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3215\
        );

    \I__5089\ : InMux
    port map (
            O => \N__36589\,
            I => \bfn_13_18_0_\
        );

    \I__5088\ : InMux
    port map (
            O => \N__36586\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__36583\,
            I => \N__36580\
        );

    \I__5086\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36577\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36574\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__36574\,
            I => \N__36571\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__36571\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_CO\
        );

    \I__5082\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36562\
        );

    \I__5081\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36562\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__36562\,
            I => \N__36558\
        );

    \I__5079\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36555\
        );

    \I__5078\ : Span4Mux_v
    port map (
            O => \N__36558\,
            I => \N__36550\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__36555\,
            I => \N__36550\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__36550\,
            I => \N__36547\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__36547\,
            I => \foc.Look_Up_Table_out1_1_0\
        );

    \I__5074\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36541\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__36541\,
            I => \N__36538\
        );

    \I__5072\ : Span12Mux_v
    port map (
            O => \N__36538\,
            I => \N__36534\
        );

    \I__5071\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36531\
        );

    \I__5070\ : Odrv12
    port map (
            O => \N__36534\,
            I => n794
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__36531\,
            I => n794
        );

    \I__5068\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36523\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__36523\,
            I => \N__36520\
        );

    \I__5066\ : Odrv4
    port map (
            O => \N__36520\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n81_adj_750\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__36517\,
            I => \N__36514\
        );

    \I__5064\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36511\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36508\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__36508\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n130_adj_748\
        );

    \I__5061\ : InMux
    port map (
            O => \N__36505\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17856\
        );

    \I__5060\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36499\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__36499\,
            I => \N__36496\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__36496\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n179_adj_746\
        );

    \I__5057\ : InMux
    port map (
            O => \N__36493\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17857\
        );

    \I__5056\ : InMux
    port map (
            O => \N__36490\,
            I => \foc.u_Park_Transform.n763_adj_2054\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__36487\,
            I => \N__36484\
        );

    \I__5054\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36481\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__36481\,
            I => \N__36478\
        );

    \I__5052\ : Span4Mux_v
    port map (
            O => \N__36478\,
            I => \N__36475\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__36475\,
            I => \foc.u_Park_Transform.n763_adj_2054_THRU_CO\
        );

    \I__5050\ : InMux
    port map (
            O => \N__36472\,
            I => \N__36464\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__36471\,
            I => \N__36461\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__36470\,
            I => \N__36458\
        );

    \I__5047\ : CascadeMux
    port map (
            O => \N__36469\,
            I => \N__36455\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__36468\,
            I => \N__36452\
        );

    \I__5045\ : CascadeMux
    port map (
            O => \N__36467\,
            I => \N__36448\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__36464\,
            I => \N__36444\
        );

    \I__5043\ : InMux
    port map (
            O => \N__36461\,
            I => \N__36439\
        );

    \I__5042\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36439\
        );

    \I__5041\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36428\
        );

    \I__5040\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36428\
        );

    \I__5039\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36428\
        );

    \I__5038\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36428\
        );

    \I__5037\ : InMux
    port map (
            O => \N__36447\,
            I => \N__36428\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__36444\,
            I => \N__36425\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__36439\,
            I => \N__36420\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__36428\,
            I => \N__36420\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__36425\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813\
        );

    \I__5032\ : Odrv12
    port map (
            O => \N__36420\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__36415\,
            I => \N__36412\
        );

    \I__5030\ : InMux
    port map (
            O => \N__36412\,
            I => \N__36409\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__36409\,
            I => \N__36406\
        );

    \I__5028\ : Span4Mux_v
    port map (
            O => \N__36406\,
            I => \N__36403\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__36403\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2411\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__36400\,
            I => \N__36397\
        );

    \I__5025\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36394\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__36394\,
            I => \N__36391\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__36391\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2414\
        );

    \I__5022\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36385\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__36385\,
            I => \N__36382\
        );

    \I__5020\ : Odrv12
    port map (
            O => \N__36382\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2511\
        );

    \I__5019\ : InMux
    port map (
            O => \N__36379\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367\
        );

    \I__5018\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36373\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__36373\,
            I => \N__36370\
        );

    \I__5016\ : Span4Mux_h
    port map (
            O => \N__36370\,
            I => \N__36367\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__36367\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2514\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__36364\,
            I => \N__36361\
        );

    \I__5013\ : InMux
    port map (
            O => \N__36361\,
            I => \N__36358\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__36358\,
            I => \N__36355\
        );

    \I__5011\ : Span4Mux_h
    port map (
            O => \N__36355\,
            I => \N__36352\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__36352\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2611\
        );

    \I__5009\ : InMux
    port map (
            O => \N__36349\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__36346\,
            I => \N__36343\
        );

    \I__5007\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36340\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36337\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__36337\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2614\
        );

    \I__5004\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36331\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__36331\,
            I => \N__36328\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__36328\,
            I => \N__36325\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__36325\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2711\
        );

    \I__5000\ : InMux
    port map (
            O => \N__36322\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369\
        );

    \I__4999\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36316\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__36316\,
            I => \N__36313\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__36313\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2714\
        );

    \I__4996\ : CascadeMux
    port map (
            O => \N__36310\,
            I => \N__36307\
        );

    \I__4995\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36304\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__36304\,
            I => \N__36301\
        );

    \I__4993\ : Odrv12
    port map (
            O => \N__36301\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2811\
        );

    \I__4992\ : InMux
    port map (
            O => \N__36298\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370\
        );

    \I__4991\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36292\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__36292\,
            I => \N__36289\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__36289\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2814\
        );

    \I__4988\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36283\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__36283\,
            I => \N__36280\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__36280\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2911\
        );

    \I__4985\ : InMux
    port map (
            O => \N__36277\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371\
        );

    \I__4984\ : InMux
    port map (
            O => \N__36274\,
            I => \N__36271\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__36268\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2914\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__36265\,
            I => \N__36262\
        );

    \I__4980\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36259\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__36259\,
            I => \N__36256\
        );

    \I__4978\ : Odrv12
    port map (
            O => \N__36256\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3011\
        );

    \I__4977\ : InMux
    port map (
            O => \N__36253\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__36250\,
            I => \N__36247\
        );

    \I__4975\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36244\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__36244\,
            I => \foc.u_Park_Transform.n412_adj_1995\
        );

    \I__4973\ : InMux
    port map (
            O => \N__36241\,
            I => \foc.u_Park_Transform.n16984\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__36238\,
            I => \N__36235\
        );

    \I__4971\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36232\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__36232\,
            I => \foc.u_Park_Transform.n415\
        );

    \I__4969\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36226\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__36226\,
            I => \N__36223\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__36223\,
            I => \foc.u_Park_Transform.n461_adj_2007\
        );

    \I__4966\ : InMux
    port map (
            O => \N__36220\,
            I => \bfn_13_16_0_\
        );

    \I__4965\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36214\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__36214\,
            I => \foc.u_Park_Transform.n464\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__36211\,
            I => \N__36208\
        );

    \I__4962\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36205\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__36205\,
            I => \N__36202\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__36202\,
            I => \foc.u_Park_Transform.n510\
        );

    \I__4959\ : InMux
    port map (
            O => \N__36199\,
            I => \foc.u_Park_Transform.n16986\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36193\
        );

    \I__4957\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36190\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__36190\,
            I => \foc.u_Park_Transform.n513\
        );

    \I__4955\ : InMux
    port map (
            O => \N__36187\,
            I => \N__36184\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__36184\,
            I => \N__36181\
        );

    \I__4953\ : Odrv4
    port map (
            O => \N__36181\,
            I => \foc.u_Park_Transform.n559\
        );

    \I__4952\ : InMux
    port map (
            O => \N__36178\,
            I => \foc.u_Park_Transform.n16987\
        );

    \I__4951\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36172\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__36172\,
            I => \foc.u_Park_Transform.n562\
        );

    \I__4949\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36166\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__36166\,
            I => \N__36163\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__36163\,
            I => \foc.u_Park_Transform.n608_adj_2067\
        );

    \I__4946\ : InMux
    port map (
            O => \N__36160\,
            I => \foc.u_Park_Transform.n16988\
        );

    \I__4945\ : InMux
    port map (
            O => \N__36157\,
            I => \N__36154\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__36154\,
            I => \foc.u_Park_Transform.n611_adj_2107\
        );

    \I__4943\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36148\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__36148\,
            I => \N__36145\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__36145\,
            I => \foc.u_Park_Transform.n657_adj_2064\
        );

    \I__4940\ : InMux
    port map (
            O => \N__36142\,
            I => \foc.u_Park_Transform.n16989\
        );

    \I__4939\ : InMux
    port map (
            O => \N__36139\,
            I => \N__36136\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__36136\,
            I => \foc.u_Park_Transform.n660_adj_2091\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__36133\,
            I => \N__36121\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__36132\,
            I => \N__36118\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__36131\,
            I => \N__36115\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__36130\,
            I => \N__36112\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__36129\,
            I => \N__36108\
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__36128\,
            I => \N__36104\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__36127\,
            I => \N__36100\
        );

    \I__4930\ : CascadeMux
    port map (
            O => \N__36126\,
            I => \N__36096\
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__36125\,
            I => \N__36092\
        );

    \I__4928\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36086\
        );

    \I__4927\ : InMux
    port map (
            O => \N__36121\,
            I => \N__36086\
        );

    \I__4926\ : InMux
    port map (
            O => \N__36118\,
            I => \N__36075\
        );

    \I__4925\ : InMux
    port map (
            O => \N__36115\,
            I => \N__36064\
        );

    \I__4924\ : InMux
    port map (
            O => \N__36112\,
            I => \N__36064\
        );

    \I__4923\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36064\
        );

    \I__4922\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36064\
        );

    \I__4921\ : InMux
    port map (
            O => \N__36107\,
            I => \N__36064\
        );

    \I__4920\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36047\
        );

    \I__4919\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36047\
        );

    \I__4918\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36047\
        );

    \I__4917\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36047\
        );

    \I__4916\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36047\
        );

    \I__4915\ : InMux
    port map (
            O => \N__36095\,
            I => \N__36047\
        );

    \I__4914\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36047\
        );

    \I__4913\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36047\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__36086\,
            I => \N__36044\
        );

    \I__4911\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36041\
        );

    \I__4910\ : CascadeMux
    port map (
            O => \N__36084\,
            I => \N__36038\
        );

    \I__4909\ : CascadeMux
    port map (
            O => \N__36083\,
            I => \N__36034\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__36082\,
            I => \N__36030\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__36081\,
            I => \N__36026\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__36080\,
            I => \N__36023\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__36079\,
            I => \N__36019\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__36078\,
            I => \N__36015\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__36075\,
            I => \N__36004\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__36064\,
            I => \N__36004\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__36047\,
            I => \N__36004\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__36044\,
            I => \N__36004\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__36004\
        );

    \I__4898\ : InMux
    port map (
            O => \N__36038\,
            I => \N__35991\
        );

    \I__4897\ : InMux
    port map (
            O => \N__36037\,
            I => \N__35991\
        );

    \I__4896\ : InMux
    port map (
            O => \N__36034\,
            I => \N__35991\
        );

    \I__4895\ : InMux
    port map (
            O => \N__36033\,
            I => \N__35991\
        );

    \I__4894\ : InMux
    port map (
            O => \N__36030\,
            I => \N__35991\
        );

    \I__4893\ : InMux
    port map (
            O => \N__36029\,
            I => \N__35991\
        );

    \I__4892\ : InMux
    port map (
            O => \N__36026\,
            I => \N__35988\
        );

    \I__4891\ : InMux
    port map (
            O => \N__36023\,
            I => \N__35977\
        );

    \I__4890\ : InMux
    port map (
            O => \N__36022\,
            I => \N__35977\
        );

    \I__4889\ : InMux
    port map (
            O => \N__36019\,
            I => \N__35977\
        );

    \I__4888\ : InMux
    port map (
            O => \N__36018\,
            I => \N__35977\
        );

    \I__4887\ : InMux
    port map (
            O => \N__36015\,
            I => \N__35977\
        );

    \I__4886\ : Span4Mux_v
    port map (
            O => \N__36004\,
            I => \N__35973\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__35991\,
            I => \N__35966\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__35988\,
            I => \N__35966\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__35977\,
            I => \N__35966\
        );

    \I__4882\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35963\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__35973\,
            I => \foc.u_Park_Transform.n607\
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__35966\,
            I => \foc.u_Park_Transform.n607\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__35963\,
            I => \foc.u_Park_Transform.n607\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__35956\,
            I => \N__35953\
        );

    \I__4877\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__35950\,
            I => \N__35947\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__35947\,
            I => \foc.u_Park_Transform.n706_adj_2044\
        );

    \I__4874\ : InMux
    port map (
            O => \N__35944\,
            I => \foc.u_Park_Transform.n16990\
        );

    \I__4873\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35935\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__35935\,
            I => \N__35931\
        );

    \I__4870\ : InMux
    port map (
            O => \N__35934\,
            I => \N__35928\
        );

    \I__4869\ : Span4Mux_v
    port map (
            O => \N__35931\,
            I => \N__35923\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__35928\,
            I => \N__35923\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__35923\,
            I => \foc.u_Park_Transform.n761\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__35920\,
            I => \N__35917\
        );

    \I__4865\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35914\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__35914\,
            I => \N__35911\
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__35911\,
            I => \foc.u_Park_Transform.n709_adj_2066\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__35908\,
            I => \N__35905\
        );

    \I__4861\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35902\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__35902\,
            I => \foc.u_Park_Transform.n762_adj_2065\
        );

    \I__4859\ : InMux
    port map (
            O => \N__35899\,
            I => \foc.u_Park_Transform.n16991\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__35896\,
            I => \N__35880\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__35895\,
            I => \N__35876\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__35894\,
            I => \N__35872\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__35893\,
            I => \N__35867\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__35892\,
            I => \N__35864\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__35891\,
            I => \N__35861\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__35890\,
            I => \N__35858\
        );

    \I__4851\ : CascadeMux
    port map (
            O => \N__35889\,
            I => \N__35855\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__35888\,
            I => \N__35851\
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__35887\,
            I => \N__35847\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__35886\,
            I => \N__35843\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__35885\,
            I => \N__35839\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__35884\,
            I => \N__35835\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__35883\,
            I => \N__35832\
        );

    \I__4844\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35819\
        );

    \I__4843\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35819\
        );

    \I__4842\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35819\
        );

    \I__4841\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35819\
        );

    \I__4840\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35819\
        );

    \I__4839\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35819\
        );

    \I__4838\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35814\
        );

    \I__4837\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35814\
        );

    \I__4836\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35807\
        );

    \I__4835\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35804\
        );

    \I__4834\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35793\
        );

    \I__4833\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35793\
        );

    \I__4832\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35793\
        );

    \I__4831\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35793\
        );

    \I__4830\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35793\
        );

    \I__4829\ : InMux
    port map (
            O => \N__35847\,
            I => \N__35778\
        );

    \I__4828\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35778\
        );

    \I__4827\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35778\
        );

    \I__4826\ : InMux
    port map (
            O => \N__35842\,
            I => \N__35778\
        );

    \I__4825\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35778\
        );

    \I__4824\ : InMux
    port map (
            O => \N__35838\,
            I => \N__35778\
        );

    \I__4823\ : InMux
    port map (
            O => \N__35835\,
            I => \N__35778\
        );

    \I__4822\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35775\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__35819\,
            I => \N__35770\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35770\
        );

    \I__4819\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35767\
        );

    \I__4818\ : CascadeMux
    port map (
            O => \N__35812\,
            I => \N__35763\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__35811\,
            I => \N__35759\
        );

    \I__4816\ : CascadeMux
    port map (
            O => \N__35810\,
            I => \N__35755\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35752\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__35804\,
            I => \N__35743\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__35793\,
            I => \N__35743\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35743\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35743\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__35770\,
            I => \N__35738\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__35767\,
            I => \N__35738\
        );

    \I__4808\ : InMux
    port map (
            O => \N__35766\,
            I => \N__35725\
        );

    \I__4807\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35725\
        );

    \I__4806\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35725\
        );

    \I__4805\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35725\
        );

    \I__4804\ : InMux
    port map (
            O => \N__35758\,
            I => \N__35725\
        );

    \I__4803\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35725\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__35752\,
            I => \N__35722\
        );

    \I__4801\ : Span12Mux_v
    port map (
            O => \N__35743\,
            I => \N__35719\
        );

    \I__4800\ : Span4Mux_h
    port map (
            O => \N__35738\,
            I => \N__35714\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35714\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__35722\,
            I => \foc.u_Park_Transform.n610\
        );

    \I__4797\ : Odrv12
    port map (
            O => \N__35719\,
            I => \foc.u_Park_Transform.n610\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__35714\,
            I => \foc.u_Park_Transform.n610\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__35707\,
            I => \N__35704\
        );

    \I__4794\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35701\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35698\
        );

    \I__4792\ : Odrv12
    port map (
            O => \N__35698\,
            I => \foc.u_Park_Transform.n69_adj_2059\
        );

    \I__4791\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35692\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__35692\,
            I => \foc.u_Park_Transform.n72_adj_2062\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__35689\,
            I => \N__35686\
        );

    \I__4788\ : InMux
    port map (
            O => \N__35686\,
            I => \N__35683\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35680\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__35680\,
            I => \foc.u_Park_Transform.n118_adj_2037\
        );

    \I__4785\ : InMux
    port map (
            O => \N__35677\,
            I => \foc.u_Park_Transform.n16978\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__35674\,
            I => \N__35671\
        );

    \I__4783\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35668\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__35668\,
            I => \foc.u_Park_Transform.n121_adj_2051\
        );

    \I__4781\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35662\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__35662\,
            I => \N__35659\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__35659\,
            I => \foc.u_Park_Transform.n167_adj_2029\
        );

    \I__4778\ : InMux
    port map (
            O => \N__35656\,
            I => \foc.u_Park_Transform.n16979\
        );

    \I__4777\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35650\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__35650\,
            I => \foc.u_Park_Transform.n170_adj_2048\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__35647\,
            I => \N__35644\
        );

    \I__4774\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35641\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35638\
        );

    \I__4772\ : Odrv12
    port map (
            O => \N__35638\,
            I => \foc.u_Park_Transform.n216_adj_2025\
        );

    \I__4771\ : InMux
    port map (
            O => \N__35635\,
            I => \foc.u_Park_Transform.n16980\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__35632\,
            I => \N__35629\
        );

    \I__4769\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35626\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__35626\,
            I => \foc.u_Park_Transform.n219_adj_2040\
        );

    \I__4767\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35620\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__35620\,
            I => \N__35617\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__35617\,
            I => \foc.u_Park_Transform.n265_adj_2023\
        );

    \I__4764\ : InMux
    port map (
            O => \N__35614\,
            I => \foc.u_Park_Transform.n16981\
        );

    \I__4763\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35608\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__35608\,
            I => \foc.u_Park_Transform.n268_adj_2027\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__35605\,
            I => \N__35602\
        );

    \I__4760\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35599\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35596\
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__35596\,
            I => \foc.u_Park_Transform.n314_adj_2010\
        );

    \I__4757\ : InMux
    port map (
            O => \N__35593\,
            I => \foc.u_Park_Transform.n16982\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__35590\,
            I => \N__35587\
        );

    \I__4755\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35584\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__35584\,
            I => \foc.u_Park_Transform.n317_adj_2021\
        );

    \I__4753\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35578\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__35578\,
            I => \N__35575\
        );

    \I__4751\ : Odrv12
    port map (
            O => \N__35575\,
            I => \foc.u_Park_Transform.n363_adj_1998\
        );

    \I__4750\ : InMux
    port map (
            O => \N__35572\,
            I => \foc.u_Park_Transform.n16983\
        );

    \I__4749\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35566\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__35566\,
            I => \foc.u_Park_Transform.n366_adj_2013\
        );

    \I__4747\ : InMux
    port map (
            O => \N__35563\,
            I => \foc.u_Park_Transform.n16999\
        );

    \I__4746\ : InMux
    port map (
            O => \N__35560\,
            I => \bfn_13_14_0_\
        );

    \I__4745\ : InMux
    port map (
            O => \N__35557\,
            I => \foc.u_Park_Transform.n17001\
        );

    \I__4744\ : InMux
    port map (
            O => \N__35554\,
            I => \foc.u_Park_Transform.n17002\
        );

    \I__4743\ : InMux
    port map (
            O => \N__35551\,
            I => \foc.u_Park_Transform.n17003\
        );

    \I__4742\ : InMux
    port map (
            O => \N__35548\,
            I => \foc.u_Park_Transform.n17004\
        );

    \I__4741\ : InMux
    port map (
            O => \N__35545\,
            I => \foc.u_Park_Transform.n17005\
        );

    \I__4740\ : InMux
    port map (
            O => \N__35542\,
            I => \N__35538\
        );

    \I__4739\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35535\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__35538\,
            I => \foc.u_Park_Transform.n757\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__35535\,
            I => \foc.u_Park_Transform.n757\
        );

    \I__4736\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35527\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__35527\,
            I => \N__35524\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__35524\,
            I => \foc.u_Park_Transform.n758\
        );

    \I__4733\ : InMux
    port map (
            O => \N__35521\,
            I => \foc.u_Park_Transform.n17006\
        );

    \I__4732\ : InMux
    port map (
            O => \N__35518\,
            I => \foc.u_Park_Transform.n759\
        );

    \I__4731\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35512\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35509\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__35509\,
            I => \N__35506\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__35506\,
            I => \foc.u_Park_Transform.n759_THRU_CO\
        );

    \I__4727\ : CascadeMux
    port map (
            O => \N__35503\,
            I => \N__35500\
        );

    \I__4726\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35497\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__35497\,
            I => \foc.u_Park_Transform.n703_adj_2160\
        );

    \I__4724\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35491\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__35491\,
            I => \N__35488\
        );

    \I__4722\ : Odrv12
    port map (
            O => \N__35488\,
            I => \foc.u_Park_Transform.n754_adj_2159\
        );

    \I__4721\ : InMux
    port map (
            O => \N__35485\,
            I => \foc.u_Park_Transform.n17204\
        );

    \I__4720\ : InMux
    port map (
            O => \N__35482\,
            I => \foc.u_Park_Transform.n755_adj_2161\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__35479\,
            I => \N__35476\
        );

    \I__4718\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35473\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__35473\,
            I => \N__35470\
        );

    \I__4716\ : Odrv12
    port map (
            O => \N__35470\,
            I => \foc.u_Park_Transform.n755_adj_2161_THRU_CO\
        );

    \I__4715\ : InMux
    port map (
            O => \N__35467\,
            I => \foc.u_Park_Transform.n16993\
        );

    \I__4714\ : InMux
    port map (
            O => \N__35464\,
            I => \foc.u_Park_Transform.n16994\
        );

    \I__4713\ : InMux
    port map (
            O => \N__35461\,
            I => \foc.u_Park_Transform.n16995\
        );

    \I__4712\ : InMux
    port map (
            O => \N__35458\,
            I => \foc.u_Park_Transform.n16996\
        );

    \I__4711\ : InMux
    port map (
            O => \N__35455\,
            I => \foc.u_Park_Transform.n16997\
        );

    \I__4710\ : InMux
    port map (
            O => \N__35452\,
            I => \foc.u_Park_Transform.n16998\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__35449\,
            I => \N__35446\
        );

    \I__4708\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35443\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__35443\,
            I => \foc.u_Park_Transform.n262_adj_1996\
        );

    \I__4706\ : InMux
    port map (
            O => \N__35440\,
            I => \foc.u_Park_Transform.n17195\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__35437\,
            I => \N__35434\
        );

    \I__4704\ : InMux
    port map (
            O => \N__35434\,
            I => \N__35431\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__35431\,
            I => \foc.u_Park_Transform.n311\
        );

    \I__4702\ : InMux
    port map (
            O => \N__35428\,
            I => \foc.u_Park_Transform.n17196\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \N__35422\
        );

    \I__4700\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35419\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__35419\,
            I => \foc.u_Park_Transform.n360\
        );

    \I__4698\ : InMux
    port map (
            O => \N__35416\,
            I => \foc.u_Park_Transform.n17197\
        );

    \I__4697\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35410\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__35410\,
            I => \foc.u_Park_Transform.n409\
        );

    \I__4695\ : InMux
    port map (
            O => \N__35407\,
            I => \bfn_13_12_0_\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__35404\,
            I => \N__35401\
        );

    \I__4693\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35398\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__35398\,
            I => \foc.u_Park_Transform.n458\
        );

    \I__4691\ : InMux
    port map (
            O => \N__35395\,
            I => \foc.u_Park_Transform.n17199\
        );

    \I__4690\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35389\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__35389\,
            I => \foc.u_Park_Transform.n507_adj_2165\
        );

    \I__4688\ : InMux
    port map (
            O => \N__35386\,
            I => \foc.u_Park_Transform.n17200\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__35383\,
            I => \N__35380\
        );

    \I__4686\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35377\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__35377\,
            I => \foc.u_Park_Transform.n556_adj_2164\
        );

    \I__4684\ : InMux
    port map (
            O => \N__35374\,
            I => \foc.u_Park_Transform.n17201\
        );

    \I__4683\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35368\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__35368\,
            I => \foc.u_Park_Transform.n605_adj_2163\
        );

    \I__4681\ : InMux
    port map (
            O => \N__35365\,
            I => \foc.u_Park_Transform.n17202\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__35362\,
            I => \N__35359\
        );

    \I__4679\ : InMux
    port map (
            O => \N__35359\,
            I => \N__35356\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__35356\,
            I => \foc.u_Park_Transform.n654_adj_2162\
        );

    \I__4677\ : InMux
    port map (
            O => \N__35353\,
            I => \foc.u_Park_Transform.n17203\
        );

    \I__4676\ : InMux
    port map (
            O => \N__35350\,
            I => \N__35347\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__35347\,
            I => \N__35344\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__35344\,
            I => \N__35341\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__35341\,
            I => \foc.u_Park_Transform.n786_adj_2152\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__35338\,
            I => \N__35335\
        );

    \I__4671\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35332\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__35332\,
            I => \N__35329\
        );

    \I__4669\ : Odrv4
    port map (
            O => \N__35329\,
            I => \foc.u_Park_Transform.n783_THRU_CO\
        );

    \I__4668\ : InMux
    port map (
            O => \N__35326\,
            I => \foc.u_Park_Transform.n17095\
        );

    \I__4667\ : InMux
    port map (
            O => \N__35323\,
            I => \N__35320\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__35320\,
            I => \N__35317\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__35317\,
            I => \N__35313\
        );

    \I__4664\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35310\
        );

    \I__4663\ : Sp12to4
    port map (
            O => \N__35313\,
            I => \N__35305\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__35310\,
            I => \N__35305\
        );

    \I__4661\ : Odrv12
    port map (
            O => \N__35305\,
            I => \foc.u_Park_Transform.n790\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__35302\,
            I => \N__35299\
        );

    \I__4659\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35296\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__35296\,
            I => \N__35293\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__35293\,
            I => \N__35290\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__35290\,
            I => \foc.u_Park_Transform.n787_adj_2149_THRU_CO\
        );

    \I__4655\ : InMux
    port map (
            O => \N__35287\,
            I => \foc.u_Park_Transform.n17096\
        );

    \I__4654\ : InMux
    port map (
            O => \N__35284\,
            I => \foc.u_Park_Transform.n17097\
        );

    \I__4653\ : InMux
    port map (
            O => \N__35281\,
            I => \N__35278\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__35278\,
            I => \foc.u_Park_Transform.n66\
        );

    \I__4651\ : InMux
    port map (
            O => \N__35275\,
            I => \foc.u_Park_Transform.n17191\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__35272\,
            I => \N__35269\
        );

    \I__4649\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35266\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__35266\,
            I => \foc.u_Park_Transform.n115\
        );

    \I__4647\ : InMux
    port map (
            O => \N__35263\,
            I => \foc.u_Park_Transform.n17192\
        );

    \I__4646\ : CascadeMux
    port map (
            O => \N__35260\,
            I => \N__35257\
        );

    \I__4645\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35254\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__35254\,
            I => \foc.u_Park_Transform.n164\
        );

    \I__4643\ : InMux
    port map (
            O => \N__35251\,
            I => \foc.u_Park_Transform.n17193\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__35248\,
            I => \N__35245\
        );

    \I__4641\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35242\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__35242\,
            I => \foc.u_Park_Transform.n213\
        );

    \I__4639\ : InMux
    port map (
            O => \N__35239\,
            I => \foc.u_Park_Transform.n17194\
        );

    \I__4638\ : InMux
    port map (
            O => \N__35236\,
            I => \foc.u_Park_Transform.n17087\
        );

    \I__4637\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35230\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__35230\,
            I => \N__35227\
        );

    \I__4635\ : Span4Mux_v
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__35224\,
            I => \foc.u_Park_Transform.n758_adj_2168\
        );

    \I__4633\ : InMux
    port map (
            O => \N__35221\,
            I => \foc.u_Park_Transform.n17088\
        );

    \I__4632\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35215\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__35215\,
            I => \N__35212\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__35212\,
            I => \N__35209\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__35209\,
            I => \foc.u_Park_Transform.n759_adj_2166_THRU_CO\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__35206\,
            I => \N__35203\
        );

    \I__4627\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35200\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__35200\,
            I => \foc.u_Park_Transform.n762\
        );

    \I__4625\ : InMux
    port map (
            O => \N__35197\,
            I => \foc.u_Park_Transform.n17089\
        );

    \I__4624\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35191\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__35191\,
            I => \N__35188\
        );

    \I__4622\ : Odrv12
    port map (
            O => \N__35188\,
            I => \foc.u_Park_Transform.n766\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__35185\,
            I => \N__35182\
        );

    \I__4620\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35179\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__35179\,
            I => \foc.u_Park_Transform.n763_THRU_CO\
        );

    \I__4618\ : InMux
    port map (
            O => \N__35176\,
            I => \bfn_13_10_0_\
        );

    \I__4617\ : InMux
    port map (
            O => \N__35173\,
            I => \N__35170\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__35167\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__35167\,
            I => \N__35164\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__35164\,
            I => \foc.u_Park_Transform.n770_adj_2030\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__35161\,
            I => \N__35158\
        );

    \I__4612\ : InMux
    port map (
            O => \N__35158\,
            I => \N__35155\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__35155\,
            I => \N__35152\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__35152\,
            I => \foc.u_Park_Transform.n767_THRU_CO\
        );

    \I__4609\ : InMux
    port map (
            O => \N__35149\,
            I => \foc.u_Park_Transform.n17091\
        );

    \I__4608\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35143\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__35143\,
            I => \N__35140\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__35140\,
            I => \N__35137\
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__35137\,
            I => \foc.u_Park_Transform.n774_adj_2045\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__35134\,
            I => \N__35131\
        );

    \I__4603\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35128\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__35128\,
            I => \N__35125\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__35125\,
            I => \N__35122\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__35122\,
            I => \foc.u_Park_Transform.n771_adj_2032_THRU_CO\
        );

    \I__4599\ : InMux
    port map (
            O => \N__35119\,
            I => \foc.u_Park_Transform.n17092\
        );

    \I__4598\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35113\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__35113\,
            I => \N__35110\
        );

    \I__4596\ : Odrv12
    port map (
            O => \N__35110\,
            I => \foc.u_Park_Transform.n778_adj_2068\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__35107\,
            I => \N__35104\
        );

    \I__4594\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35101\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__35101\,
            I => \N__35098\
        );

    \I__4592\ : Span4Mux_v
    port map (
            O => \N__35098\,
            I => \N__35095\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__35095\,
            I => \foc.u_Park_Transform.n775_adj_2047_THRU_CO\
        );

    \I__4590\ : InMux
    port map (
            O => \N__35092\,
            I => \foc.u_Park_Transform.n17093\
        );

    \I__4589\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35086\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__35086\,
            I => \N__35083\
        );

    \I__4587\ : Odrv4
    port map (
            O => \N__35083\,
            I => \foc.u_Park_Transform.n782_adj_2109\
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__35080\,
            I => \N__35077\
        );

    \I__4585\ : InMux
    port map (
            O => \N__35077\,
            I => \N__35074\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__35074\,
            I => \N__35071\
        );

    \I__4583\ : Odrv12
    port map (
            O => \N__35071\,
            I => \foc.u_Park_Transform.n779_adj_2070_THRU_CO\
        );

    \I__4582\ : InMux
    port map (
            O => \N__35068\,
            I => \foc.u_Park_Transform.n17094\
        );

    \I__4581\ : InMux
    port map (
            O => \N__35065\,
            I => \foc.u_Park_Transform.n17083\
        );

    \I__4580\ : InMux
    port map (
            O => \N__35062\,
            I => \foc.u_Park_Transform.n17084\
        );

    \I__4579\ : InMux
    port map (
            O => \N__35059\,
            I => \foc.u_Park_Transform.n17085\
        );

    \I__4578\ : InMux
    port map (
            O => \N__35056\,
            I => \foc.u_Park_Transform.n17086\
        );

    \I__4577\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35050\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35047\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__35047\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n470\
        );

    \I__4574\ : InMux
    port map (
            O => \N__35044\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18115\
        );

    \I__4573\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35038\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__35035\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__35035\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n519\
        );

    \I__4570\ : InMux
    port map (
            O => \N__35032\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18116\
        );

    \I__4569\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35026\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__35026\,
            I => \N__35023\
        );

    \I__4567\ : Odrv12
    port map (
            O => \N__35023\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n568\
        );

    \I__4566\ : InMux
    port map (
            O => \N__35020\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18117\
        );

    \I__4565\ : InMux
    port map (
            O => \N__35017\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18118\
        );

    \I__4564\ : InMux
    port map (
            O => \N__35014\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18119\
        );

    \I__4563\ : CascadeMux
    port map (
            O => \N__35011\,
            I => \N__35007\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__35010\,
            I => \N__35004\
        );

    \I__4561\ : InMux
    port map (
            O => \N__35007\,
            I => \N__35000\
        );

    \I__4560\ : InMux
    port map (
            O => \N__35004\,
            I => \N__34995\
        );

    \I__4559\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34995\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__35000\,
            I => \N__34990\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__34995\,
            I => \N__34990\
        );

    \I__4556\ : Odrv4
    port map (
            O => \N__34990\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n617\
        );

    \I__4555\ : InMux
    port map (
            O => \N__34987\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18120\
        );

    \I__4554\ : InMux
    port map (
            O => \N__34984\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598\
        );

    \I__4553\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34978\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34975\
        );

    \I__4551\ : Odrv12
    port map (
            O => \N__34975\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n78_adj_617\
        );

    \I__4550\ : InMux
    port map (
            O => \N__34972\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18107\
        );

    \I__4549\ : InMux
    port map (
            O => \N__34969\,
            I => \N__34966\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34963\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__34963\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n127_adj_615\
        );

    \I__4546\ : InMux
    port map (
            O => \N__34960\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18108\
        );

    \I__4545\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34954\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__34954\,
            I => \N__34951\
        );

    \I__4543\ : Odrv12
    port map (
            O => \N__34951\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n176_adj_613\
        );

    \I__4542\ : InMux
    port map (
            O => \N__34948\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18109\
        );

    \I__4541\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34942\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__34942\,
            I => \N__34939\
        );

    \I__4539\ : Odrv12
    port map (
            O => \N__34939\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n225_adj_611\
        );

    \I__4538\ : InMux
    port map (
            O => \N__34936\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18110\
        );

    \I__4537\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34930\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34927\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__34927\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n274_adj_609\
        );

    \I__4534\ : InMux
    port map (
            O => \N__34924\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18111\
        );

    \I__4533\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34918\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__34918\,
            I => \N__34915\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__34915\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n323_adj_607\
        );

    \I__4530\ : InMux
    port map (
            O => \N__34912\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18112\
        );

    \I__4529\ : InMux
    port map (
            O => \N__34909\,
            I => \N__34906\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__34906\,
            I => \N__34903\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__34903\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n372\
        );

    \I__4526\ : InMux
    port map (
            O => \N__34900\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18113\
        );

    \I__4525\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34894\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__34894\,
            I => \N__34891\
        );

    \I__4523\ : Odrv12
    port map (
            O => \N__34891\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n421\
        );

    \I__4522\ : InMux
    port map (
            O => \N__34888\,
            I => \bfn_12_25_0_\
        );

    \I__4521\ : InMux
    port map (
            O => \N__34885\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17661\
        );

    \I__4520\ : InMux
    port map (
            O => \N__34882\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17662\
        );

    \I__4519\ : InMux
    port map (
            O => \N__34879\,
            I => \bfn_12_23_0_\
        );

    \I__4518\ : InMux
    port map (
            O => \N__34876\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17664\
        );

    \I__4517\ : InMux
    port map (
            O => \N__34873\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17665\
        );

    \I__4516\ : InMux
    port map (
            O => \N__34870\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17666\
        );

    \I__4515\ : InMux
    port map (
            O => \N__34867\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17667\
        );

    \I__4514\ : InMux
    port map (
            O => \N__34864\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775\
        );

    \I__4513\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34858\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__34858\,
            I => \N__34855\
        );

    \I__4511\ : Odrv12
    port map (
            O => \N__34855\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3017\
        );

    \I__4510\ : InMux
    port map (
            O => \N__34852\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382\
        );

    \I__4509\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34846\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__34846\,
            I => \N__34843\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__34843\,
            I => \N__34840\
        );

    \I__4506\ : Odrv4
    port map (
            O => \N__34840\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3117\
        );

    \I__4505\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34834\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__34834\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3219\
        );

    \I__4503\ : InMux
    port map (
            O => \N__34831\,
            I => \bfn_12_20_0_\
        );

    \I__4502\ : InMux
    port map (
            O => \N__34828\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__34825\,
            I => \N__34822\
        );

    \I__4500\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34819\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__34819\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_CO\
        );

    \I__4498\ : InMux
    port map (
            O => \N__34816\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17656\
        );

    \I__4497\ : InMux
    port map (
            O => \N__34813\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17657\
        );

    \I__4496\ : InMux
    port map (
            O => \N__34810\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17658\
        );

    \I__4495\ : InMux
    port map (
            O => \N__34807\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17659\
        );

    \I__4494\ : InMux
    port map (
            O => \N__34804\,
            I => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17660\
        );

    \I__4493\ : InMux
    port map (
            O => \N__34801\,
            I => \foc.u_Park_Transform.n16914\
        );

    \I__4492\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34792\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__34797\,
            I => \N__34788\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__34796\,
            I => \N__34784\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__34795\,
            I => \N__34780\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__34792\,
            I => \N__34776\
        );

    \I__4487\ : InMux
    port map (
            O => \N__34791\,
            I => \N__34761\
        );

    \I__4486\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34761\
        );

    \I__4485\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34761\
        );

    \I__4484\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34761\
        );

    \I__4483\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34761\
        );

    \I__4482\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34761\
        );

    \I__4481\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34761\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__34776\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__34761\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__34756\,
            I => \N__34753\
        );

    \I__4477\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34750\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__34750\,
            I => \N__34747\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__34747\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2417\
        );

    \I__4474\ : InMux
    port map (
            O => \N__34744\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376\
        );

    \I__4473\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34738\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__34738\,
            I => \N__34735\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__34735\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2517\
        );

    \I__4470\ : InMux
    port map (
            O => \N__34732\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__34729\,
            I => \N__34726\
        );

    \I__4468\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34723\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__34723\,
            I => \N__34720\
        );

    \I__4466\ : Odrv12
    port map (
            O => \N__34720\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2617\
        );

    \I__4465\ : InMux
    port map (
            O => \N__34717\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378\
        );

    \I__4464\ : InMux
    port map (
            O => \N__34714\,
            I => \N__34711\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__34711\,
            I => \N__34708\
        );

    \I__4462\ : Odrv12
    port map (
            O => \N__34708\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2717\
        );

    \I__4461\ : InMux
    port map (
            O => \N__34705\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379\
        );

    \I__4460\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34699\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__34699\,
            I => \N__34696\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__34696\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2817\
        );

    \I__4457\ : InMux
    port map (
            O => \N__34693\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380\
        );

    \I__4456\ : InMux
    port map (
            O => \N__34690\,
            I => \N__34687\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__34687\,
            I => \N__34684\
        );

    \I__4454\ : Odrv12
    port map (
            O => \N__34684\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2917\
        );

    \I__4453\ : InMux
    port map (
            O => \N__34681\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381\
        );

    \I__4452\ : InMux
    port map (
            O => \N__34678\,
            I => \foc.u_Park_Transform.n16905\
        );

    \I__4451\ : InMux
    port map (
            O => \N__34675\,
            I => \foc.u_Park_Transform.n16906\
        );

    \I__4450\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34669\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34666\
        );

    \I__4448\ : Odrv12
    port map (
            O => \N__34666\,
            I => \foc.u_Park_Transform.n766_adj_2053\
        );

    \I__4447\ : InMux
    port map (
            O => \N__34663\,
            I => \bfn_12_18_0_\
        );

    \I__4446\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34657\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__34657\,
            I => \N__34654\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__34654\,
            I => \foc.u_Park_Transform.n770\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__34651\,
            I => \N__34648\
        );

    \I__4442\ : InMux
    port map (
            O => \N__34648\,
            I => \N__34645\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__34645\,
            I => \N__34642\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__34642\,
            I => \foc.u_Park_Transform.n767_adj_2041_THRU_CO\
        );

    \I__4439\ : InMux
    port map (
            O => \N__34639\,
            I => \foc.u_Park_Transform.n16908\
        );

    \I__4438\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34633\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__4436\ : Span4Mux_h
    port map (
            O => \N__34630\,
            I => \N__34627\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__34627\,
            I => \foc.u_Park_Transform.n774\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__4433\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34618\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34615\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__34615\,
            I => \foc.u_Park_Transform.n771_THRU_CO\
        );

    \I__4430\ : InMux
    port map (
            O => \N__34612\,
            I => \foc.u_Park_Transform.n16909\
        );

    \I__4429\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34606\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34603\
        );

    \I__4427\ : Odrv12
    port map (
            O => \N__34603\,
            I => \foc.u_Park_Transform.n778\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__34600\,
            I => \N__34597\
        );

    \I__4425\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34594\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__34594\,
            I => \N__34591\
        );

    \I__4423\ : Span12Mux_v
    port map (
            O => \N__34591\,
            I => \N__34588\
        );

    \I__4422\ : Odrv12
    port map (
            O => \N__34588\,
            I => \foc.u_Park_Transform.n775_THRU_CO\
        );

    \I__4421\ : InMux
    port map (
            O => \N__34585\,
            I => \foc.u_Park_Transform.n16910\
        );

    \I__4420\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34579\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__34579\,
            I => \N__34576\
        );

    \I__4418\ : Span4Mux_h
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__34573\,
            I => \foc.u_Park_Transform.n782\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__4415\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34564\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34561\
        );

    \I__4413\ : Odrv12
    port map (
            O => \N__34561\,
            I => \foc.u_Park_Transform.n779_THRU_CO\
        );

    \I__4412\ : InMux
    port map (
            O => \N__34558\,
            I => \foc.u_Park_Transform.n16911\
        );

    \I__4411\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34552\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__34552\,
            I => \N__34549\
        );

    \I__4409\ : Span12Mux_v
    port map (
            O => \N__34549\,
            I => \N__34546\
        );

    \I__4408\ : Odrv12
    port map (
            O => \N__34546\,
            I => \foc.u_Park_Transform.n786\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__34543\,
            I => \N__34540\
        );

    \I__4406\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34537\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__34537\,
            I => \N__34534\
        );

    \I__4404\ : Span4Mux_v
    port map (
            O => \N__34534\,
            I => \N__34531\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__34531\,
            I => \foc.u_Park_Transform.n783_adj_2167_THRU_CO\
        );

    \I__4402\ : InMux
    port map (
            O => \N__34528\,
            I => \foc.u_Park_Transform.n16912\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__34525\,
            I => \N__34522\
        );

    \I__4400\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34519\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__34519\,
            I => \N__34516\
        );

    \I__4398\ : Span4Mux_v
    port map (
            O => \N__34516\,
            I => \N__34513\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__34513\,
            I => \foc.u_Park_Transform.n787_THRU_CO\
        );

    \I__4396\ : InMux
    port map (
            O => \N__34510\,
            I => \foc.u_Park_Transform.n16913\
        );

    \I__4395\ : InMux
    port map (
            O => \N__34507\,
            I => \foc.u_Park_Transform.n16975\
        );

    \I__4394\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34501\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__34501\,
            I => \N__34497\
        );

    \I__4392\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34494\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__34497\,
            I => \N__34491\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__34494\,
            I => \N__34488\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__34491\,
            I => \foc.u_Park_Transform.n765\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__34488\,
            I => \foc.u_Park_Transform.n765\
        );

    \I__4387\ : CascadeMux
    port map (
            O => \N__34483\,
            I => \N__34480\
        );

    \I__4386\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34477\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__34477\,
            I => \foc.u_Park_Transform.n712\
        );

    \I__4384\ : InMux
    port map (
            O => \N__34474\,
            I => \foc.u_Park_Transform.n16976\
        );

    \I__4383\ : InMux
    port map (
            O => \N__34471\,
            I => \foc.u_Park_Transform.n767_adj_2041\
        );

    \I__4382\ : InMux
    port map (
            O => \N__34468\,
            I => \foc.u_Park_Transform.n16900\
        );

    \I__4381\ : InMux
    port map (
            O => \N__34465\,
            I => \foc.u_Park_Transform.n16901\
        );

    \I__4380\ : InMux
    port map (
            O => \N__34462\,
            I => \foc.u_Park_Transform.n16902\
        );

    \I__4379\ : InMux
    port map (
            O => \N__34459\,
            I => \foc.u_Park_Transform.n16903\
        );

    \I__4378\ : InMux
    port map (
            O => \N__34456\,
            I => \foc.u_Park_Transform.n16904\
        );

    \I__4377\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34450\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__34450\,
            I => \foc.u_Park_Transform.n271_adj_2043\
        );

    \I__4375\ : InMux
    port map (
            O => \N__34447\,
            I => \foc.u_Park_Transform.n16967\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__4373\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34438\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__34438\,
            I => \foc.u_Park_Transform.n320_adj_2036\
        );

    \I__4371\ : InMux
    port map (
            O => \N__34435\,
            I => \foc.u_Park_Transform.n16968\
        );

    \I__4370\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34429\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__34429\,
            I => \foc.u_Park_Transform.n369_adj_2026\
        );

    \I__4368\ : InMux
    port map (
            O => \N__34426\,
            I => \foc.u_Park_Transform.n16969\
        );

    \I__4367\ : CascadeMux
    port map (
            O => \N__34423\,
            I => \N__34420\
        );

    \I__4366\ : InMux
    port map (
            O => \N__34420\,
            I => \N__34417\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__34417\,
            I => \foc.u_Park_Transform.n418\
        );

    \I__4364\ : InMux
    port map (
            O => \N__34414\,
            I => \bfn_12_16_0_\
        );

    \I__4363\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34408\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__34408\,
            I => \foc.u_Park_Transform.n467\
        );

    \I__4361\ : InMux
    port map (
            O => \N__34405\,
            I => \foc.u_Park_Transform.n16971\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__34402\,
            I => \N__34399\
        );

    \I__4359\ : InMux
    port map (
            O => \N__34399\,
            I => \N__34396\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__34396\,
            I => \foc.u_Park_Transform.n516\
        );

    \I__4357\ : InMux
    port map (
            O => \N__34393\,
            I => \foc.u_Park_Transform.n16972\
        );

    \I__4356\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34387\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__34387\,
            I => \foc.u_Park_Transform.n565_adj_2020\
        );

    \I__4354\ : InMux
    port map (
            O => \N__34384\,
            I => \foc.u_Park_Transform.n16973\
        );

    \I__4353\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34378\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__34378\,
            I => \foc.u_Park_Transform.n614\
        );

    \I__4351\ : InMux
    port map (
            O => \N__34375\,
            I => \foc.u_Park_Transform.n16974\
        );

    \I__4350\ : InMux
    port map (
            O => \N__34372\,
            I => \N__34369\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__34369\,
            I => \foc.u_Park_Transform.n663\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__34366\,
            I => \n4_cascade_\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__34363\,
            I => \N__34357\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__34362\,
            I => \N__34353\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__34361\,
            I => \N__34350\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__34360\,
            I => \N__34346\
        );

    \I__4343\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34339\
        );

    \I__4342\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34339\
        );

    \I__4341\ : InMux
    port map (
            O => \N__34353\,
            I => \N__34339\
        );

    \I__4340\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34332\
        );

    \I__4339\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34332\
        );

    \I__4338\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34332\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__34339\,
            I => \N__34329\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__34332\,
            I => \N__34326\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__34329\,
            I => \foc.u_Park_Transform.n237\
        );

    \I__4334\ : Odrv12
    port map (
            O => \N__34326\,
            I => \foc.u_Park_Transform.n237\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__34321\,
            I => \N__34318\
        );

    \I__4332\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34314\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__34317\,
            I => \N__34311\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__34314\,
            I => \N__34308\
        );

    \I__4329\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34305\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__34308\,
            I => \N__34302\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__34305\,
            I => \N__34299\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__34302\,
            I => \foc.u_Park_Transform.n188\
        );

    \I__4325\ : Odrv12
    port map (
            O => \N__34299\,
            I => \foc.u_Park_Transform.n188\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__34294\,
            I => \N__34288\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__34293\,
            I => \N__34285\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__34292\,
            I => \N__34281\
        );

    \I__4321\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34267\
        );

    \I__4320\ : InMux
    port map (
            O => \N__34288\,
            I => \N__34267\
        );

    \I__4319\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34258\
        );

    \I__4318\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34258\
        );

    \I__4317\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34258\
        );

    \I__4316\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34258\
        );

    \I__4315\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34255\
        );

    \I__4314\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34252\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__34277\,
            I => \N__34246\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__34276\,
            I => \N__34240\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__34275\,
            I => \N__34237\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__34274\,
            I => \N__34233\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__34273\,
            I => \N__34229\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__34272\,
            I => \N__34224\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__34267\,
            I => \N__34216\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__34258\,
            I => \N__34216\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34213\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__34252\,
            I => \N__34210\
        );

    \I__4303\ : InMux
    port map (
            O => \N__34251\,
            I => \N__34201\
        );

    \I__4302\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34201\
        );

    \I__4301\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34201\
        );

    \I__4300\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34201\
        );

    \I__4299\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34192\
        );

    \I__4298\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34192\
        );

    \I__4297\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34192\
        );

    \I__4296\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34192\
        );

    \I__4295\ : InMux
    port map (
            O => \N__34237\,
            I => \N__34179\
        );

    \I__4294\ : InMux
    port map (
            O => \N__34236\,
            I => \N__34179\
        );

    \I__4293\ : InMux
    port map (
            O => \N__34233\,
            I => \N__34179\
        );

    \I__4292\ : InMux
    port map (
            O => \N__34232\,
            I => \N__34179\
        );

    \I__4291\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34179\
        );

    \I__4290\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34179\
        );

    \I__4289\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34174\
        );

    \I__4288\ : InMux
    port map (
            O => \N__34224\,
            I => \N__34174\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__34223\,
            I => \N__34170\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__34222\,
            I => \N__34166\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__34221\,
            I => \N__34162\
        );

    \I__4284\ : Span4Mux_v
    port map (
            O => \N__34216\,
            I => \N__34151\
        );

    \I__4283\ : Span4Mux_h
    port map (
            O => \N__34213\,
            I => \N__34151\
        );

    \I__4282\ : Span4Mux_v
    port map (
            O => \N__34210\,
            I => \N__34151\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__34201\,
            I => \N__34151\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__34192\,
            I => \N__34151\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__34179\,
            I => \N__34146\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__34146\
        );

    \I__4277\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34133\
        );

    \I__4276\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34133\
        );

    \I__4275\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34133\
        );

    \I__4274\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34133\
        );

    \I__4273\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34133\
        );

    \I__4272\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34133\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__34151\,
            I => \foc.u_Park_Transform.n613\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__34146\,
            I => \foc.u_Park_Transform.n613\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__34133\,
            I => \foc.u_Park_Transform.n613\
        );

    \I__4268\ : InMux
    port map (
            O => \N__34126\,
            I => \N__34123\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__34123\,
            I => \foc.u_Park_Transform.n75_adj_2123\
        );

    \I__4266\ : InMux
    port map (
            O => \N__34120\,
            I => \foc.u_Park_Transform.n16963\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__34117\,
            I => \N__34114\
        );

    \I__4264\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__34111\,
            I => \foc.u_Park_Transform.n124_adj_2090\
        );

    \I__4262\ : InMux
    port map (
            O => \N__34108\,
            I => \foc.u_Park_Transform.n16964\
        );

    \I__4261\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34102\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__34102\,
            I => \foc.u_Park_Transform.n173_adj_2061\
        );

    \I__4259\ : InMux
    port map (
            O => \N__34099\,
            I => \foc.u_Park_Transform.n16965\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__34096\,
            I => \N__34093\
        );

    \I__4257\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34090\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__34090\,
            I => \foc.u_Park_Transform.n222_adj_2049\
        );

    \I__4255\ : InMux
    port map (
            O => \N__34087\,
            I => \foc.u_Park_Transform.n16966\
        );

    \I__4254\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34078\
        );

    \I__4253\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34078\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__34078\,
            I => \foc.Look_Up_Table_out1_1_3\
        );

    \I__4251\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34069\
        );

    \I__4250\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34069\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__34069\,
            I => \foc.Look_Up_Table_out1_1_5\
        );

    \I__4248\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34060\
        );

    \I__4247\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34060\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__34060\,
            I => \foc.Look_Up_Table_out1_1_4\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__34057\,
            I => \N__34054\
        );

    \I__4244\ : InMux
    port map (
            O => \N__34054\,
            I => \N__34051\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__34051\,
            I => \N__34048\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__34048\,
            I => \foc.u_Park_Transform.n412\
        );

    \I__4241\ : InMux
    port map (
            O => \N__34045\,
            I => \bfn_12_12_0_\
        );

    \I__4240\ : InMux
    port map (
            O => \N__34042\,
            I => \N__34039\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__34039\,
            I => \N__34036\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__34036\,
            I => \foc.u_Park_Transform.n461\
        );

    \I__4237\ : InMux
    port map (
            O => \N__34033\,
            I => \foc.u_Park_Transform.n17184\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__34030\,
            I => \N__34027\
        );

    \I__4235\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34024\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__34024\,
            I => \N__34021\
        );

    \I__4233\ : Odrv12
    port map (
            O => \N__34021\,
            I => \foc.u_Park_Transform.n510_adj_2004\
        );

    \I__4232\ : InMux
    port map (
            O => \N__34018\,
            I => \foc.u_Park_Transform.n17185\
        );

    \I__4231\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34012\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__34012\,
            I => \N__34009\
        );

    \I__4229\ : Odrv12
    port map (
            O => \N__34009\,
            I => \foc.u_Park_Transform.n559_adj_2001\
        );

    \I__4228\ : InMux
    port map (
            O => \N__34006\,
            I => \foc.u_Park_Transform.n17186\
        );

    \I__4227\ : InMux
    port map (
            O => \N__34003\,
            I => \N__34000\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__34000\,
            I => \N__33997\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__33997\,
            I => \foc.u_Park_Transform.n608\
        );

    \I__4224\ : InMux
    port map (
            O => \N__33994\,
            I => \foc.u_Park_Transform.n17187\
        );

    \I__4223\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33988\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33985\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__33985\,
            I => \foc.u_Park_Transform.n657\
        );

    \I__4220\ : InMux
    port map (
            O => \N__33982\,
            I => \foc.u_Park_Transform.n17188\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__33979\,
            I => \N__33976\
        );

    \I__4218\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33970\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__33970\,
            I => \foc.u_Park_Transform.n706\
        );

    \I__4215\ : InMux
    port map (
            O => \N__33967\,
            I => \foc.u_Park_Transform.n17189\
        );

    \I__4214\ : InMux
    port map (
            O => \N__33964\,
            I => \foc.u_Park_Transform.n759_adj_2166\
        );

    \I__4213\ : InMux
    port map (
            O => \N__33961\,
            I => \foc.u_Park_Transform.n763\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__33958\,
            I => \N__33955\
        );

    \I__4211\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33952\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__33952\,
            I => \N__33949\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__33949\,
            I => \foc.u_Park_Transform.n69\
        );

    \I__4208\ : InMux
    port map (
            O => \N__33946\,
            I => \foc.u_Park_Transform.n17176\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__33943\,
            I => \N__33940\
        );

    \I__4206\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33937\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__33937\,
            I => \N__33934\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__33934\,
            I => \foc.u_Park_Transform.n118\
        );

    \I__4203\ : InMux
    port map (
            O => \N__33931\,
            I => \foc.u_Park_Transform.n17177\
        );

    \I__4202\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33925\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33922\
        );

    \I__4200\ : Odrv12
    port map (
            O => \N__33922\,
            I => \foc.u_Park_Transform.n167\
        );

    \I__4199\ : InMux
    port map (
            O => \N__33919\,
            I => \foc.u_Park_Transform.n17178\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__33916\,
            I => \N__33913\
        );

    \I__4197\ : InMux
    port map (
            O => \N__33913\,
            I => \N__33910\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__33910\,
            I => \N__33907\
        );

    \I__4195\ : Odrv12
    port map (
            O => \N__33907\,
            I => \foc.u_Park_Transform.n216\
        );

    \I__4194\ : InMux
    port map (
            O => \N__33904\,
            I => \foc.u_Park_Transform.n17179\
        );

    \I__4193\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33898\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33895\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__33895\,
            I => \foc.u_Park_Transform.n265\
        );

    \I__4190\ : InMux
    port map (
            O => \N__33892\,
            I => \foc.u_Park_Transform.n17180\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__33889\,
            I => \N__33886\
        );

    \I__4188\ : InMux
    port map (
            O => \N__33886\,
            I => \N__33883\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__33883\,
            I => \N__33880\
        );

    \I__4186\ : Odrv4
    port map (
            O => \N__33880\,
            I => \foc.u_Park_Transform.n314\
        );

    \I__4185\ : InMux
    port map (
            O => \N__33877\,
            I => \foc.u_Park_Transform.n17181\
        );

    \I__4184\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33871\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33868\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__33868\,
            I => \foc.u_Park_Transform.n363\
        );

    \I__4181\ : InMux
    port map (
            O => \N__33865\,
            I => \foc.u_Park_Transform.n17182\
        );

    \I__4180\ : InMux
    port map (
            O => \N__33862\,
            I => \N__33859\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__33859\,
            I => \N__33856\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__33856\,
            I => \foc.u_Park_Transform.n366\
        );

    \I__4177\ : InMux
    port map (
            O => \N__33853\,
            I => \foc.u_Park_Transform.n17167\
        );

    \I__4176\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33847\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33844\
        );

    \I__4174\ : Span4Mux_v
    port map (
            O => \N__33844\,
            I => \N__33841\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__33841\,
            I => \foc.u_Park_Transform.n415_adj_2008\
        );

    \I__4172\ : InMux
    port map (
            O => \N__33838\,
            I => \bfn_12_10_0_\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__33835\,
            I => \N__33832\
        );

    \I__4170\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33829\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__33829\,
            I => \N__33826\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__33826\,
            I => \foc.u_Park_Transform.n464_adj_2005\
        );

    \I__4167\ : InMux
    port map (
            O => \N__33823\,
            I => \foc.u_Park_Transform.n17169\
        );

    \I__4166\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33817\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__33817\,
            I => \N__33814\
        );

    \I__4164\ : Odrv4
    port map (
            O => \N__33814\,
            I => \foc.u_Park_Transform.n513_adj_2002\
        );

    \I__4163\ : InMux
    port map (
            O => \N__33811\,
            I => \foc.u_Park_Transform.n17170\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__33808\,
            I => \N__33805\
        );

    \I__4161\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33802\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__33802\,
            I => \N__33799\
        );

    \I__4159\ : Odrv12
    port map (
            O => \N__33799\,
            I => \foc.u_Park_Transform.n562_adj_2000\
        );

    \I__4158\ : InMux
    port map (
            O => \N__33796\,
            I => \foc.u_Park_Transform.n17171\
        );

    \I__4157\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33790\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__4155\ : Odrv12
    port map (
            O => \N__33787\,
            I => \foc.u_Park_Transform.n611\
        );

    \I__4154\ : InMux
    port map (
            O => \N__33784\,
            I => \foc.u_Park_Transform.n17172\
        );

    \I__4153\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33778\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__33778\,
            I => \N__33775\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__33775\,
            I => \foc.u_Park_Transform.n660\
        );

    \I__4150\ : InMux
    port map (
            O => \N__33772\,
            I => \foc.u_Park_Transform.n17173\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__33769\,
            I => \N__33766\
        );

    \I__4148\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33763\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__33763\,
            I => \N__33760\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__33760\,
            I => \foc.u_Park_Transform.n709\
        );

    \I__4145\ : InMux
    port map (
            O => \N__33757\,
            I => \foc.u_Park_Transform.n17174\
        );

    \I__4144\ : InMux
    port map (
            O => \N__33754\,
            I => \bfn_11_24_0_\
        );

    \I__4143\ : InMux
    port map (
            O => \N__33751\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__33748\,
            I => \N__33745\
        );

    \I__4141\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33742\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__33742\,
            I => \N__33739\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__33739\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_CO\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__33736\,
            I => \N__33733\
        );

    \I__4137\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33730\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__33730\,
            I => \N__33727\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__33727\,
            I => \foc.u_Park_Transform.n72\
        );

    \I__4134\ : InMux
    port map (
            O => \N__33724\,
            I => \foc.u_Park_Transform.n17161\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__4132\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33715\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__33715\,
            I => \N__33712\
        );

    \I__4130\ : Odrv12
    port map (
            O => \N__33712\,
            I => \foc.u_Park_Transform.n121\
        );

    \I__4129\ : InMux
    port map (
            O => \N__33709\,
            I => \foc.u_Park_Transform.n17162\
        );

    \I__4128\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33703\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__33703\,
            I => \N__33700\
        );

    \I__4126\ : Odrv12
    port map (
            O => \N__33700\,
            I => \foc.u_Park_Transform.n170\
        );

    \I__4125\ : InMux
    port map (
            O => \N__33697\,
            I => \foc.u_Park_Transform.n17163\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__33694\,
            I => \N__33691\
        );

    \I__4123\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33688\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__33688\,
            I => \N__33685\
        );

    \I__4121\ : Odrv12
    port map (
            O => \N__33685\,
            I => \foc.u_Park_Transform.n219\
        );

    \I__4120\ : InMux
    port map (
            O => \N__33682\,
            I => \foc.u_Park_Transform.n17164\
        );

    \I__4119\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33676\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__33676\,
            I => \N__33673\
        );

    \I__4117\ : Odrv12
    port map (
            O => \N__33673\,
            I => \foc.u_Park_Transform.n268\
        );

    \I__4116\ : InMux
    port map (
            O => \N__33670\,
            I => \foc.u_Park_Transform.n17165\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__33667\,
            I => \N__33664\
        );

    \I__4114\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33661\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33658\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__33658\,
            I => \foc.u_Park_Transform.n317\
        );

    \I__4111\ : InMux
    port map (
            O => \N__33655\,
            I => \foc.u_Park_Transform.n17166\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__4109\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33646\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__33646\,
            I => \N__33643\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__33643\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2426\
        );

    \I__4106\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33637\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__33637\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2523\
        );

    \I__4104\ : InMux
    port map (
            O => \N__33634\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403\
        );

    \I__4103\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33628\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33625\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__33625\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2526\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__33622\,
            I => \N__33619\
        );

    \I__4099\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33616\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__33616\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2623\
        );

    \I__4097\ : InMux
    port map (
            O => \N__33613\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__4095\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33604\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__33604\,
            I => \N__33601\
        );

    \I__4093\ : Odrv12
    port map (
            O => \N__33601\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2626\
        );

    \I__4092\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33595\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__33595\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2723\
        );

    \I__4090\ : InMux
    port map (
            O => \N__33592\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405\
        );

    \I__4089\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33586\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33583\
        );

    \I__4087\ : Odrv4
    port map (
            O => \N__33583\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2726\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__4085\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__33574\,
            I => \N__33571\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__33571\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2823\
        );

    \I__4082\ : InMux
    port map (
            O => \N__33568\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406\
        );

    \I__4081\ : InMux
    port map (
            O => \N__33565\,
            I => \N__33562\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__33562\,
            I => \N__33559\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__33559\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2826\
        );

    \I__4078\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33553\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__33553\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2923\
        );

    \I__4076\ : InMux
    port map (
            O => \N__33550\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407\
        );

    \I__4075\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33544\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33541\
        );

    \I__4073\ : Odrv12
    port map (
            O => \N__33541\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2926\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__33538\,
            I => \N__33535\
        );

    \I__4071\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33532\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__33532\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3023\
        );

    \I__4069\ : InMux
    port map (
            O => \N__33529\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408\
        );

    \I__4068\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33523\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33520\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__33520\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3026\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__33517\,
            I => \N__33510\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__33516\,
            I => \N__33507\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__33515\,
            I => \N__33504\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__33514\,
            I => \N__33501\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__33513\,
            I => \N__33497\
        );

    \I__4060\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33490\
        );

    \I__4059\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33490\
        );

    \I__4058\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33479\
        );

    \I__4057\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33479\
        );

    \I__4056\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33479\
        );

    \I__4055\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33479\
        );

    \I__4054\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33479\
        );

    \I__4053\ : InMux
    port map (
            O => \N__33495\,
            I => \N__33476\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__33490\,
            I => \N__33471\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33471\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__33476\,
            I => \N__33468\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__33471\,
            I => \N__33465\
        );

    \I__4048\ : Span4Mux_v
    port map (
            O => \N__33468\,
            I => \N__33462\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__33465\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__33462\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822\
        );

    \I__4045\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33454\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__33454\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3123\
        );

    \I__4043\ : InMux
    port map (
            O => \N__33451\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409\
        );

    \I__4042\ : InMux
    port map (
            O => \N__33448\,
            I => \N__33445\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__33445\,
            I => \N__33442\
        );

    \I__4040\ : Odrv12
    port map (
            O => \N__33442\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3126\
        );

    \I__4039\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33436\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33433\
        );

    \I__4037\ : Odrv12
    port map (
            O => \N__33433\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3231\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__33430\,
            I => \N__33427\
        );

    \I__4035\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33424\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__33424\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2629\
        );

    \I__4033\ : InMux
    port map (
            O => \N__33421\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414\
        );

    \I__4032\ : InMux
    port map (
            O => \N__33418\,
            I => \N__33415\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__33415\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2729\
        );

    \I__4030\ : InMux
    port map (
            O => \N__33412\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415\
        );

    \I__4029\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33406\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__33406\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2829\
        );

    \I__4027\ : InMux
    port map (
            O => \N__33403\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416\
        );

    \I__4026\ : InMux
    port map (
            O => \N__33400\,
            I => \N__33397\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__33397\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2929\
        );

    \I__4024\ : InMux
    port map (
            O => \N__33394\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417\
        );

    \I__4023\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33388\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__33388\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3029\
        );

    \I__4021\ : InMux
    port map (
            O => \N__33385\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418\
        );

    \I__4020\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33379\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__33379\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3129\
        );

    \I__4018\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33373\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33370\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__33370\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3235\
        );

    \I__4015\ : InMux
    port map (
            O => \N__33367\,
            I => \bfn_11_22_0_\
        );

    \I__4014\ : InMux
    port map (
            O => \N__33364\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__33361\,
            I => \N__33358\
        );

    \I__4012\ : InMux
    port map (
            O => \N__33358\,
            I => \N__33355\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__33355\,
            I => \N__33352\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__33352\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_CO\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__33349\,
            I => \N__33341\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__33348\,
            I => \N__33338\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__33347\,
            I => \N__33335\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__33346\,
            I => \N__33332\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__33345\,
            I => \N__33328\
        );

    \I__4004\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33324\
        );

    \I__4003\ : InMux
    port map (
            O => \N__33341\,
            I => \N__33319\
        );

    \I__4002\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33319\
        );

    \I__4001\ : InMux
    port map (
            O => \N__33335\,
            I => \N__33308\
        );

    \I__4000\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33308\
        );

    \I__3999\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33308\
        );

    \I__3998\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33308\
        );

    \I__3997\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33308\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__33324\,
            I => \N__33301\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33301\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__33308\,
            I => \N__33301\
        );

    \I__3993\ : Span4Mux_v
    port map (
            O => \N__33301\,
            I => \N__33298\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__33298\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2825\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__33295\,
            I => \N__33292\
        );

    \I__3990\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33289\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__33289\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2423\
        );

    \I__3988\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33283\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__33283\,
            I => \N__33280\
        );

    \I__3986\ : Odrv12
    port map (
            O => \N__33280\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3247\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__33277\,
            I => \N__33274\
        );

    \I__3984\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33271\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__33271\,
            I => \N__33268\
        );

    \I__3982\ : Span4Mux_v
    port map (
            O => \N__33268\,
            I => \N__33265\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__33265\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_CO\
        );

    \I__3980\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33259\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__33259\,
            I => \N__33256\
        );

    \I__3978\ : Odrv12
    port map (
            O => \N__33256\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_43\
        );

    \I__3977\ : InMux
    port map (
            O => \N__33253\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500\
        );

    \I__3976\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33247\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__33247\,
            I => \N__33244\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__33244\,
            I => \N__33241\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__33241\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3251\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__3971\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33232\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__33232\,
            I => \N__33229\
        );

    \I__3969\ : Odrv12
    port map (
            O => \N__33229\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_CO\
        );

    \I__3968\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33223\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__33223\,
            I => \N__33220\
        );

    \I__3966\ : Span4Mux_v
    port map (
            O => \N__33220\,
            I => \N__33217\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__33217\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_44\
        );

    \I__3964\ : InMux
    port map (
            O => \N__33214\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501\
        );

    \I__3963\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33208\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__33208\,
            I => \N__33205\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__33205\,
            I => \N__33202\
        );

    \I__3960\ : Span4Mux_h
    port map (
            O => \N__33202\,
            I => \N__33199\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__33199\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3255\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__33196\,
            I => \N__33193\
        );

    \I__3957\ : InMux
    port map (
            O => \N__33193\,
            I => \N__33190\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__33190\,
            I => \N__33187\
        );

    \I__3955\ : Span4Mux_v
    port map (
            O => \N__33187\,
            I => \N__33184\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__33184\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_CO\
        );

    \I__3953\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33178\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__33178\,
            I => \N__33175\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__33175\,
            I => \N__33172\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__33172\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_45\
        );

    \I__3949\ : InMux
    port map (
            O => \N__33169\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502\
        );

    \I__3948\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33163\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__33160\,
            I => \N__33157\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__33157\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3259\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__33154\,
            I => \N__33151\
        );

    \I__3943\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__33148\,
            I => \N__33145\
        );

    \I__3941\ : Span4Mux_v
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__33142\,
            I => \N__33139\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__33139\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_CO\
        );

    \I__3938\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33133\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__33133\,
            I => \N__33130\
        );

    \I__3936\ : Span4Mux_v
    port map (
            O => \N__33130\,
            I => \N__33127\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__33127\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_46\
        );

    \I__3934\ : InMux
    port map (
            O => \N__33124\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503\
        );

    \I__3933\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33118\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33115\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__33115\,
            I => \N__33112\
        );

    \I__3930\ : Span4Mux_v
    port map (
            O => \N__33112\,
            I => \N__33109\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__33109\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3263\
        );

    \I__3928\ : InMux
    port map (
            O => \N__33106\,
            I => \N__33103\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__33103\,
            I => \N__33100\
        );

    \I__3926\ : Span4Mux_h
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__33097\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_CO\
        );

    \I__3924\ : InMux
    port map (
            O => \N__33094\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17504\
        );

    \I__3923\ : InMux
    port map (
            O => \N__33091\,
            I => \N__33088\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__33088\,
            I => \N__33085\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__33085\,
            I => \N__33082\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__33082\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_47\
        );

    \I__3919\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33076\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__33076\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2329\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__33073\,
            I => \N__33070\
        );

    \I__3916\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33067\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__33067\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2429\
        );

    \I__3914\ : InMux
    port map (
            O => \N__33064\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412\
        );

    \I__3913\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33058\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__33058\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2529\
        );

    \I__3911\ : InMux
    port map (
            O => \N__33055\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__33052\,
            I => \N__33049\
        );

    \I__3909\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33046\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__33046\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_CO\
        );

    \I__3907\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33040\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__33040\,
            I => \N__33037\
        );

    \I__3905\ : Odrv12
    port map (
            O => \N__33037\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_35\
        );

    \I__3904\ : InMux
    port map (
            O => \N__33034\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492\
        );

    \I__3903\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__33025\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__33025\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_36\
        );

    \I__3900\ : InMux
    port map (
            O => \N__33022\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493\
        );

    \I__3899\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33016\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__33016\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3223\
        );

    \I__3897\ : InMux
    port map (
            O => \N__33013\,
            I => \N__33010\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__3895\ : Odrv12
    port map (
            O => \N__33007\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_37\
        );

    \I__3894\ : InMux
    port map (
            O => \N__33004\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494\
        );

    \I__3893\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__3891\ : Span4Mux_v
    port map (
            O => \N__32995\,
            I => \N__32992\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__32992\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3227\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__32989\,
            I => \N__32986\
        );

    \I__3888\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32983\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__32983\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_CO\
        );

    \I__3886\ : InMux
    port map (
            O => \N__32980\,
            I => \N__32977\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__32971\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_38\
        );

    \I__3882\ : InMux
    port map (
            O => \N__32968\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__32965\,
            I => \N__32962\
        );

    \I__3880\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32959\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__32959\,
            I => \N__32956\
        );

    \I__3878\ : Span4Mux_v
    port map (
            O => \N__32956\,
            I => \N__32953\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__32953\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_CO\
        );

    \I__3876\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32947\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__32944\,
            I => \N__32941\
        );

    \I__3873\ : Odrv4
    port map (
            O => \N__32941\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_39\
        );

    \I__3872\ : InMux
    port map (
            O => \N__32938\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496\
        );

    \I__3871\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32932\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32929\
        );

    \I__3869\ : Odrv12
    port map (
            O => \N__32929\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_40\
        );

    \I__3868\ : InMux
    port map (
            O => \N__32926\,
            I => \bfn_11_20_0_\
        );

    \I__3867\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32917\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__32917\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3239\
        );

    \I__3864\ : InMux
    port map (
            O => \N__32914\,
            I => \N__32911\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__32911\,
            I => \N__32908\
        );

    \I__3862\ : Odrv12
    port map (
            O => \N__32908\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_41\
        );

    \I__3861\ : InMux
    port map (
            O => \N__32905\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498\
        );

    \I__3860\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32899\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__32899\,
            I => \N__32896\
        );

    \I__3858\ : Span4Mux_v
    port map (
            O => \N__32896\,
            I => \N__32893\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__32893\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3243\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__32890\,
            I => \N__32887\
        );

    \I__3855\ : InMux
    port map (
            O => \N__32887\,
            I => \N__32884\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__32884\,
            I => \N__32881\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__32881\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_CO\
        );

    \I__3852\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32875\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__32875\,
            I => \N__32872\
        );

    \I__3850\ : Odrv12
    port map (
            O => \N__32872\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_42\
        );

    \I__3849\ : InMux
    port map (
            O => \N__32869\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499\
        );

    \I__3848\ : InMux
    port map (
            O => \N__32866\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__32863\,
            I => \N__32857\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__32862\,
            I => \N__32853\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__32861\,
            I => \N__32849\
        );

    \I__3844\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32833\
        );

    \I__3843\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32833\
        );

    \I__3842\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32833\
        );

    \I__3841\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32833\
        );

    \I__3840\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32833\
        );

    \I__3839\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32833\
        );

    \I__3838\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32833\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__32833\,
            I => \N__32830\
        );

    \I__3836\ : Span4Mux_v
    port map (
            O => \N__32830\,
            I => \N__32827\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__32827\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2807\
        );

    \I__3834\ : InMux
    port map (
            O => \N__32824\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364\
        );

    \I__3833\ : InMux
    port map (
            O => \N__32821\,
            I => \bfn_11_18_0_\
        );

    \I__3832\ : InMux
    port map (
            O => \N__32818\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212\
        );

    \I__3831\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32812\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32809\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__32809\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3008\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__32806\,
            I => \N__32801\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__32805\,
            I => \N__32793\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__32804\,
            I => \N__32790\
        );

    \I__3825\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32787\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__32800\,
            I => \N__32784\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__32799\,
            I => \N__32780\
        );

    \I__3822\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32777\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__32797\,
            I => \N__32774\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__32796\,
            I => \N__32771\
        );

    \I__3819\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32767\
        );

    \I__3818\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32762\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32759\
        );

    \I__3816\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32756\
        );

    \I__3815\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32751\
        );

    \I__3814\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32751\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__32777\,
            I => \N__32748\
        );

    \I__3812\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32745\
        );

    \I__3811\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32742\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__32770\,
            I => \N__32739\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__32767\,
            I => \N__32735\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__32766\,
            I => \N__32732\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__32765\,
            I => \N__32729\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__32762\,
            I => \N__32725\
        );

    \I__3805\ : Span4Mux_v
    port map (
            O => \N__32759\,
            I => \N__32714\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__32756\,
            I => \N__32714\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__32751\,
            I => \N__32714\
        );

    \I__3802\ : Span4Mux_h
    port map (
            O => \N__32748\,
            I => \N__32714\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__32745\,
            I => \N__32714\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__32742\,
            I => \N__32711\
        );

    \I__3799\ : InMux
    port map (
            O => \N__32739\,
            I => \N__32708\
        );

    \I__3798\ : CascadeMux
    port map (
            O => \N__32738\,
            I => \N__32705\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__32735\,
            I => \N__32702\
        );

    \I__3796\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32697\
        );

    \I__3795\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32697\
        );

    \I__3794\ : InMux
    port map (
            O => \N__32728\,
            I => \N__32694\
        );

    \I__3793\ : Span4Mux_v
    port map (
            O => \N__32725\,
            I => \N__32688\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__32714\,
            I => \N__32688\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__32711\,
            I => \N__32683\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32683\
        );

    \I__3789\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32680\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__32702\,
            I => \N__32673\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__32697\,
            I => \N__32673\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__32694\,
            I => \N__32673\
        );

    \I__3785\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32670\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__32688\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__32683\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__32680\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__32673\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__32670\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\
        );

    \I__3779\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32656\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__32656\,
            I => \N__32653\
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__32653\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3108\
        );

    \I__3776\ : InMux
    port map (
            O => \N__32650\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490\
        );

    \I__3775\ : InMux
    port map (
            O => \N__32647\,
            I => \N__32644\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__32644\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3211\
        );

    \I__3773\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32638\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32635\
        );

    \I__3771\ : Odrv12
    port map (
            O => \N__32635\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_34\
        );

    \I__3770\ : InMux
    port map (
            O => \N__32632\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491\
        );

    \I__3769\ : InMux
    port map (
            O => \N__32629\,
            I => \foc.u_Park_Transform.n16959\
        );

    \I__3768\ : InMux
    port map (
            O => \N__32626\,
            I => \foc.u_Park_Transform.n16960\
        );

    \I__3767\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32620\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__32620\,
            I => \N__32616\
        );

    \I__3765\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32613\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__32616\,
            I => \foc.u_Park_Transform.n769\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__32613\,
            I => \foc.u_Park_Transform.n769\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__32608\,
            I => \N__32604\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__32607\,
            I => \N__32601\
        );

    \I__3760\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32597\
        );

    \I__3759\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32592\
        );

    \I__3758\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32592\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__32597\,
            I => \N__32587\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32587\
        );

    \I__3755\ : Odrv12
    port map (
            O => \N__32587\,
            I => \foc.u_Park_Transform.n617\
        );

    \I__3754\ : InMux
    port map (
            O => \N__32584\,
            I => \foc.u_Park_Transform.n16961\
        );

    \I__3753\ : InMux
    port map (
            O => \N__32581\,
            I => \foc.u_Park_Transform.n771\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__32578\,
            I => \N__32575\
        );

    \I__3751\ : InMux
    port map (
            O => \N__32575\,
            I => \N__32572\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__32572\,
            I => \N__32569\
        );

    \I__3749\ : Odrv12
    port map (
            O => \N__32569\,
            I => \foc.u_Park_Transform.n176_adj_2104\
        );

    \I__3748\ : InMux
    port map (
            O => \N__32566\,
            I => \foc.u_Park_Transform.n16950\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__32563\,
            I => \N__32560\
        );

    \I__3746\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32557\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__32557\,
            I => \N__32554\
        );

    \I__3744\ : Odrv12
    port map (
            O => \N__32554\,
            I => \foc.u_Park_Transform.n225_adj_2075\
        );

    \I__3743\ : InMux
    port map (
            O => \N__32551\,
            I => \foc.u_Park_Transform.n16951\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__32548\,
            I => \N__32545\
        );

    \I__3741\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32542\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32539\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__32539\,
            I => \foc.u_Park_Transform.n274_adj_2058\
        );

    \I__3738\ : InMux
    port map (
            O => \N__32536\,
            I => \foc.u_Park_Transform.n16952\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__32533\,
            I => \N__32530\
        );

    \I__3736\ : InMux
    port map (
            O => \N__32530\,
            I => \N__32527\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__32527\,
            I => \N__32524\
        );

    \I__3734\ : Odrv12
    port map (
            O => \N__32524\,
            I => \foc.u_Park_Transform.n323_adj_2057\
        );

    \I__3733\ : InMux
    port map (
            O => \N__32521\,
            I => \foc.u_Park_Transform.n16953\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__32518\,
            I => \N__32515\
        );

    \I__3731\ : InMux
    port map (
            O => \N__32515\,
            I => \N__32512\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32509\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__32509\,
            I => \foc.u_Park_Transform.n372_adj_2042\
        );

    \I__3728\ : InMux
    port map (
            O => \N__32506\,
            I => \foc.u_Park_Transform.n16954\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__32503\,
            I => \N__32500\
        );

    \I__3726\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32497\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__32497\,
            I => \N__32494\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__32494\,
            I => \N__32491\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__32491\,
            I => \foc.u_Park_Transform.n421\
        );

    \I__3722\ : InMux
    port map (
            O => \N__32488\,
            I => \bfn_11_16_0_\
        );

    \I__3721\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32482\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__32482\,
            I => \N__32479\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__32479\,
            I => \foc.u_Park_Transform.n470\
        );

    \I__3718\ : InMux
    port map (
            O => \N__32476\,
            I => \foc.u_Park_Transform.n16956\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__32473\,
            I => \N__32470\
        );

    \I__3716\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32467\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__32467\,
            I => \N__32464\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__32464\,
            I => \foc.u_Park_Transform.n519\
        );

    \I__3713\ : InMux
    port map (
            O => \N__32461\,
            I => \foc.u_Park_Transform.n16957\
        );

    \I__3712\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32455\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__32455\,
            I => \N__32452\
        );

    \I__3710\ : Odrv12
    port map (
            O => \N__32452\,
            I => \foc.u_Park_Transform.n568\
        );

    \I__3709\ : InMux
    port map (
            O => \N__32449\,
            I => \foc.u_Park_Transform.n16958\
        );

    \I__3708\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32440\
        );

    \I__3707\ : InMux
    port map (
            O => \N__32445\,
            I => \N__32440\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__32440\,
            I => \N__32437\
        );

    \I__3705\ : Odrv12
    port map (
            O => \N__32437\,
            I => \foc.Look_Up_Table_out1_1_11\
        );

    \I__3704\ : InMux
    port map (
            O => \N__32434\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952\
        );

    \I__3703\ : InMux
    port map (
            O => \N__32431\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953\
        );

    \I__3702\ : InMux
    port map (
            O => \N__32428\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954\
        );

    \I__3701\ : InMux
    port map (
            O => \N__32425\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955\
        );

    \I__3700\ : InMux
    port map (
            O => \N__32422\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15956\
        );

    \I__3699\ : InMux
    port map (
            O => \N__32419\,
            I => \N__32416\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32412\
        );

    \I__3697\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32409\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__32412\,
            I => \foc.Look_Up_Table_out1_1_12\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__32409\,
            I => \foc.Look_Up_Table_out1_1_12\
        );

    \I__3694\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32401\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__32401\,
            I => \N__32398\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__32398\,
            I => \N__32394\
        );

    \I__3691\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32391\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__32394\,
            I => \foc.u_Park_Transform.n785\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__32391\,
            I => \foc.u_Park_Transform.n785\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__32386\,
            I => \N__32377\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__32385\,
            I => \N__32373\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__32384\,
            I => \N__32360\
        );

    \I__3685\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32353\
        );

    \I__3684\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32353\
        );

    \I__3683\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32353\
        );

    \I__3682\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32343\
        );

    \I__3681\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32343\
        );

    \I__3680\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32343\
        );

    \I__3679\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32343\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__32372\,
            I => \N__32340\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__32371\,
            I => \N__32336\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__32370\,
            I => \N__32332\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__32369\,
            I => \N__32327\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__32368\,
            I => \N__32324\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__32367\,
            I => \N__32320\
        );

    \I__3672\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32307\
        );

    \I__3671\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32307\
        );

    \I__3670\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32307\
        );

    \I__3669\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32307\
        );

    \I__3668\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32307\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__32353\,
            I => \N__32304\
        );

    \I__3666\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32301\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32298\
        );

    \I__3664\ : InMux
    port map (
            O => \N__32340\,
            I => \N__32285\
        );

    \I__3663\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32285\
        );

    \I__3662\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32285\
        );

    \I__3661\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32285\
        );

    \I__3660\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32285\
        );

    \I__3659\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32285\
        );

    \I__3658\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32280\
        );

    \I__3657\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32280\
        );

    \I__3656\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32271\
        );

    \I__3655\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32271\
        );

    \I__3654\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32271\
        );

    \I__3653\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32271\
        );

    \I__3652\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32268\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32265\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__32304\,
            I => \N__32260\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__32301\,
            I => \N__32260\
        );

    \I__3648\ : Span4Mux_v
    port map (
            O => \N__32298\,
            I => \N__32249\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__32285\,
            I => \N__32249\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__32280\,
            I => \N__32249\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__32271\,
            I => \N__32249\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__32268\,
            I => \N__32249\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__32265\,
            I => \foc.u_Park_Transform.n616\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__32260\,
            I => \foc.u_Park_Transform.n616\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__32249\,
            I => \foc.u_Park_Transform.n616\
        );

    \I__3640\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32239\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32236\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__32236\,
            I => \foc.u_Park_Transform.n78_adj_2145\
        );

    \I__3637\ : InMux
    port map (
            O => \N__32233\,
            I => \foc.u_Park_Transform.n16948\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__32230\,
            I => \N__32227\
        );

    \I__3635\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32224\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32221\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__32221\,
            I => \foc.u_Park_Transform.n127_adj_2119\
        );

    \I__3632\ : InMux
    port map (
            O => \N__32218\,
            I => \foc.u_Park_Transform.n16949\
        );

    \I__3631\ : InMux
    port map (
            O => \N__32215\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944\
        );

    \I__3630\ : InMux
    port map (
            O => \N__32212\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945\
        );

    \I__3629\ : InMux
    port map (
            O => \N__32209\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946\
        );

    \I__3628\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32200\
        );

    \I__3627\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32200\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__32200\,
            I => \foc.Look_Up_Table_out1_1_6\
        );

    \I__3625\ : InMux
    port map (
            O => \N__32197\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947\
        );

    \I__3624\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32188\
        );

    \I__3623\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32188\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__32188\,
            I => \foc.Look_Up_Table_out1_1_7\
        );

    \I__3621\ : InMux
    port map (
            O => \N__32185\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948\
        );

    \I__3620\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32176\
        );

    \I__3619\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32176\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__32176\,
            I => \foc.Look_Up_Table_out1_1_8\
        );

    \I__3617\ : InMux
    port map (
            O => \N__32173\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949\
        );

    \I__3616\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32164\
        );

    \I__3615\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32164\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__32164\,
            I => \foc.Look_Up_Table_out1_1_9\
        );

    \I__3613\ : InMux
    port map (
            O => \N__32161\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950\
        );

    \I__3612\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32152\
        );

    \I__3611\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32152\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__32152\,
            I => \N__32149\
        );

    \I__3609\ : Odrv4
    port map (
            O => \N__32149\,
            I => \foc.Look_Up_Table_out1_1_10\
        );

    \I__3608\ : InMux
    port map (
            O => \N__32146\,
            I => \bfn_11_14_0_\
        );

    \I__3607\ : InMux
    port map (
            O => \N__32143\,
            I => \foc.u_Park_Transform.n787_adj_2149\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__32140\,
            I => \N__32137\
        );

    \I__3605\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32126\
        );

    \I__3604\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32126\
        );

    \I__3603\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32126\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__32134\,
            I => \N__32121\
        );

    \I__3601\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32118\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__32126\,
            I => \N__32110\
        );

    \I__3599\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32103\
        );

    \I__3598\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32103\
        );

    \I__3597\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32103\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__32118\,
            I => \N__32100\
        );

    \I__3595\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32097\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__32116\,
            I => \N__32094\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__32115\,
            I => \N__32090\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__32114\,
            I => \N__32086\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__32113\,
            I => \N__32083\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__32110\,
            I => \N__32078\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32078\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__32100\,
            I => \N__32073\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N__32073\
        );

    \I__3586\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32066\
        );

    \I__3585\ : InMux
    port map (
            O => \N__32093\,
            I => \N__32066\
        );

    \I__3584\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32066\
        );

    \I__3583\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32059\
        );

    \I__3582\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32059\
        );

    \I__3581\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32059\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__32078\,
            I => \foc.u_Park_Transform.n625\
        );

    \I__3579\ : Odrv4
    port map (
            O => \N__32073\,
            I => \foc.u_Park_Transform.n625\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__32066\,
            I => \foc.u_Park_Transform.n625\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__32059\,
            I => \foc.u_Park_Transform.n625\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__32050\,
            I => \n21486_cascade_\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__32047\,
            I => \N__32044\
        );

    \I__3574\ : InMux
    port map (
            O => \N__32044\,
            I => \N__32041\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__32041\,
            I => \N__32037\
        );

    \I__3572\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32034\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__32037\,
            I => n139
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__32034\,
            I => n139
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__32029\,
            I => \N__32026\
        );

    \I__3568\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32023\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__32023\,
            I => \N__32019\
        );

    \I__3566\ : InMux
    port map (
            O => \N__32022\,
            I => \N__32016\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__32019\,
            I => \foc.u_Park_Transform.n90\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__32016\,
            I => \foc.u_Park_Transform.n90\
        );

    \I__3563\ : InMux
    port map (
            O => \N__32011\,
            I => \N__32008\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__32008\,
            I => \N__32005\
        );

    \I__3561\ : Span4Mux_v
    port map (
            O => \N__32005\,
            I => \N__32001\
        );

    \I__3560\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31998\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__32001\,
            I => \foc.u_Park_Transform.n781\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__31998\,
            I => \foc.u_Park_Transform.n781\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__31993\,
            I => \N__31990\
        );

    \I__3556\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31987\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__31987\,
            I => \N__31984\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__31984\,
            I => \foc.u_Park_Transform.n87_adj_2138\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__31981\,
            I => \N__31978\
        );

    \I__3552\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31975\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__31975\,
            I => \N__31972\
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__31972\,
            I => \foc.u_Park_Transform.n136_adj_2127\
        );

    \I__3549\ : InMux
    port map (
            O => \N__31969\,
            I => \foc.u_Park_Transform.n17980\
        );

    \I__3548\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31963\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__31963\,
            I => \N__31960\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__31960\,
            I => \foc.u_Park_Transform.n185_adj_2126\
        );

    \I__3545\ : InMux
    port map (
            O => \N__31957\,
            I => \foc.u_Park_Transform.n17981\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__31954\,
            I => \N__31951\
        );

    \I__3543\ : InMux
    port map (
            O => \N__31951\,
            I => \N__31948\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__31948\,
            I => \N__31945\
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__31945\,
            I => \foc.u_Park_Transform.n234_adj_2125\
        );

    \I__3540\ : InMux
    port map (
            O => \N__31942\,
            I => \foc.u_Park_Transform.n17982\
        );

    \I__3539\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31936\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31933\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__31933\,
            I => \foc.u_Park_Transform.n283_adj_2122\
        );

    \I__3536\ : InMux
    port map (
            O => \N__31930\,
            I => \foc.u_Park_Transform.n17983\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__31927\,
            I => \N__31923\
        );

    \I__3534\ : InMux
    port map (
            O => \N__31926\,
            I => \N__31917\
        );

    \I__3533\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31917\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__31922\,
            I => \N__31914\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__31917\,
            I => \N__31911\
        );

    \I__3530\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31908\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__31911\,
            I => \foc.u_Park_Transform.n332_adj_2110\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__31908\,
            I => \foc.u_Park_Transform.n332_adj_2110\
        );

    \I__3527\ : InMux
    port map (
            O => \N__31903\,
            I => \foc.u_Park_Transform.n17984\
        );

    \I__3526\ : InMux
    port map (
            O => \N__31900\,
            I => \foc.u_Park_Transform.n17985\
        );

    \I__3525\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31894\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__31894\,
            I => \N__31891\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__31891\,
            I => \foc.u_Park_Transform.n182_adj_2094\
        );

    \I__3522\ : InMux
    port map (
            O => \N__31888\,
            I => \foc.u_Park_Transform.n17099\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__31885\,
            I => \N__31882\
        );

    \I__3520\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31879\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__31879\,
            I => \N__31876\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__31876\,
            I => \foc.u_Park_Transform.n231_adj_2089\
        );

    \I__3517\ : InMux
    port map (
            O => \N__31873\,
            I => \foc.u_Park_Transform.n17100\
        );

    \I__3516\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31867\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__31867\,
            I => \N__31864\
        );

    \I__3514\ : Span4Mux_v
    port map (
            O => \N__31864\,
            I => \N__31861\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__31861\,
            I => \foc.u_Park_Transform.n280_adj_2087\
        );

    \I__3512\ : InMux
    port map (
            O => \N__31858\,
            I => \foc.u_Park_Transform.n17101\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__31855\,
            I => \N__31852\
        );

    \I__3510\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31849\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31846\
        );

    \I__3508\ : Span4Mux_v
    port map (
            O => \N__31846\,
            I => \N__31843\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__31843\,
            I => \foc.u_Park_Transform.n329_adj_2080\
        );

    \I__3506\ : InMux
    port map (
            O => \N__31840\,
            I => \foc.u_Park_Transform.n17102\
        );

    \I__3505\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31834\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__3503\ : Odrv12
    port map (
            O => \N__31831\,
            I => \foc.u_Park_Transform.n378_adj_2078\
        );

    \I__3502\ : InMux
    port map (
            O => \N__31828\,
            I => \foc.u_Park_Transform.n17103\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__31825\,
            I => \N__31821\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__31824\,
            I => \N__31817\
        );

    \I__3499\ : InMux
    port map (
            O => \N__31821\,
            I => \N__31810\
        );

    \I__3498\ : InMux
    port map (
            O => \N__31820\,
            I => \N__31810\
        );

    \I__3497\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31810\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31807\
        );

    \I__3495\ : Span4Mux_h
    port map (
            O => \N__31807\,
            I => \N__31804\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__31804\,
            I => \foc.u_Park_Transform.n427_adj_2069\
        );

    \I__3493\ : InMux
    port map (
            O => \N__31801\,
            I => \foc.u_Park_Transform.n17104\
        );

    \I__3492\ : InMux
    port map (
            O => \N__31798\,
            I => \bfn_11_10_0_\
        );

    \I__3491\ : InMux
    port map (
            O => \N__31795\,
            I => \foc.u_Park_Transform.n783\
        );

    \I__3490\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31785\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__31791\,
            I => \N__31782\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__31790\,
            I => \N__31778\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__31789\,
            I => \N__31774\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__31788\,
            I => \N__31769\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__31785\,
            I => \N__31766\
        );

    \I__3484\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31753\
        );

    \I__3483\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31753\
        );

    \I__3482\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31753\
        );

    \I__3481\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31753\
        );

    \I__3480\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31753\
        );

    \I__3479\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31753\
        );

    \I__3478\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31748\
        );

    \I__3477\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31748\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__31766\,
            I => \N__31740\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__31753\,
            I => \N__31740\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__31748\,
            I => \N__31740\
        );

    \I__3473\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31737\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__31740\,
            I => \N__31730\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__31737\,
            I => \N__31727\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__31736\,
            I => \N__31724\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__31735\,
            I => \N__31720\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__31734\,
            I => \N__31716\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__31733\,
            I => \N__31711\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__31730\,
            I => \N__31706\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__31727\,
            I => \N__31706\
        );

    \I__3464\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31693\
        );

    \I__3463\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31693\
        );

    \I__3462\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31693\
        );

    \I__3461\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31693\
        );

    \I__3460\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31693\
        );

    \I__3459\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31693\
        );

    \I__3458\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31688\
        );

    \I__3457\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31688\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__31706\,
            I => \foc.u_Park_Transform.n622\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__31693\,
            I => \foc.u_Park_Transform.n622\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__31688\,
            I => \foc.u_Park_Transform.n622\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__31681\,
            I => \N__31678\
        );

    \I__3452\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31675\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__31675\,
            I => \N__31672\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__31672\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7552\
        );

    \I__3449\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31666\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__31666\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7470\
        );

    \I__3447\ : InMux
    port map (
            O => \N__31663\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352\
        );

    \I__3446\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31657\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__31657\,
            I => \N__31654\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__31654\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7551\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__31651\,
            I => \N__31648\
        );

    \I__3442\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31645\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__31645\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7469\
        );

    \I__3440\ : InMux
    port map (
            O => \N__31642\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353\
        );

    \I__3439\ : InMux
    port map (
            O => \N__31639\,
            I => \N__31636\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__31633\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7550\
        );

    \I__3436\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31627\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__31627\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7468\
        );

    \I__3434\ : InMux
    port map (
            O => \N__31624\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354\
        );

    \I__3433\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31618\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__31618\,
            I => \N__31615\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__31615\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7549\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__3429\ : InMux
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__31606\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7467\
        );

    \I__3427\ : InMux
    port map (
            O => \N__31603\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355\
        );

    \I__3426\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__31597\,
            I => \N__31594\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__31594\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7548\
        );

    \I__3423\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31588\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__31588\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7466\
        );

    \I__3421\ : InMux
    port map (
            O => \N__31585\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356\
        );

    \I__3420\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__31576\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7547\
        );

    \I__3417\ : CascadeMux
    port map (
            O => \N__31573\,
            I => \N__31564\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__31572\,
            I => \N__31558\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__31571\,
            I => \N__31555\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__31570\,
            I => \N__31551\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__31569\,
            I => \N__31548\
        );

    \I__3412\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31536\
        );

    \I__3411\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31536\
        );

    \I__3410\ : InMux
    port map (
            O => \N__31564\,
            I => \N__31536\
        );

    \I__3409\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31536\
        );

    \I__3408\ : InMux
    port map (
            O => \N__31562\,
            I => \N__31536\
        );

    \I__3407\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31529\
        );

    \I__3406\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31529\
        );

    \I__3405\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31529\
        );

    \I__3404\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31520\
        );

    \I__3403\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31520\
        );

    \I__3402\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31520\
        );

    \I__3401\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31520\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__31536\,
            I => \N__31511\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31511\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__31520\,
            I => \N__31511\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__31519\,
            I => \N__31506\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__31518\,
            I => \N__31502\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__31511\,
            I => \N__31488\
        );

    \I__3394\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31473\
        );

    \I__3393\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31473\
        );

    \I__3392\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31473\
        );

    \I__3391\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31473\
        );

    \I__3390\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31473\
        );

    \I__3389\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31473\
        );

    \I__3388\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31473\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__31499\,
            I => \N__31469\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__31498\,
            I => \N__31465\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__31497\,
            I => \N__31461\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__31496\,
            I => \N__31458\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__31495\,
            I => \N__31454\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__31494\,
            I => \N__31451\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__31493\,
            I => \N__31448\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__31492\,
            I => \N__31444\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__31491\,
            I => \N__31441\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__31488\,
            I => \N__31434\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__31473\,
            I => \N__31434\
        );

    \I__3376\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31419\
        );

    \I__3375\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31419\
        );

    \I__3374\ : InMux
    port map (
            O => \N__31468\,
            I => \N__31419\
        );

    \I__3373\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31419\
        );

    \I__3372\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31419\
        );

    \I__3371\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31419\
        );

    \I__3370\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31419\
        );

    \I__3369\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31416\
        );

    \I__3368\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31413\
        );

    \I__3367\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31406\
        );

    \I__3366\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31406\
        );

    \I__3365\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31406\
        );

    \I__3364\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31397\
        );

    \I__3363\ : InMux
    port map (
            O => \N__31441\,
            I => \N__31397\
        );

    \I__3362\ : InMux
    port map (
            O => \N__31440\,
            I => \N__31397\
        );

    \I__3361\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31397\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__31434\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__31419\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__31416\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__31413\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__31406\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__31397\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\
        );

    \I__3354\ : InMux
    port map (
            O => \N__31384\,
            I => \bfn_10_26_0_\
        );

    \I__3353\ : InMux
    port map (
            O => \N__31381\,
            I => \N__31378\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__31378\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7465\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__3350\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31369\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__31369\,
            I => \N__31366\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__31366\,
            I => \foc.u_Park_Transform.n84\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__31363\,
            I => \N__31360\
        );

    \I__3346\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31357\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__31357\,
            I => \N__31354\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__31354\,
            I => \foc.u_Park_Transform.n133_adj_2101\
        );

    \I__3343\ : InMux
    port map (
            O => \N__31351\,
            I => \foc.u_Park_Transform.n17098\
        );

    \I__3342\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31345\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__31345\,
            I => \N__31342\
        );

    \I__3340\ : Odrv12
    port map (
            O => \N__31342\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2920\
        );

    \I__3339\ : InMux
    port map (
            O => \N__31339\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__31336\,
            I => \N__31333\
        );

    \I__3337\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31330\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__31330\,
            I => \N__31327\
        );

    \I__3335\ : Odrv12
    port map (
            O => \N__31327\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3020\
        );

    \I__3334\ : InMux
    port map (
            O => \N__31324\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__31321\,
            I => \N__31315\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__31320\,
            I => \N__31311\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__31319\,
            I => \N__31307\
        );

    \I__3330\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31291\
        );

    \I__3329\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31291\
        );

    \I__3328\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31291\
        );

    \I__3327\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31291\
        );

    \I__3326\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31291\
        );

    \I__3325\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31291\
        );

    \I__3324\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31291\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31288\
        );

    \I__3322\ : Span4Mux_v
    port map (
            O => \N__31288\,
            I => \N__31284\
        );

    \I__3321\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31281\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__31284\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__31281\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819\
        );

    \I__3318\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31273\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__31273\,
            I => \N__31270\
        );

    \I__3316\ : Odrv12
    port map (
            O => \N__31270\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3120\
        );

    \I__3315\ : InMux
    port map (
            O => \N__31267\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400\
        );

    \I__3314\ : InMux
    port map (
            O => \N__31264\,
            I => \bfn_10_24_0_\
        );

    \I__3313\ : InMux
    port map (
            O => \N__31261\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228\
        );

    \I__3312\ : InMux
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__31255\,
            I => \N__31252\
        );

    \I__3310\ : Span4Mux_v
    port map (
            O => \N__31252\,
            I => \N__31249\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__31249\,
            I => \N__31246\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__31246\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7554\
        );

    \I__3307\ : InMux
    port map (
            O => \N__31243\,
            I => \N__31240\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__31240\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7472\
        );

    \I__3305\ : InMux
    port map (
            O => \N__31237\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__31234\,
            I => \N__31231\
        );

    \I__3303\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31228\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__31228\,
            I => \N__31225\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__31225\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7553\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__31222\,
            I => \N__31219\
        );

    \I__3299\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31216\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__31216\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7471\
        );

    \I__3297\ : InMux
    port map (
            O => \N__31213\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351\
        );

    \I__3296\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31207\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__31207\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2932\
        );

    \I__3294\ : InMux
    port map (
            O => \N__31204\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427\
        );

    \I__3293\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31198\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__31198\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3032\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__31195\,
            I => \N__31188\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__31194\,
            I => \N__31185\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__31193\,
            I => \N__31182\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__31192\,
            I => \N__31179\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__31191\,
            I => \N__31175\
        );

    \I__3286\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31170\
        );

    \I__3285\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31167\
        );

    \I__3284\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31154\
        );

    \I__3283\ : InMux
    port map (
            O => \N__31179\,
            I => \N__31154\
        );

    \I__3282\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31154\
        );

    \I__3281\ : InMux
    port map (
            O => \N__31175\,
            I => \N__31154\
        );

    \I__3280\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31154\
        );

    \I__3279\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31154\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__31170\,
            I => \N__31147\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31147\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__31154\,
            I => \N__31147\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__31147\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2828\
        );

    \I__3274\ : InMux
    port map (
            O => \N__31144\,
            I => \bfn_10_22_0_\
        );

    \I__3273\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31138\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__31138\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3132\
        );

    \I__3271\ : InMux
    port map (
            O => \N__31135\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429\
        );

    \I__3270\ : InMux
    port map (
            O => \N__31132\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__31129\,
            I => \N__31126\
        );

    \I__3268\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31123\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__31123\,
            I => \N__31120\
        );

    \I__3266\ : Span12Mux_h
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__3265\ : Odrv12
    port map (
            O => \N__31117\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2420\
        );

    \I__3264\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31111\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__31111\,
            I => \N__31108\
        );

    \I__3262\ : Span4Mux_v
    port map (
            O => \N__31108\,
            I => \N__31105\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__31105\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2520\
        );

    \I__3260\ : InMux
    port map (
            O => \N__31102\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__31099\,
            I => \N__31096\
        );

    \I__3258\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31093\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31090\
        );

    \I__3256\ : Span4Mux_v
    port map (
            O => \N__31090\,
            I => \N__31087\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__31087\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2620\
        );

    \I__3254\ : InMux
    port map (
            O => \N__31084\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395\
        );

    \I__3253\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31078\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__31078\,
            I => \N__31075\
        );

    \I__3251\ : Odrv12
    port map (
            O => \N__31075\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2720\
        );

    \I__3250\ : InMux
    port map (
            O => \N__31072\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__31069\,
            I => \N__31066\
        );

    \I__3248\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31063\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__31063\,
            I => \N__31060\
        );

    \I__3246\ : Odrv12
    port map (
            O => \N__31060\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2820\
        );

    \I__3245\ : InMux
    port map (
            O => \N__31057\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397\
        );

    \I__3244\ : InMux
    port map (
            O => \N__31054\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224\
        );

    \I__3243\ : InMux
    port map (
            O => \N__31051\,
            I => \N__31048\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__31048\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2332\
        );

    \I__3241\ : InMux
    port map (
            O => \N__31045\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__31042\,
            I => \N__31039\
        );

    \I__3239\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31036\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__31036\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2432\
        );

    \I__3237\ : InMux
    port map (
            O => \N__31033\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422\
        );

    \I__3236\ : InMux
    port map (
            O => \N__31030\,
            I => \N__31027\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__31027\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2532\
        );

    \I__3234\ : InMux
    port map (
            O => \N__31024\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__3232\ : InMux
    port map (
            O => \N__31018\,
            I => \N__31015\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__31015\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2632\
        );

    \I__3230\ : InMux
    port map (
            O => \N__31012\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424\
        );

    \I__3229\ : InMux
    port map (
            O => \N__31009\,
            I => \N__31006\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__31006\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2732\
        );

    \I__3227\ : InMux
    port map (
            O => \N__31003\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425\
        );

    \I__3226\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30997\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__30997\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2832\
        );

    \I__3224\ : InMux
    port map (
            O => \N__30994\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426\
        );

    \I__3223\ : InMux
    port map (
            O => \N__30991\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385\
        );

    \I__3222\ : InMux
    port map (
            O => \N__30988\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386\
        );

    \I__3221\ : InMux
    port map (
            O => \N__30985\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387\
        );

    \I__3220\ : InMux
    port map (
            O => \N__30982\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388\
        );

    \I__3219\ : InMux
    port map (
            O => \N__30979\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389\
        );

    \I__3218\ : InMux
    port map (
            O => \N__30976\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390\
        );

    \I__3217\ : InMux
    port map (
            O => \N__30973\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391\
        );

    \I__3216\ : InMux
    port map (
            O => \N__30970\,
            I => \bfn_10_20_0_\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__30967\,
            I => \N__30964\
        );

    \I__3214\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30961\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30958\
        );

    \I__3212\ : Odrv12
    port map (
            O => \N__30958\,
            I => \foc.u_Park_Transform.n231\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__30955\,
            I => \N__30952\
        );

    \I__3210\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30949\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__30949\,
            I => \N__30946\
        );

    \I__3208\ : Span4Mux_v
    port map (
            O => \N__30946\,
            I => \N__30943\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__30943\,
            I => \foc.u_Park_Transform.n277\
        );

    \I__3206\ : InMux
    port map (
            O => \N__30940\,
            I => \foc.u_Park_Transform.n16927\
        );

    \I__3205\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30934\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__30934\,
            I => \N__30931\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__30931\,
            I => \foc.u_Park_Transform.n280\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__30928\,
            I => \N__30925\
        );

    \I__3201\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30922\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__30922\,
            I => \N__30919\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__30919\,
            I => \foc.u_Park_Transform.n326\
        );

    \I__3198\ : InMux
    port map (
            O => \N__30916\,
            I => \foc.u_Park_Transform.n16928\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__30913\,
            I => \N__30910\
        );

    \I__3196\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30907\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__30904\,
            I => \foc.u_Park_Transform.n329\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__30901\,
            I => \N__30898\
        );

    \I__3192\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30895\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30892\
        );

    \I__3190\ : Span4Mux_v
    port map (
            O => \N__30892\,
            I => \N__30889\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__30889\,
            I => \foc.u_Park_Transform.n375\
        );

    \I__3188\ : InMux
    port map (
            O => \N__30886\,
            I => \foc.u_Park_Transform.n16929\
        );

    \I__3187\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30880\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30877\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__30877\,
            I => \foc.u_Park_Transform.n378\
        );

    \I__3184\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30871\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__30871\,
            I => \foc.u_Park_Transform.n424\
        );

    \I__3182\ : InMux
    port map (
            O => \N__30868\,
            I => \foc.u_Park_Transform.n16930\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__30865\,
            I => \N__30862\
        );

    \I__3180\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30859\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__30856\,
            I => \foc.u_Park_Transform.n473\
        );

    \I__3177\ : InMux
    port map (
            O => \N__30853\,
            I => \bfn_10_18_0_\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__30850\,
            I => \N__30841\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \N__30834\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__30848\,
            I => \N__30830\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__30847\,
            I => \N__30826\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__30846\,
            I => \N__30822\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__30845\,
            I => \N__30817\
        );

    \I__3170\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30812\
        );

    \I__3169\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30812\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__30840\,
            I => \N__30809\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__30839\,
            I => \N__30805\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__30838\,
            I => \N__30801\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__30837\,
            I => \N__30797\
        );

    \I__3164\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30791\
        );

    \I__3163\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30791\
        );

    \I__3162\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30778\
        );

    \I__3161\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30778\
        );

    \I__3160\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30778\
        );

    \I__3159\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30778\
        );

    \I__3158\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30778\
        );

    \I__3157\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30778\
        );

    \I__3156\ : InMux
    port map (
            O => \N__30820\,
            I => \N__30773\
        );

    \I__3155\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30773\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__30812\,
            I => \N__30770\
        );

    \I__3153\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30765\
        );

    \I__3152\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30765\
        );

    \I__3151\ : InMux
    port map (
            O => \N__30805\,
            I => \N__30751\
        );

    \I__3150\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30751\
        );

    \I__3149\ : InMux
    port map (
            O => \N__30801\,
            I => \N__30751\
        );

    \I__3148\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30751\
        );

    \I__3147\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30751\
        );

    \I__3146\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30751\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__30791\,
            I => \N__30748\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30743\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__30773\,
            I => \N__30743\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__30770\,
            I => \N__30738\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30738\
        );

    \I__3140\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30735\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30731\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__30748\,
            I => \N__30722\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__30743\,
            I => \N__30722\
        );

    \I__3136\ : Span4Mux_h
    port map (
            O => \N__30738\,
            I => \N__30722\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30722\
        );

    \I__3134\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30719\
        );

    \I__3133\ : Odrv12
    port map (
            O => \N__30731\,
            I => \foc.u_Park_Transform.n619\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__30722\,
            I => \foc.u_Park_Transform.n619\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__30719\,
            I => \foc.u_Park_Transform.n619\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__30712\,
            I => \N__30708\
        );

    \I__3129\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30700\
        );

    \I__3128\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30700\
        );

    \I__3127\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30700\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__30700\,
            I => \N__30697\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__30697\,
            I => \foc.u_Park_Transform.n522\
        );

    \I__3124\ : InMux
    port map (
            O => \N__30694\,
            I => \foc.u_Park_Transform.n16932\
        );

    \I__3123\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30688\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__30688\,
            I => \N__30684\
        );

    \I__3121\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30681\
        );

    \I__3120\ : Span12Mux_h
    port map (
            O => \N__30684\,
            I => \N__30676\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30676\
        );

    \I__3118\ : Odrv12
    port map (
            O => \N__30676\,
            I => \foc.u_Park_Transform.n777\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__30673\,
            I => \N__30669\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__30672\,
            I => \N__30665\
        );

    \I__3115\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30658\
        );

    \I__3114\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30658\
        );

    \I__3113\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30658\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N__30655\
        );

    \I__3111\ : Odrv12
    port map (
            O => \N__30655\,
            I => \foc.u_Park_Transform.n427\
        );

    \I__3110\ : InMux
    port map (
            O => \N__30652\,
            I => \foc.u_Park_Transform.n16933\
        );

    \I__3109\ : InMux
    port map (
            O => \N__30649\,
            I => \foc.u_Park_Transform.n779\
        );

    \I__3108\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30643\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__30643\,
            I => \foc.u_Park_Transform.n283\
        );

    \I__3106\ : InMux
    port map (
            O => \N__30640\,
            I => \foc.u_Park_Transform.n16919\
        );

    \I__3105\ : InMux
    port map (
            O => \N__30637\,
            I => \foc.u_Park_Transform.n16920\
        );

    \I__3104\ : InMux
    port map (
            O => \N__30634\,
            I => \foc.u_Park_Transform.n16921\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__30631\,
            I => \N__30628\
        );

    \I__3102\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30624\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__30627\,
            I => \N__30620\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__30624\,
            I => \N__30617\
        );

    \I__3099\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30612\
        );

    \I__3098\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30612\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__30617\,
            I => \foc.u_Park_Transform.n332\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__30612\,
            I => \foc.u_Park_Transform.n332\
        );

    \I__3095\ : InMux
    port map (
            O => \N__30607\,
            I => \bfn_10_16_0_\
        );

    \I__3094\ : InMux
    port map (
            O => \N__30604\,
            I => \foc.u_Park_Transform.n783_adj_2167\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__30601\,
            I => \N__30598\
        );

    \I__3092\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30595\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__30595\,
            I => \N__30592\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__30592\,
            I => \foc.u_Park_Transform.n81_adj_2120\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__30589\,
            I => \N__30586\
        );

    \I__3088\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30583\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__30583\,
            I => \N__30580\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__30580\,
            I => \foc.u_Park_Transform.n84_adj_2118\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__30577\,
            I => \N__30574\
        );

    \I__3084\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30571\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30568\
        );

    \I__3082\ : Span4Mux_h
    port map (
            O => \N__30568\,
            I => \N__30565\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__30565\,
            I => \foc.u_Park_Transform.n130_adj_2105\
        );

    \I__3080\ : InMux
    port map (
            O => \N__30562\,
            I => \foc.u_Park_Transform.n16924\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__30559\,
            I => \N__30556\
        );

    \I__3078\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30553\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__30553\,
            I => \N__30550\
        );

    \I__3076\ : Odrv12
    port map (
            O => \N__30550\,
            I => \foc.u_Park_Transform.n133\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__30547\,
            I => \N__30544\
        );

    \I__3074\ : InMux
    port map (
            O => \N__30544\,
            I => \N__30541\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__30541\,
            I => \N__30538\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__30538\,
            I => \foc.u_Park_Transform.n179_adj_2076\
        );

    \I__3071\ : InMux
    port map (
            O => \N__30535\,
            I => \foc.u_Park_Transform.n16925\
        );

    \I__3070\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30529\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30526\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__30526\,
            I => \foc.u_Park_Transform.n182\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__30523\,
            I => \N__30520\
        );

    \I__3066\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30517\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30514\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__30514\,
            I => \foc.u_Park_Transform.n228\
        );

    \I__3063\ : InMux
    port map (
            O => \N__30511\,
            I => \foc.u_Park_Transform.n16926\
        );

    \I__3062\ : InMux
    port map (
            O => \N__30508\,
            I => \foc.u_Park_Transform.n18164\
        );

    \I__3061\ : InMux
    port map (
            O => \N__30505\,
            I => \foc.u_Park_Transform.n18165\
        );

    \I__3060\ : InMux
    port map (
            O => \N__30502\,
            I => \foc.u_Park_Transform.n787\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__30499\,
            I => \N__30496\
        );

    \I__3058\ : InMux
    port map (
            O => \N__30496\,
            I => \N__30493\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__30493\,
            I => \foc.u_Park_Transform.n87\
        );

    \I__3056\ : InMux
    port map (
            O => \N__30490\,
            I => \foc.u_Park_Transform.n16915\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__30487\,
            I => \N__30484\
        );

    \I__3054\ : InMux
    port map (
            O => \N__30484\,
            I => \N__30481\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__30481\,
            I => \foc.u_Park_Transform.n136\
        );

    \I__3052\ : InMux
    port map (
            O => \N__30478\,
            I => \foc.u_Park_Transform.n16916\
        );

    \I__3051\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30472\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__30472\,
            I => \foc.u_Park_Transform.n185\
        );

    \I__3049\ : InMux
    port map (
            O => \N__30469\,
            I => \foc.u_Park_Transform.n16917\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__30466\,
            I => \N__30463\
        );

    \I__3047\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30460\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__30460\,
            I => \foc.u_Park_Transform.n234\
        );

    \I__3045\ : InMux
    port map (
            O => \N__30457\,
            I => \foc.u_Park_Transform.n16918\
        );

    \I__3044\ : InMux
    port map (
            O => \N__30454\,
            I => \foc.u_Park_Transform.n771_adj_2032\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__30451\,
            I => \N__30448\
        );

    \I__3042\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30444\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__30447\,
            I => \N__30441\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__30444\,
            I => \N__30438\
        );

    \I__3039\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30435\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__30438\,
            I => \foc.u_Park_Transform.n773\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__30435\,
            I => \foc.u_Park_Transform.n773\
        );

    \I__3036\ : InMux
    port map (
            O => \N__30430\,
            I => \foc.u_Park_Transform.n18160\
        );

    \I__3035\ : InMux
    port map (
            O => \N__30427\,
            I => \foc.u_Park_Transform.n18161\
        );

    \I__3034\ : InMux
    port map (
            O => \N__30424\,
            I => \foc.u_Park_Transform.n18162\
        );

    \I__3033\ : InMux
    port map (
            O => \N__30421\,
            I => \foc.u_Park_Transform.n18163\
        );

    \I__3032\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30415\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__30415\,
            I => \foc.u_Park_Transform.n372\
        );

    \I__3030\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30409\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__30409\,
            I => \foc.u_Park_Transform.n418_adj_2024\
        );

    \I__3028\ : InMux
    port map (
            O => \N__30406\,
            I => \foc.u_Park_Transform.n17137\
        );

    \I__3027\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30400\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__30400\,
            I => \foc.u_Park_Transform.n421_adj_2039\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__30397\,
            I => \N__30394\
        );

    \I__3024\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30391\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__30391\,
            I => \N__30388\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__30388\,
            I => \foc.u_Park_Transform.n467_adj_2019\
        );

    \I__3021\ : InMux
    port map (
            O => \N__30385\,
            I => \bfn_10_12_0_\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__30382\,
            I => \N__30379\
        );

    \I__3019\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30376\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__30376\,
            I => \foc.u_Park_Transform.n470_adj_2038\
        );

    \I__3017\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30370\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__30370\,
            I => \N__30367\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__30367\,
            I => \foc.u_Park_Transform.n516_adj_2018\
        );

    \I__3014\ : InMux
    port map (
            O => \N__30364\,
            I => \foc.u_Park_Transform.n17139\
        );

    \I__3013\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30358\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__30358\,
            I => \foc.u_Park_Transform.n519_adj_2035\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__30355\,
            I => \N__30352\
        );

    \I__3010\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30349\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__30349\,
            I => \N__30346\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__30346\,
            I => \foc.u_Park_Transform.n565\
        );

    \I__3007\ : InMux
    port map (
            O => \N__30343\,
            I => \foc.u_Park_Transform.n17140\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__30340\,
            I => \N__30337\
        );

    \I__3005\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30334\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__30334\,
            I => \foc.u_Park_Transform.n568_adj_2034\
        );

    \I__3003\ : InMux
    port map (
            O => \N__30331\,
            I => \N__30328\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__30328\,
            I => \N__30325\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__30325\,
            I => \foc.u_Park_Transform.n614_adj_2017\
        );

    \I__3000\ : InMux
    port map (
            O => \N__30322\,
            I => \foc.u_Park_Transform.n17141\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__30319\,
            I => \N__30316\
        );

    \I__2998\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30313\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30310\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__30310\,
            I => \foc.u_Park_Transform.n663_adj_2016\
        );

    \I__2995\ : InMux
    port map (
            O => \N__30307\,
            I => \foc.u_Park_Transform.n17142\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__30304\,
            I => \N__30301\
        );

    \I__2993\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30298\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__30298\,
            I => \N__30295\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__30295\,
            I => \foc.u_Park_Transform.n712_adj_2015\
        );

    \I__2990\ : InMux
    port map (
            O => \N__30292\,
            I => \foc.u_Park_Transform.n17143\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__30289\,
            I => \N__30285\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__30288\,
            I => \N__30282\
        );

    \I__2987\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30278\
        );

    \I__2986\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30273\
        );

    \I__2985\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30273\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__30278\,
            I => \foc.u_Park_Transform.n617_adj_2031\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__30273\,
            I => \foc.u_Park_Transform.n617_adj_2031\
        );

    \I__2982\ : InMux
    port map (
            O => \N__30268\,
            I => \foc.u_Park_Transform.n17144\
        );

    \I__2981\ : InMux
    port map (
            O => \N__30265\,
            I => \foc.u_Park_Transform.n767\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__30262\,
            I => \N__30259\
        );

    \I__2979\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30256\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__30256\,
            I => \N__30253\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__30253\,
            I => \foc.u_Park_Transform.n75\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__30250\,
            I => \N__30247\
        );

    \I__2975\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30244\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__30244\,
            I => \foc.u_Park_Transform.n78\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__30241\,
            I => \N__30238\
        );

    \I__2972\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30235\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30232\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__30232\,
            I => \foc.u_Park_Transform.n124\
        );

    \I__2969\ : InMux
    port map (
            O => \N__30229\,
            I => \foc.u_Park_Transform.n17131\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__2967\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__30220\,
            I => \foc.u_Park_Transform.n127\
        );

    \I__2965\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30214\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__30214\,
            I => \N__30211\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__30211\,
            I => \foc.u_Park_Transform.n173\
        );

    \I__2962\ : InMux
    port map (
            O => \N__30208\,
            I => \foc.u_Park_Transform.n17132\
        );

    \I__2961\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__30202\,
            I => \foc.u_Park_Transform.n176\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__30199\,
            I => \N__30196\
        );

    \I__2958\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30190\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__30190\,
            I => \foc.u_Park_Transform.n222\
        );

    \I__2955\ : InMux
    port map (
            O => \N__30187\,
            I => \foc.u_Park_Transform.n17133\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__30184\,
            I => \N__30181\
        );

    \I__2953\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__30178\,
            I => \foc.u_Park_Transform.n225\
        );

    \I__2951\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30172\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30169\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__30169\,
            I => \foc.u_Park_Transform.n271\
        );

    \I__2948\ : InMux
    port map (
            O => \N__30166\,
            I => \foc.u_Park_Transform.n17134\
        );

    \I__2947\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__30160\,
            I => \foc.u_Park_Transform.n274\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__2944\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30151\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__30151\,
            I => \N__30148\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__30148\,
            I => \foc.u_Park_Transform.n320\
        );

    \I__2941\ : InMux
    port map (
            O => \N__30145\,
            I => \foc.u_Park_Transform.n17135\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__30142\,
            I => \N__30139\
        );

    \I__2939\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30136\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__30136\,
            I => \foc.u_Park_Transform.n323\
        );

    \I__2937\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30130\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__30130\,
            I => \N__30127\
        );

    \I__2935\ : Odrv12
    port map (
            O => \N__30127\,
            I => \foc.u_Park_Transform.n369\
        );

    \I__2934\ : InMux
    port map (
            O => \N__30124\,
            I => \foc.u_Park_Transform.n17136\
        );

    \I__2933\ : InMux
    port map (
            O => \N__30121\,
            I => \foc.u_Park_Transform.n17151\
        );

    \I__2932\ : InMux
    port map (
            O => \N__30118\,
            I => \foc.u_Park_Transform.n17152\
        );

    \I__2931\ : InMux
    port map (
            O => \N__30115\,
            I => \bfn_10_10_0_\
        );

    \I__2930\ : InMux
    port map (
            O => \N__30112\,
            I => \foc.u_Park_Transform.n17154\
        );

    \I__2929\ : InMux
    port map (
            O => \N__30109\,
            I => \foc.u_Park_Transform.n17155\
        );

    \I__2928\ : InMux
    port map (
            O => \N__30106\,
            I => \foc.u_Park_Transform.n17156\
        );

    \I__2927\ : InMux
    port map (
            O => \N__30103\,
            I => \foc.u_Park_Transform.n17157\
        );

    \I__2926\ : InMux
    port map (
            O => \N__30100\,
            I => \foc.u_Park_Transform.n17158\
        );

    \I__2925\ : InMux
    port map (
            O => \N__30097\,
            I => \foc.u_Park_Transform.n17159\
        );

    \I__2924\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30091\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30088\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__30088\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3047\
        );

    \I__2921\ : InMux
    port map (
            O => \N__30085\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487\
        );

    \I__2920\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30079\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__30079\,
            I => \N__30076\
        );

    \I__2918\ : Span4Mux_v
    port map (
            O => \N__30076\,
            I => \N__30073\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__30073\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3147\
        );

    \I__2916\ : InMux
    port map (
            O => \N__30070\,
            I => \bfn_9_25_0_\
        );

    \I__2915\ : InMux
    port map (
            O => \N__30067\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17489\
        );

    \I__2914\ : InMux
    port map (
            O => \N__30064\,
            I => \foc.u_Park_Transform.n17146\
        );

    \I__2913\ : InMux
    port map (
            O => \N__30061\,
            I => \foc.u_Park_Transform.n17147\
        );

    \I__2912\ : InMux
    port map (
            O => \N__30058\,
            I => \foc.u_Park_Transform.n17148\
        );

    \I__2911\ : InMux
    port map (
            O => \N__30055\,
            I => \foc.u_Park_Transform.n17149\
        );

    \I__2910\ : InMux
    port map (
            O => \N__30052\,
            I => \foc.u_Park_Transform.n17150\
        );

    \I__2909\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__30046\,
            I => \N__30043\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__30043\,
            I => \N__30040\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__30040\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7891\
        );

    \I__2905\ : InMux
    port map (
            O => \N__30037\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17343\
        );

    \I__2904\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__30028\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__30028\,
            I => \N__30025\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__30025\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2347\
        );

    \I__2900\ : InMux
    port map (
            O => \N__30022\,
            I => \N__30019\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__30019\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7473\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__30016\,
            I => \N__30013\
        );

    \I__2897\ : InMux
    port map (
            O => \N__30013\,
            I => \N__30010\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__30010\,
            I => \N__30007\
        );

    \I__2895\ : Span4Mux_v
    port map (
            O => \N__30007\,
            I => \N__30004\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__30004\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2447\
        );

    \I__2893\ : InMux
    port map (
            O => \N__30001\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481\
        );

    \I__2892\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29995\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__29995\,
            I => \N__29992\
        );

    \I__2890\ : Span4Mux_h
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__29989\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2547\
        );

    \I__2888\ : InMux
    port map (
            O => \N__29986\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__29983\,
            I => \N__29980\
        );

    \I__2886\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29977\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__29977\,
            I => \N__29974\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__29974\,
            I => \N__29971\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__29971\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2647\
        );

    \I__2882\ : InMux
    port map (
            O => \N__29968\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483\
        );

    \I__2881\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29962\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__29962\,
            I => \N__29959\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__29959\,
            I => \N__29956\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__29956\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2747\
        );

    \I__2877\ : InMux
    port map (
            O => \N__29953\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484\
        );

    \I__2876\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29947\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__29947\,
            I => \N__29944\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__29944\,
            I => \N__29941\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__29941\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2847\
        );

    \I__2872\ : InMux
    port map (
            O => \N__29938\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485\
        );

    \I__2871\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29932\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__29932\,
            I => \N__29929\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__29929\,
            I => \N__29926\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__29926\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2947\
        );

    \I__2867\ : InMux
    port map (
            O => \N__29923\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486\
        );

    \I__2866\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29917\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__29917\,
            I => \N__29914\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__29914\,
            I => \N__29911\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__29911\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3135\
        );

    \I__2862\ : InMux
    port map (
            O => \N__29908\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439\
        );

    \I__2861\ : InMux
    port map (
            O => \N__29905\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244\
        );

    \I__2860\ : InMux
    port map (
            O => \N__29902\,
            I => \N__29899\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__29899\,
            I => \N__29896\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__29896\,
            I => \N__29893\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__29893\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7897\
        );

    \I__2856\ : InMux
    port map (
            O => \N__29890\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29884\
        );

    \I__2854\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29881\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29878\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__29878\,
            I => \N__29875\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__29875\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7896\
        );

    \I__2850\ : InMux
    port map (
            O => \N__29872\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338\
        );

    \I__2849\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29866\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29863\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__29863\,
            I => \N__29860\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__29860\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7895\
        );

    \I__2845\ : InMux
    port map (
            O => \N__29857\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__29854\,
            I => \N__29851\
        );

    \I__2843\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29848\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__29848\,
            I => \N__29845\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__29845\,
            I => \N__29842\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__29842\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7894\
        );

    \I__2839\ : InMux
    port map (
            O => \N__29839\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340\
        );

    \I__2838\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29833\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N__29830\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__29830\,
            I => \N__29827\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__29827\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7893\
        );

    \I__2834\ : InMux
    port map (
            O => \N__29824\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__29821\,
            I => \N__29818\
        );

    \I__2832\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29815\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__29815\,
            I => \N__29812\
        );

    \I__2830\ : Span12Mux_s11_v
    port map (
            O => \N__29812\,
            I => \N__29809\
        );

    \I__2829\ : Odrv12
    port map (
            O => \N__29809\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7892\
        );

    \I__2828\ : InMux
    port map (
            O => \N__29806\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342\
        );

    \I__2827\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29800\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__29800\,
            I => \N__29797\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__29797\,
            I => \N__29794\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__29794\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2335\
        );

    \I__2823\ : InMux
    port map (
            O => \N__29791\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431\
        );

    \I__2822\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29785\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__29785\,
            I => \N__29782\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__29782\,
            I => \N__29779\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__29779\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2435\
        );

    \I__2818\ : InMux
    port map (
            O => \N__29776\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__29773\,
            I => \N__29770\
        );

    \I__2816\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29767\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29764\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__29764\,
            I => \N__29761\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__29761\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2535\
        );

    \I__2812\ : InMux
    port map (
            O => \N__29758\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433\
        );

    \I__2811\ : InMux
    port map (
            O => \N__29755\,
            I => \N__29752\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__29752\,
            I => \N__29749\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__29746\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2635\
        );

    \I__2807\ : InMux
    port map (
            O => \N__29743\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__29740\,
            I => \N__29737\
        );

    \I__2805\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29734\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__29734\,
            I => \N__29731\
        );

    \I__2803\ : Span4Mux_v
    port map (
            O => \N__29731\,
            I => \N__29728\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__29728\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2735\
        );

    \I__2801\ : InMux
    port map (
            O => \N__29725\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435\
        );

    \I__2800\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29719\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N__29716\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__29716\,
            I => \N__29713\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__29713\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2835\
        );

    \I__2796\ : InMux
    port map (
            O => \N__29710\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436\
        );

    \I__2795\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29704\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29701\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__29701\,
            I => \N__29698\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__29698\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2935\
        );

    \I__2791\ : InMux
    port map (
            O => \N__29695\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437\
        );

    \I__2790\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29689\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__29689\,
            I => \N__29686\
        );

    \I__2788\ : Span4Mux_h
    port map (
            O => \N__29686\,
            I => \N__29683\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__29683\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3035\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__2785\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29669\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \N__29666\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__29675\,
            I => \N__29663\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__29674\,
            I => \N__29659\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \N__29655\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__29672\,
            I => \N__29652\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__29669\,
            I => \N__29649\
        );

    \I__2778\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29646\
        );

    \I__2777\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29633\
        );

    \I__2776\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29633\
        );

    \I__2775\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29633\
        );

    \I__2774\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29633\
        );

    \I__2773\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29633\
        );

    \I__2772\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29633\
        );

    \I__2771\ : Odrv12
    port map (
            O => \N__29649\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__29646\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__29633\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831\
        );

    \I__2768\ : InMux
    port map (
            O => \N__29626\,
            I => \bfn_9_22_0_\
        );

    \I__2767\ : InMux
    port map (
            O => \N__29623\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464\
        );

    \I__2766\ : InMux
    port map (
            O => \N__29620\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465\
        );

    \I__2765\ : InMux
    port map (
            O => \N__29617\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466\
        );

    \I__2764\ : InMux
    port map (
            O => \N__29614\,
            I => \bfn_9_20_0_\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__29611\,
            I => \N__29606\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__29610\,
            I => \N__29602\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__29609\,
            I => \N__29598\
        );

    \I__2760\ : InMux
    port map (
            O => \N__29606\,
            I => \N__29580\
        );

    \I__2759\ : InMux
    port map (
            O => \N__29605\,
            I => \N__29580\
        );

    \I__2758\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29580\
        );

    \I__2757\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29580\
        );

    \I__2756\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29580\
        );

    \I__2755\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29580\
        );

    \I__2754\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29580\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__29595\,
            I => \N__29577\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__29580\,
            I => \N__29574\
        );

    \I__2751\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29571\
        );

    \I__2750\ : Span4Mux_v
    port map (
            O => \N__29574\,
            I => \N__29566\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__29571\,
            I => \N__29566\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__29566\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2834\
        );

    \I__2747\ : InMux
    port map (
            O => \N__29563\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__29560\,
            I => \N__29557\
        );

    \I__2745\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29554\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__29554\,
            I => \N__29548\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__29553\,
            I => \N__29544\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__29552\,
            I => \N__29540\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__29551\,
            I => \N__29536\
        );

    \I__2740\ : Span4Mux_h
    port map (
            O => \N__29548\,
            I => \N__29528\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29525\
        );

    \I__2738\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29510\
        );

    \I__2737\ : InMux
    port map (
            O => \N__29543\,
            I => \N__29510\
        );

    \I__2736\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29510\
        );

    \I__2735\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29510\
        );

    \I__2734\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29510\
        );

    \I__2733\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29510\
        );

    \I__2732\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29510\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__29533\,
            I => \N__29507\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \N__29503\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__29531\,
            I => \N__29499\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__29528\,
            I => \N__29494\
        );

    \I__2727\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29491\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__29510\,
            I => \N__29488\
        );

    \I__2725\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29473\
        );

    \I__2724\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29473\
        );

    \I__2723\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29473\
        );

    \I__2722\ : InMux
    port map (
            O => \N__29502\,
            I => \N__29473\
        );

    \I__2721\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29473\
        );

    \I__2720\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29473\
        );

    \I__2719\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29473\
        );

    \I__2718\ : Sp12to4
    port map (
            O => \N__29494\,
            I => \N__29468\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29468\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__29488\,
            I => \N__29465\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__29473\,
            I => \N__29462\
        );

    \I__2714\ : Span12Mux_s8_h
    port map (
            O => \N__29468\,
            I => \N__29459\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__29465\,
            I => \N__29454\
        );

    \I__2712\ : Span4Mux_h
    port map (
            O => \N__29462\,
            I => \N__29454\
        );

    \I__2711\ : Odrv12
    port map (
            O => \N__29459\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__29454\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840\
        );

    \I__2709\ : InMux
    port map (
            O => \N__29449\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__29446\,
            I => \N__29443\
        );

    \I__2707\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29436\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__29442\,
            I => \N__29433\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__29441\,
            I => \N__29430\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__29440\,
            I => \N__29427\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__29439\,
            I => \N__29423\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__29436\,
            I => \N__29418\
        );

    \I__2701\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29415\
        );

    \I__2700\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29402\
        );

    \I__2699\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29402\
        );

    \I__2698\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29402\
        );

    \I__2697\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29402\
        );

    \I__2696\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29402\
        );

    \I__2695\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29402\
        );

    \I__2694\ : Span4Mux_v
    port map (
            O => \N__29418\,
            I => \N__29399\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__29415\,
            I => \N__29394\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__29402\,
            I => \N__29394\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29391\
        );

    \I__2690\ : Span4Mux_h
    port map (
            O => \N__29394\,
            I => \N__29388\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__29391\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__29388\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843\
        );

    \I__2687\ : InMux
    port map (
            O => \N__29383\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470\
        );

    \I__2686\ : InMux
    port map (
            O => \N__29380\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15471\
        );

    \I__2685\ : InMux
    port map (
            O => \N__29377\,
            I => \foc.u_Park_Transform.n16944\
        );

    \I__2684\ : InMux
    port map (
            O => \N__29374\,
            I => \foc.u_Park_Transform.n16945\
        );

    \I__2683\ : InMux
    port map (
            O => \N__29371\,
            I => \foc.u_Park_Transform.n16946\
        );

    \I__2682\ : InMux
    port map (
            O => \N__29368\,
            I => \foc.u_Park_Transform.n775\
        );

    \I__2681\ : InMux
    port map (
            O => \N__29365\,
            I => \bfn_9_19_0_\
        );

    \I__2680\ : InMux
    port map (
            O => \N__29362\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460\
        );

    \I__2679\ : InMux
    port map (
            O => \N__29359\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461\
        );

    \I__2678\ : InMux
    port map (
            O => \N__29356\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462\
        );

    \I__2677\ : InMux
    port map (
            O => \N__29353\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463\
        );

    \I__2676\ : InMux
    port map (
            O => \N__29350\,
            I => \foc.u_Park_Transform.n16935\
        );

    \I__2675\ : InMux
    port map (
            O => \N__29347\,
            I => \foc.u_Park_Transform.n16936\
        );

    \I__2674\ : InMux
    port map (
            O => \N__29344\,
            I => \foc.u_Park_Transform.n16937\
        );

    \I__2673\ : InMux
    port map (
            O => \N__29341\,
            I => \foc.u_Park_Transform.n16938\
        );

    \I__2672\ : InMux
    port map (
            O => \N__29338\,
            I => \foc.u_Park_Transform.n16939\
        );

    \I__2671\ : InMux
    port map (
            O => \N__29335\,
            I => \foc.u_Park_Transform.n16940\
        );

    \I__2670\ : InMux
    port map (
            O => \N__29332\,
            I => \foc.u_Park_Transform.n16941\
        );

    \I__2669\ : InMux
    port map (
            O => \N__29329\,
            I => \bfn_9_16_0_\
        );

    \I__2668\ : InMux
    port map (
            O => \N__29326\,
            I => \foc.u_Park_Transform.n16943\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__29323\,
            I => \N__29320\
        );

    \I__2666\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29317\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__29317\,
            I => \N__29314\
        );

    \I__2664\ : Odrv12
    port map (
            O => \N__29314\,
            I => \foc.u_Park_Transform.n424_adj_2052\
        );

    \I__2663\ : InMux
    port map (
            O => \N__29311\,
            I => \bfn_9_12_0_\
        );

    \I__2662\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29305\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__29305\,
            I => \N__29302\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__29302\,
            I => \foc.u_Park_Transform.n473_adj_2050\
        );

    \I__2659\ : InMux
    port map (
            O => \N__29299\,
            I => \foc.u_Park_Transform.n17126\
        );

    \I__2658\ : InMux
    port map (
            O => \N__29296\,
            I => \foc.u_Park_Transform.n17127\
        );

    \I__2657\ : InMux
    port map (
            O => \N__29293\,
            I => \foc.u_Park_Transform.n17128\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__29290\,
            I => \N__29285\
        );

    \I__2655\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29282\
        );

    \I__2654\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29277\
        );

    \I__2653\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29277\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__29282\,
            I => \N__29272\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__29277\,
            I => \N__29272\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__29272\,
            I => \foc.u_Park_Transform.n522_adj_2046\
        );

    \I__2649\ : InMux
    port map (
            O => \N__29269\,
            I => \foc.u_Park_Transform.n17129\
        );

    \I__2648\ : InMux
    port map (
            O => \N__29266\,
            I => \foc.u_Park_Transform.n775_adj_2047\
        );

    \I__2647\ : InMux
    port map (
            O => \N__29263\,
            I => \foc.u_Park_Transform.n779_adj_2070\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__29260\,
            I => \N__29257\
        );

    \I__2645\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29251\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__29251\,
            I => \foc.u_Park_Transform.n81\
        );

    \I__2642\ : InMux
    port map (
            O => \N__29248\,
            I => \foc.u_Park_Transform.n17118\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__29245\,
            I => \N__29242\
        );

    \I__2640\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29239\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__29239\,
            I => \N__29236\
        );

    \I__2638\ : Odrv12
    port map (
            O => \N__29236\,
            I => \foc.u_Park_Transform.n130\
        );

    \I__2637\ : InMux
    port map (
            O => \N__29233\,
            I => \foc.u_Park_Transform.n17119\
        );

    \I__2636\ : InMux
    port map (
            O => \N__29230\,
            I => \N__29227\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29224\
        );

    \I__2634\ : Odrv12
    port map (
            O => \N__29224\,
            I => \foc.u_Park_Transform.n179\
        );

    \I__2633\ : InMux
    port map (
            O => \N__29221\,
            I => \foc.u_Park_Transform.n17120\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__29218\,
            I => \N__29215\
        );

    \I__2631\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29212\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__29212\,
            I => \N__29209\
        );

    \I__2629\ : Odrv12
    port map (
            O => \N__29209\,
            I => \foc.u_Park_Transform.n228_adj_2063\
        );

    \I__2628\ : InMux
    port map (
            O => \N__29206\,
            I => \foc.u_Park_Transform.n17121\
        );

    \I__2627\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29200\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29197\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__29197\,
            I => \foc.u_Park_Transform.n277_adj_2060\
        );

    \I__2624\ : InMux
    port map (
            O => \N__29194\,
            I => \foc.u_Park_Transform.n17122\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__29191\,
            I => \N__29188\
        );

    \I__2622\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29185\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29182\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__29182\,
            I => \foc.u_Park_Transform.n326_adj_2056\
        );

    \I__2619\ : InMux
    port map (
            O => \N__29179\,
            I => \foc.u_Park_Transform.n17123\
        );

    \I__2618\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29173\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__29173\,
            I => \N__29170\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__29170\,
            I => \foc.u_Park_Transform.n375_adj_2055\
        );

    \I__2615\ : InMux
    port map (
            O => \N__29167\,
            I => \foc.u_Park_Transform.n17124\
        );

    \I__2614\ : InMux
    port map (
            O => \N__29164\,
            I => \foc.u_Park_Transform.n17108\
        );

    \I__2613\ : InMux
    port map (
            O => \N__29161\,
            I => \foc.u_Park_Transform.n17109\
        );

    \I__2612\ : InMux
    port map (
            O => \N__29158\,
            I => \foc.u_Park_Transform.n17110\
        );

    \I__2611\ : InMux
    port map (
            O => \N__29155\,
            I => \foc.u_Park_Transform.n17111\
        );

    \I__2610\ : InMux
    port map (
            O => \N__29152\,
            I => \foc.u_Park_Transform.n17112\
        );

    \I__2609\ : InMux
    port map (
            O => \N__29149\,
            I => \foc.u_Park_Transform.n17113\
        );

    \I__2608\ : InMux
    port map (
            O => \N__29146\,
            I => \bfn_9_10_0_\
        );

    \I__2607\ : InMux
    port map (
            O => \N__29143\,
            I => \foc.u_Park_Transform.n17115\
        );

    \I__2606\ : InMux
    port map (
            O => \N__29140\,
            I => \foc.u_Park_Transform.n17116\
        );

    \I__2605\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29134\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__29134\,
            I => \N__29131\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__29131\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2744\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__29128\,
            I => \N__29125\
        );

    \I__2601\ : InMux
    port map (
            O => \N__29125\,
            I => \N__29122\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__29122\,
            I => \N__29119\
        );

    \I__2599\ : Odrv12
    port map (
            O => \N__29119\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2841\
        );

    \I__2598\ : InMux
    port map (
            O => \N__29116\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__29113\,
            I => \N__29110\
        );

    \I__2596\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29107\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__29107\,
            I => \N__29104\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__29104\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2844\
        );

    \I__2593\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29098\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29095\
        );

    \I__2591\ : Odrv12
    port map (
            O => \N__29095\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2941\
        );

    \I__2590\ : InMux
    port map (
            O => \N__29092\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466\
        );

    \I__2589\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29086\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__29083\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2944\
        );

    \I__2586\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29077\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__29077\,
            I => \N__29074\
        );

    \I__2584\ : Odrv12
    port map (
            O => \N__29074\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3041\
        );

    \I__2583\ : InMux
    port map (
            O => \N__29071\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467\
        );

    \I__2582\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29065\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__29062\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3044\
        );

    \I__2579\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29056\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__29056\,
            I => \N__29053\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__29053\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3141\
        );

    \I__2576\ : InMux
    port map (
            O => \N__29050\,
            I => \bfn_7_26_0_\
        );

    \I__2575\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29044\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__29044\,
            I => \N__29041\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__29041\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3144\
        );

    \I__2572\ : InMux
    port map (
            O => \N__29038\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469\
        );

    \I__2571\ : InMux
    port map (
            O => \N__29035\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256\
        );

    \I__2570\ : InMux
    port map (
            O => \N__29032\,
            I => \foc.u_Park_Transform.n17107\
        );

    \I__2569\ : InMux
    port map (
            O => \N__29029\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477\
        );

    \I__2568\ : InMux
    port map (
            O => \N__29026\,
            I => \bfn_7_24_0_\
        );

    \I__2567\ : InMux
    port map (
            O => \N__29023\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479\
        );

    \I__2566\ : InMux
    port map (
            O => \N__29020\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260\
        );

    \I__2565\ : InMux
    port map (
            O => \N__29017\,
            I => \N__29014\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__29011\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__29011\,
            I => \N__29008\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__29008\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2341\
        );

    \I__2561\ : InMux
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__28999\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2344\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__2557\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__28984\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2441\
        );

    \I__2553\ : InMux
    port map (
            O => \N__28981\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__28978\,
            I => \N__28975\
        );

    \I__2551\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28969\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__28969\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2444\
        );

    \I__2548\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28963\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28960\
        );

    \I__2546\ : Sp12to4
    port map (
            O => \N__28960\,
            I => \N__28957\
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__28957\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2541\
        );

    \I__2544\ : InMux
    port map (
            O => \N__28954\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462\
        );

    \I__2543\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28948\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28945\
        );

    \I__2541\ : Odrv12
    port map (
            O => \N__28945\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2544\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__28942\,
            I => \N__28939\
        );

    \I__2539\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28936\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28933\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__28933\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2641\
        );

    \I__2536\ : InMux
    port map (
            O => \N__28930\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__28927\,
            I => \N__28924\
        );

    \I__2534\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28921\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__28921\,
            I => \N__28918\
        );

    \I__2532\ : Odrv12
    port map (
            O => \N__28918\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2644\
        );

    \I__2531\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28912\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__28912\,
            I => \N__28909\
        );

    \I__2529\ : Odrv12
    port map (
            O => \N__28909\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2741\
        );

    \I__2528\ : InMux
    port map (
            O => \N__28906\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464\
        );

    \I__2527\ : InMux
    port map (
            O => \N__28903\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459\
        );

    \I__2526\ : InMux
    port map (
            O => \N__28900\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252\
        );

    \I__2525\ : InMux
    port map (
            O => \N__28897\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471\
        );

    \I__2524\ : InMux
    port map (
            O => \N__28894\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472\
        );

    \I__2523\ : InMux
    port map (
            O => \N__28891\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473\
        );

    \I__2522\ : InMux
    port map (
            O => \N__28888\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474\
        );

    \I__2521\ : InMux
    port map (
            O => \N__28885\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475\
        );

    \I__2520\ : InMux
    port map (
            O => \N__28882\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__28879\,
            I => \N__28876\
        );

    \I__2518\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28870\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__28870\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2438\
        );

    \I__2515\ : InMux
    port map (
            O => \N__28867\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451\
        );

    \I__2514\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28861\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__28858\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2538\
        );

    \I__2511\ : InMux
    port map (
            O => \N__28855\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__28852\,
            I => \N__28849\
        );

    \I__2509\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__28846\,
            I => \N__28843\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__28843\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2638\
        );

    \I__2506\ : InMux
    port map (
            O => \N__28840\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453\
        );

    \I__2505\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28834\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28831\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__28831\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2738\
        );

    \I__2502\ : InMux
    port map (
            O => \N__28828\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__28825\,
            I => \N__28822\
        );

    \I__2500\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28816\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__28816\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2838\
        );

    \I__2497\ : InMux
    port map (
            O => \N__28813\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455\
        );

    \I__2496\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28807\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__28807\,
            I => \N__28804\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__28804\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2938\
        );

    \I__2493\ : InMux
    port map (
            O => \N__28801\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456\
        );

    \I__2492\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28795\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__28795\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3038\
        );

    \I__2490\ : InMux
    port map (
            O => \N__28792\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457\
        );

    \I__2489\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28786\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28783\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__28783\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3138\
        );

    \I__2486\ : InMux
    port map (
            O => \N__28780\,
            I => \bfn_7_22_0_\
        );

    \I__2485\ : InMux
    port map (
            O => \N__28777\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444\
        );

    \I__2484\ : InMux
    port map (
            O => \N__28774\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445\
        );

    \I__2483\ : InMux
    port map (
            O => \N__28771\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446\
        );

    \I__2482\ : InMux
    port map (
            O => \N__28768\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447\
        );

    \I__2481\ : InMux
    port map (
            O => \N__28765\,
            I => \bfn_7_20_0_\
        );

    \I__2480\ : InMux
    port map (
            O => \N__28762\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449\
        );

    \I__2479\ : InMux
    port map (
            O => \N__28759\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__28756\,
            I => \N__28752\
        );

    \I__2477\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28741\
        );

    \I__2476\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28741\
        );

    \I__2475\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28741\
        );

    \I__2474\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28741\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__28741\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8490\
        );

    \I__2472\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28735\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__28735\,
            I => \N__28732\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__28732\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2338\
        );

    \I__2469\ : InMux
    port map (
            O => \N__28729\,
            I => \N__28726\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__28726\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8175\
        );

    \I__2467\ : InMux
    port map (
            O => \N__28723\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346\
        );

    \I__2466\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28717\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__28717\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8174\
        );

    \I__2464\ : InMux
    port map (
            O => \N__28714\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347\
        );

    \I__2463\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28708\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__28708\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8173\
        );

    \I__2461\ : InMux
    port map (
            O => \N__28705\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348\
        );

    \I__2460\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28699\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__28699\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8172\
        );

    \I__2458\ : InMux
    port map (
            O => \N__28696\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17349\
        );

    \I__2457\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__28690\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8177\
        );

    \I__2455\ : InMux
    port map (
            O => \N__28687\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441\
        );

    \I__2454\ : InMux
    port map (
            O => \N__28684\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442\
        );

    \I__2453\ : InMux
    port map (
            O => \N__28681\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443\
        );

    \I__2452\ : InMux
    port map (
            O => \N__28678\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332\
        );

    \I__2451\ : InMux
    port map (
            O => \N__28675\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333\
        );

    \I__2450\ : InMux
    port map (
            O => \N__28672\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334\
        );

    \I__2449\ : InMux
    port map (
            O => \N__28669\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335\
        );

    \I__2448\ : InMux
    port map (
            O => \N__28666\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17336\
        );

    \I__2447\ : InMux
    port map (
            O => \N__28663\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344\
        );

    \I__2446\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28657\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__28657\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8176\
        );

    \I__2444\ : InMux
    port map (
            O => \N__28654\,
            I => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345\
        );

    \I__2443\ : IoInMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__28648\,
            I => \N__28645\
        );

    \I__2441\ : Span12Mux_s8_h
    port map (
            O => \N__28645\,
            I => \N__28642\
        );

    \I__2440\ : Span12Mux_v
    port map (
            O => \N__28642\,
            I => \N__28639\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__28639\,
            I => pin3_clk_16mhz_pad_gb_input
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17365\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17090\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16907\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_19_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_21_0_\
        );

    \IN_MUX_bfv_19_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18151\,
            carryinitout => \bfn_19_22_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18159\,
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17964\,
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17972\,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15727\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15735\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15743\,
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_18_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_26_0_\
        );

    \IN_MUX_bfv_18_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18361\,
            carryinitout => \bfn_18_27_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_19_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17718\,
            carryinitout => \bfn_19_18_0_\
        );

    \IN_MUX_bfv_19_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17726\,
            carryinitout => \bfn_19_19_0_\
        );

    \IN_MUX_bfv_20_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_14_0_\
        );

    \IN_MUX_bfv_20_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17512\,
            carryinitout => \bfn_20_15_0_\
        );

    \IN_MUX_bfv_20_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17520\,
            carryinitout => \bfn_20_16_0_\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15782\,
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15790\,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15798\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_19_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_9_0_\
        );

    \IN_MUX_bfv_19_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17934\,
            carryinitout => \bfn_19_10_0_\
        );

    \IN_MUX_bfv_6_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17419\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17410\,
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17401\,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17392\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17383\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17374\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15951\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17497\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15467\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_10_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17357\,
            carryinitout => \bfn_10_26_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17488\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_7_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_23_0_\
        );

    \IN_MUX_bfv_7_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17478\,
            carryinitout => \bfn_7_24_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17468\,
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17458\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17448\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17438\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17428\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n15755\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n15763\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n15771\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17284\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17292\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17300\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16922\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16931\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16942\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16955\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16970\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n16985\,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17000\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17015\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17030\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17045\,
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17060\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17075\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17105\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17114\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17125\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17138\,
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17153\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17168\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17183\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17198\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17213\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17228\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17243\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_Park_Transform.n17258\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17734\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17863\,
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_12_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17663\,
            carryinitout => \bfn_12_23_0_\
        );

    \IN_MUX_bfv_12_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_24_0_\
        );

    \IN_MUX_bfv_12_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18114\,
            carryinitout => \bfn_12_25_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18099\,
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18084\,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18069\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18054\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18039\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_16_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18024\,
            carryinitout => \bfn_16_26_0_\
        );

    \IN_MUX_bfv_16_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_27_0_\
        );

    \IN_MUX_bfv_16_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18009\,
            carryinitout => \bfn_16_28_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17994\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_21_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_23_0_\
        );

    \IN_MUX_bfv_21_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15920\,
            carryinitout => \bfn_21_24_0_\
        );

    \IN_MUX_bfv_21_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15928\,
            carryinitout => \bfn_21_25_0_\
        );

    \IN_MUX_bfv_21_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15936\,
            carryinitout => \bfn_21_26_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15890\,
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_18_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15898\,
            carryinitout => \bfn_18_24_0_\
        );

    \IN_MUX_bfv_18_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15906\,
            carryinitout => \bfn_18_25_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_25_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18376\,
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_19_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_26_0_\
        );

    \IN_MUX_bfv_19_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18346\,
            carryinitout => \bfn_19_27_0_\
        );

    \IN_MUX_bfv_19_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_28_0_\
        );

    \IN_MUX_bfv_19_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18331\,
            carryinitout => \bfn_19_29_0_\
        );

    \IN_MUX_bfv_20_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_28_0_\
        );

    \IN_MUX_bfv_20_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18316\,
            carryinitout => \bfn_20_29_0_\
        );

    \IN_MUX_bfv_21_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_28_0_\
        );

    \IN_MUX_bfv_21_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18301\,
            carryinitout => \bfn_21_29_0_\
        );

    \IN_MUX_bfv_22_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_28_0_\
        );

    \IN_MUX_bfv_22_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18286\,
            carryinitout => \bfn_22_29_0_\
        );

    \IN_MUX_bfv_23_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_27_0_\
        );

    \IN_MUX_bfv_23_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18271\,
            carryinitout => \bfn_23_28_0_\
        );

    \IN_MUX_bfv_23_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_25_0_\
        );

    \IN_MUX_bfv_23_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18256\,
            carryinitout => \bfn_23_26_0_\
        );

    \IN_MUX_bfv_22_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_25_0_\
        );

    \IN_MUX_bfv_22_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18241\,
            carryinitout => \bfn_22_26_0_\
        );

    \IN_MUX_bfv_20_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_25_0_\
        );

    \IN_MUX_bfv_20_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18226\,
            carryinitout => \bfn_20_26_0_\
        );

    \IN_MUX_bfv_20_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_23_0_\
        );

    \IN_MUX_bfv_20_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18211\,
            carryinitout => \bfn_20_24_0_\
        );

    \IN_MUX_bfv_19_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_24_0_\
        );

    \IN_MUX_bfv_19_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18196\,
            carryinitout => \bfn_19_25_0_\
        );

    \IN_MUX_bfv_21_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_21_0_\
        );

    \IN_MUX_bfv_21_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18181\,
            carryinitout => \bfn_21_22_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_5_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18142\,
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_18_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_5_0_\
        );

    \IN_MUX_bfv_18_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17273\,
            carryinitout => \bfn_18_6_0_\
        );

    \IN_MUX_bfv_20_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_5_0_\
        );

    \IN_MUX_bfv_20_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18129\,
            carryinitout => \bfn_20_6_0_\
        );

    \IN_MUX_bfv_19_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_5_0_\
        );

    \IN_MUX_bfv_19_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17648\,
            carryinitout => \bfn_19_6_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17633\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_20_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_7_0_\
        );

    \IN_MUX_bfv_20_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17618\,
            carryinitout => \bfn_20_8_0_\
        );

    \IN_MUX_bfv_21_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_7_0_\
        );

    \IN_MUX_bfv_21_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17603\,
            carryinitout => \bfn_21_8_0_\
        );

    \IN_MUX_bfv_20_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_9_0_\
        );

    \IN_MUX_bfv_20_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17588\,
            carryinitout => \bfn_20_10_0_\
        );

    \IN_MUX_bfv_21_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_9_0_\
        );

    \IN_MUX_bfv_21_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17573\,
            carryinitout => \bfn_21_10_0_\
        );

    \IN_MUX_bfv_21_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_11_0_\
        );

    \IN_MUX_bfv_21_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17558\,
            carryinitout => \bfn_21_12_0_\
        );

    \IN_MUX_bfv_22_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_11_0_\
        );

    \IN_MUX_bfv_22_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17543\,
            carryinitout => \bfn_22_12_0_\
        );

    \IN_MUX_bfv_23_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_11_0_\
        );

    \IN_MUX_bfv_23_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17528\,
            carryinitout => \bfn_23_12_0_\
        );

    \IN_MUX_bfv_22_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_19_0_\
        );

    \IN_MUX_bfv_22_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15980\,
            carryinitout => \bfn_22_20_0_\
        );

    \IN_MUX_bfv_22_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15988\,
            carryinitout => \bfn_22_21_0_\
        );

    \IN_MUX_bfv_22_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15996\,
            carryinitout => \bfn_22_22_0_\
        );

    \IN_MUX_bfv_24_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_16_0_\
        );

    \IN_MUX_bfv_24_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_24_17_0_\
        );

    \IN_MUX_bfv_24_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15580_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_24_18_0_\
        );

    \IN_MUX_bfv_24_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15588\,
            carryinitout => \bfn_24_19_0_\
        );

    \IN_MUX_bfv_24_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15596\,
            carryinitout => \bfn_24_20_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17949\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_19_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_11_0_\
        );

    \IN_MUX_bfv_19_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17919\,
            carryinitout => \bfn_19_12_0_\
        );

    \IN_MUX_bfv_20_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_11_0_\
        );

    \IN_MUX_bfv_20_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17904\,
            carryinitout => \bfn_20_12_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17889\,
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17874\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17848\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17833\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_19_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_13_0_\
        );

    \IN_MUX_bfv_19_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17818\,
            carryinitout => \bfn_19_14_0_\
        );

    \IN_MUX_bfv_19_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_15_0_\
        );

    \IN_MUX_bfv_19_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17803\,
            carryinitout => \bfn_19_16_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17788\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17773\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17758\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_21_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_17_0_\
        );

    \IN_MUX_bfv_21_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17743\,
            carryinitout => \bfn_21_18_0_\
        );

    \pin3_clk_16mhz_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__28651\,
            GLOBALBUFFEROUTPUT => \pin3_clk_16mhz_N\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_2_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31562\,
            in2 => \N__32765\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7897\,
            ltout => OPEN,
            carryin => \bfn_6_20_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_3_lut_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28750\,
            in2 => \_gnd_net_\,
            in3 => \N__28678\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8176\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_4_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31563\,
            in2 => \N__32766\,
            in3 => \N__28675\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8175\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_5_lut_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28751\,
            in2 => \N__31573\,
            in3 => \N__28672\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8174\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_6_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31567\,
            in2 => \N__28756\,
            in3 => \N__28669\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8173\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17336\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_7_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31568\,
            in1 => \N__28755\,
            in2 => \_gnd_net_\,
            in3 => \N__28666\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_2_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31547\,
            in2 => \N__32799\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7554\,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28693\,
            in2 => \_gnd_net_\,
            in3 => \N__28663\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7896\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_4_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28660\,
            in2 => \N__31571\,
            in3 => \N__28654\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7895\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_5_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28729\,
            in2 => \N__31569\,
            in3 => \N__28723\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7894\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_6_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28720\,
            in2 => \N__31572\,
            in3 => \N__28714\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7893\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_7_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28711\,
            in2 => \N__31570\,
            in3 => \N__28705\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7892\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17349\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_8_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28702\,
            in1 => \N__31554\,
            in2 => \_gnd_net_\,
            in3 => \N__28696\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7891\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_2_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31561\,
            in2 => \_gnd_net_\,
            in3 => \N__32783\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_2_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29596\,
            in2 => \N__32796\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2335\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_3_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28738\,
            in2 => \_gnd_net_\,
            in3 => \N__28687\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2435\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_4_lut_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29597\,
            in2 => \N__28879\,
            in3 => \N__28684\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2535\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_5_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28864\,
            in2 => \N__29609\,
            in3 => \N__28681\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2635\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_6_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29601\,
            in2 => \N__28852\,
            in3 => \N__28777\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2735\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_7_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28837\,
            in2 => \N__29610\,
            in3 => \N__28774\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2835\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_8_lut_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29605\,
            in2 => \N__28825\,
            in3 => \N__28771\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2935\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_9_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28810\,
            in2 => \N__29611\,
            in3 => \N__28768\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3035\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17448\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_10_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28798\,
            in2 => \N__29595\,
            in3 => \N__28765\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3135\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_11_lut_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28789\,
            in2 => \_gnd_net_\,
            in3 => \N__28762\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3247\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_LUT4_0_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28759\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.i13555_2_lut_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32728\,
            in2 => \_gnd_net_\,
            in3 => \N__44911\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_2_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29497\,
            in2 => \N__32797\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2338\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_3_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29017\,
            in2 => \_gnd_net_\,
            in3 => \N__28867\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2438\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_4_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29498\,
            in2 => \N__28996\,
            in3 => \N__28855\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2538\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_5_lut_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28966\,
            in2 => \N__29531\,
            in3 => \N__28840\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2638\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_6_lut_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29502\,
            in2 => \N__28942\,
            in3 => \N__28828\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2738\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_7_lut_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28915\,
            in2 => \N__29532\,
            in3 => \N__28813\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2838\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_8_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29506\,
            in2 => \N__29128\,
            in3 => \N__28801\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2938\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_9_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29101\,
            in2 => \N__29533\,
            in3 => \N__28792\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3038\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17458\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_10_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29080\,
            in2 => \N__29547\,
            in3 => \N__28780\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3138\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_11_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29059\,
            in2 => \_gnd_net_\,
            in3 => \N__28903\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3251\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_LUT4_0_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28900\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_2_lut_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29421\,
            in2 => \N__32800\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2344\,
            ltout => OPEN,
            carryin => \bfn_7_23_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_3_lut_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30034\,
            in2 => \_gnd_net_\,
            in3 => \N__28897\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2444\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_4_lut_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29422\,
            in2 => \N__30016\,
            in3 => \N__28894\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2544\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_5_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29998\,
            in2 => \N__29439\,
            in3 => \N__28891\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2644\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_6_lut_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29426\,
            in2 => \N__29983\,
            in3 => \N__28888\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2744\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_7_lut_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29965\,
            in2 => \N__29440\,
            in3 => \N__28885\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2844\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_8_lut_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29950\,
            in2 => \N__29442\,
            in3 => \N__28882\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2944\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_9_lut_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29935\,
            in2 => \N__29441\,
            in3 => \N__29029\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3044\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17478\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_10_lut_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30094\,
            in2 => \N__29446\,
            in3 => \N__29026\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3144\,
            ltout => OPEN,
            carryin => \bfn_7_24_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_11_lut_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30082\,
            in2 => \_gnd_net_\,
            in3 => \N__29023\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3259\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_LUT4_0_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29020\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_2_lut_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29534\,
            in2 => \N__32806\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2341\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_3_lut_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29005\,
            in2 => \_gnd_net_\,
            in3 => \N__28981\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2441\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_4_lut_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29535\,
            in2 => \N__28978\,
            in3 => \N__28954\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2541\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_5_lut_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28951\,
            in2 => \N__29551\,
            in3 => \N__28930\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2641\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_6_lut_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29539\,
            in2 => \N__28927\,
            in3 => \N__28906\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2741\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_7_lut_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29137\,
            in2 => \N__29552\,
            in3 => \N__29116\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2841\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_8_lut_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29543\,
            in2 => \N__29113\,
            in3 => \N__29092\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2941\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_9_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29089\,
            in2 => \N__29553\,
            in3 => \N__29071\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3041\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17468\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_10_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29068\,
            in2 => \N__29560\,
            in3 => \N__29050\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3141\,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_11_lut_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29047\,
            in2 => \_gnd_net_\,
            in3 => \N__29038\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3255\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_LUT4_0_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29035\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_2_lut_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31747\,
            in2 => \N__30850\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n81\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \foc.u_Park_Transform.n17107\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_3_lut_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30844\,
            in2 => \N__31375\,
            in3 => \N__29032\,
            lcout => \foc.u_Park_Transform.n130\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17107\,
            carryout => \foc.u_Park_Transform.n17108\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_4_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30796\,
            in2 => \N__31363\,
            in3 => \N__29164\,
            lcout => \foc.u_Park_Transform.n179\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17108\,
            carryout => \foc.u_Park_Transform.n17109\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_5_lut_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31897\,
            in2 => \N__30837\,
            in3 => \N__29161\,
            lcout => \foc.u_Park_Transform.n228_adj_2063\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17109\,
            carryout => \foc.u_Park_Transform.n17110\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_6_lut_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30800\,
            in2 => \N__31885\,
            in3 => \N__29158\,
            lcout => \foc.u_Park_Transform.n277_adj_2060\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17110\,
            carryout => \foc.u_Park_Transform.n17111\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_7_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31870\,
            in2 => \N__30838\,
            in3 => \N__29155\,
            lcout => \foc.u_Park_Transform.n326_adj_2056\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17111\,
            carryout => \foc.u_Park_Transform.n17112\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_8_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30804\,
            in2 => \N__31855\,
            in3 => \N__29152\,
            lcout => \foc.u_Park_Transform.n375_adj_2055\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17112\,
            carryout => \foc.u_Park_Transform.n17113\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_9_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31837\,
            in2 => \N__30839\,
            in3 => \N__29149\,
            lcout => \foc.u_Park_Transform.n424_adj_2052\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17113\,
            carryout => \foc.u_Park_Transform.n17114\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_10_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30808\,
            in2 => \N__31824\,
            in3 => \N__29146\,
            lcout => \foc.u_Park_Transform.n473_adj_2050\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \foc.u_Park_Transform.n17115\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_11_lut_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31820\,
            in2 => \N__30840\,
            in3 => \N__29143\,
            lcout => \foc.u_Park_Transform.n522_adj_2046\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17115\,
            carryout => \foc.u_Park_Transform.n17116\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_12_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30687\,
            in2 => \N__31825\,
            in3 => \N__29140\,
            lcout => \foc.u_Park_Transform.n778_adj_2068\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17116\,
            carryout => \foc.u_Park_Transform.n779_adj_2070\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n779_adj_2070_THRU_LUT4_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29263\,
            lcout => \foc.u_Park_Transform.n779_adj_2070_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_2_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30764\,
            in2 => \N__32369\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n78\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \foc.u_Park_Transform.n17118\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_3_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32330\,
            in2 => \N__29260\,
            in3 => \N__29248\,
            lcout => \foc.u_Park_Transform.n127\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17118\,
            carryout => \foc.u_Park_Transform.n17119\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_4_lut_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32331\,
            in2 => \N__29245\,
            in3 => \N__29233\,
            lcout => \foc.u_Park_Transform.n176\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17119\,
            carryout => \foc.u_Park_Transform.n17120\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_5_lut_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29230\,
            in2 => \N__32370\,
            in3 => \N__29221\,
            lcout => \foc.u_Park_Transform.n225\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17120\,
            carryout => \foc.u_Park_Transform.n17121\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_6_lut_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32335\,
            in2 => \N__29218\,
            in3 => \N__29206\,
            lcout => \foc.u_Park_Transform.n274\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17121\,
            carryout => \foc.u_Park_Transform.n17122\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_7_lut_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29203\,
            in2 => \N__32371\,
            in3 => \N__29194\,
            lcout => \foc.u_Park_Transform.n323\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17122\,
            carryout => \foc.u_Park_Transform.n17123\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_8_lut_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32339\,
            in2 => \N__29191\,
            in3 => \N__29179\,
            lcout => \foc.u_Park_Transform.n372\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17123\,
            carryout => \foc.u_Park_Transform.n17124\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_9_lut_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29176\,
            in2 => \N__32372\,
            in3 => \N__29167\,
            lcout => \foc.u_Park_Transform.n421_adj_2039\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17124\,
            carryout => \foc.u_Park_Transform.n17125\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_10_lut_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32319\,
            in2 => \N__29323\,
            in3 => \N__29311\,
            lcout => \foc.u_Park_Transform.n470_adj_2038\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \foc.u_Park_Transform.n17126\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_11_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29308\,
            in2 => \N__32367\,
            in3 => \N__29299\,
            lcout => \foc.u_Park_Transform.n519_adj_2035\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17126\,
            carryout => \foc.u_Park_Transform.n17127\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_12_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32323\,
            in2 => \N__29290\,
            in3 => \N__29296\,
            lcout => \foc.u_Park_Transform.n568_adj_2034\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17127\,
            carryout => \foc.u_Park_Transform.n17128\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_13_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29288\,
            in2 => \N__32368\,
            in3 => \N__29293\,
            lcout => \foc.u_Park_Transform.n617_adj_2031\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17128\,
            carryout => \foc.u_Park_Transform.n17129\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_14_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29289\,
            in2 => \N__30447\,
            in3 => \N__29269\,
            lcout => \foc.u_Park_Transform.n774_adj_2045\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17129\,
            carryout => \foc.u_Park_Transform.n775_adj_2047\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n775_adj_2047_THRU_LUT4_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29266\,
            lcout => \foc.u_Park_Transform.n775_adj_2047_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i22_2_lut_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__32157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i528_2_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32158\,
            lcout => \foc.u_Park_Transform.n777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_2_lut_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30734\,
            in2 => \N__32384\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n78_adj_2145\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \foc.u_Park_Transform.n16935\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_3_lut_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32363\,
            in2 => \N__30601\,
            in3 => \N__29350\,
            lcout => \foc.u_Park_Transform.n127_adj_2119\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16935\,
            carryout => \foc.u_Park_Transform.n16936\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_4_lut_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32381\,
            in2 => \N__30577\,
            in3 => \N__29347\,
            lcout => \foc.u_Park_Transform.n176_adj_2104\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16936\,
            carryout => \foc.u_Park_Transform.n16937\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_5_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32364\,
            in2 => \N__30547\,
            in3 => \N__29344\,
            lcout => \foc.u_Park_Transform.n225_adj_2075\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16937\,
            carryout => \foc.u_Park_Transform.n16938\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_6_lut_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32382\,
            in2 => \N__30523\,
            in3 => \N__29341\,
            lcout => \foc.u_Park_Transform.n274_adj_2058\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16938\,
            carryout => \foc.u_Park_Transform.n16939\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_7_lut_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32365\,
            in2 => \N__30955\,
            in3 => \N__29338\,
            lcout => \foc.u_Park_Transform.n323_adj_2057\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16939\,
            carryout => \foc.u_Park_Transform.n16940\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_8_lut_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32383\,
            in2 => \N__30928\,
            in3 => \N__29335\,
            lcout => \foc.u_Park_Transform.n372_adj_2042\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16940\,
            carryout => \foc.u_Park_Transform.n16941\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_9_lut_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32366\,
            in2 => \N__30901\,
            in3 => \N__29332\,
            lcout => \foc.u_Park_Transform.n421\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16941\,
            carryout => \foc.u_Park_Transform.n16942\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_10_lut_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30874\,
            in2 => \N__32385\,
            in3 => \N__29329\,
            lcout => \foc.u_Park_Transform.n470\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \foc.u_Park_Transform.n16943\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_11_lut_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32376\,
            in2 => \N__30865\,
            in3 => \N__29326\,
            lcout => \foc.u_Park_Transform.n519\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16943\,
            carryout => \foc.u_Park_Transform.n16944\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_12_lut_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30707\,
            in2 => \N__32386\,
            in3 => \N__29377\,
            lcout => \foc.u_Park_Transform.n568\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16944\,
            carryout => \foc.u_Park_Transform.n16945\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_13_lut_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32380\,
            in2 => \N__30712\,
            in3 => \N__29374\,
            lcout => \foc.u_Park_Transform.n617\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16945\,
            carryout => \foc.u_Park_Transform.n16946\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_570_14_lut_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30711\,
            in2 => \N__30451\,
            in3 => \N__29371\,
            lcout => \foc.u_Park_Transform.n774\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16946\,
            carryout => \foc.u_Park_Transform.n775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n775_THRU_LUT4_0_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29368\,
            lcout => \foc.u_Park_Transform.n775_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44946\,
            in2 => \_gnd_net_\,
            in3 => \N__29365\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2807\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44949\,
            in2 => \_gnd_net_\,
            in3 => \N__29362\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68428\,
            in2 => \_gnd_net_\,
            in3 => \N__29359\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44950\,
            in2 => \_gnd_net_\,
            in3 => \N__29356\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44947\,
            in2 => \_gnd_net_\,
            in3 => \N__29353\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44951\,
            in2 => \_gnd_net_\,
            in3 => \N__29623\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44948\,
            in2 => \_gnd_net_\,
            in3 => \N__29620\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2825\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44952\,
            in2 => \_gnd_net_\,
            in3 => \N__29617\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2828\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15467\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44954\,
            in2 => \_gnd_net_\,
            in3 => \N__29614\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44953\,
            in2 => \_gnd_net_\,
            in3 => \N__29563\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2834\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44955\,
            in2 => \_gnd_net_\,
            in3 => \N__29449\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68436\,
            in2 => \_gnd_net_\,
            in3 => \N__29383\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15471\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__68437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29380\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_2_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32693\,
            in2 => \N__29672\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2332\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_3_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29803\,
            in2 => \_gnd_net_\,
            in3 => \N__29791\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2432\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_4_lut_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29788\,
            in2 => \N__29673\,
            in3 => \N__29776\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2532\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_5_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29658\,
            in2 => \N__29773\,
            in3 => \N__29758\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2632\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_6_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29755\,
            in2 => \N__29674\,
            in3 => \N__29743\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2732\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_7_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29662\,
            in2 => \N__29740\,
            in3 => \N__29725\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2832\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_8_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29722\,
            in2 => \N__29675\,
            in3 => \N__29710\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2932\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_9_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29707\,
            in2 => \N__29676\,
            in3 => \N__29695\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3032\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17438\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_10_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29692\,
            in2 => \N__29680\,
            in3 => \N__29626\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3132\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_11_lut_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29920\,
            in2 => \_gnd_net_\,
            in3 => \N__29908\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3243\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_LUT4_0_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29905\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_2_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31500\,
            in2 => \N__32770\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7473\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_3_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29902\,
            in2 => \_gnd_net_\,
            in3 => \N__29890\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7553\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_4_lut_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31501\,
            in2 => \N__29887\,
            in3 => \N__29872\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7552\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_5_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29869\,
            in2 => \N__31518\,
            in3 => \N__29857\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7551\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_6_lut_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31505\,
            in2 => \N__29854\,
            in3 => \N__29839\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7550\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_7_lut_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29836\,
            in2 => \N__31519\,
            in3 => \N__29824\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7549\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_8_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31509\,
            in2 => \N__29821\,
            in3 => \N__29806\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7548\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17343\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_9_lut_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31510\,
            in1 => \N__30049\,
            in2 => \_gnd_net_\,
            in3 => \N__30037\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_2_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32798\,
            in2 => \N__31496\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2347\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_3_lut_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30022\,
            in2 => \_gnd_net_\,
            in3 => \N__30001\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2447\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_4_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31243\,
            in2 => \N__31497\,
            in3 => \N__29986\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2547\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_5_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31464\,
            in2 => \N__31222\,
            in3 => \N__29968\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2647\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_6_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31669\,
            in2 => \N__31498\,
            in3 => \N__29953\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2747\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_7_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31468\,
            in2 => \N__31651\,
            in3 => \N__29938\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2847\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_8_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31630\,
            in2 => \N__31499\,
            in3 => \N__29923\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2947\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_9_lut_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31472\,
            in2 => \N__31612\,
            in3 => \N__30085\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3047\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17488\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_10_lut_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31591\,
            in2 => \N__31495\,
            in3 => \N__30070\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3147\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17489\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_11_lut_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__31381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30067\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_2_lut_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34278\,
            in2 => \N__35893\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n72\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \foc.u_Park_Transform.n17146\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_3_lut_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35870\,
            in2 => \N__30262\,
            in3 => \N__30064\,
            lcout => \foc.u_Park_Transform.n121\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17146\,
            carryout => \foc.u_Park_Transform.n17147\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_4_lut_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35871\,
            in2 => \N__30241\,
            in3 => \N__30061\,
            lcout => \foc.u_Park_Transform.n170\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17147\,
            carryout => \foc.u_Park_Transform.n17148\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_5_lut_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30217\,
            in2 => \N__35894\,
            in3 => \N__30058\,
            lcout => \foc.u_Park_Transform.n219\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17148\,
            carryout => \foc.u_Park_Transform.n17149\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_6_lut_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35875\,
            in2 => \N__30199\,
            in3 => \N__30055\,
            lcout => \foc.u_Park_Transform.n268\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17149\,
            carryout => \foc.u_Park_Transform.n17150\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_7_lut_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30175\,
            in2 => \N__35895\,
            in3 => \N__30052\,
            lcout => \foc.u_Park_Transform.n317\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17150\,
            carryout => \foc.u_Park_Transform.n17151\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_8_lut_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35879\,
            in2 => \N__30157\,
            in3 => \N__30121\,
            lcout => \foc.u_Park_Transform.n366\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17151\,
            carryout => \foc.u_Park_Transform.n17152\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_9_lut_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30133\,
            in2 => \N__35896\,
            in3 => \N__30118\,
            lcout => \foc.u_Park_Transform.n415_adj_2008\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17152\,
            carryout => \foc.u_Park_Transform.n17153\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_10_lut_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30412\,
            in2 => \N__35810\,
            in3 => \N__30115\,
            lcout => \foc.u_Park_Transform.n464_adj_2005\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \foc.u_Park_Transform.n17154\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_11_lut_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35758\,
            in2 => \N__30397\,
            in3 => \N__30112\,
            lcout => \foc.u_Park_Transform.n513_adj_2002\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17154\,
            carryout => \foc.u_Park_Transform.n17155\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_12_lut_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30373\,
            in2 => \N__35811\,
            in3 => \N__30109\,
            lcout => \foc.u_Park_Transform.n562_adj_2000\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17155\,
            carryout => \foc.u_Park_Transform.n17156\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_13_lut_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35762\,
            in2 => \N__30355\,
            in3 => \N__30106\,
            lcout => \foc.u_Park_Transform.n611\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17156\,
            carryout => \foc.u_Park_Transform.n17157\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_14_lut_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30331\,
            in2 => \N__35812\,
            in3 => \N__30103\,
            lcout => \foc.u_Park_Transform.n660\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17157\,
            carryout => \foc.u_Park_Transform.n17158\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_15_lut_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35766\,
            in2 => \N__30319\,
            in3 => \N__30100\,
            lcout => \foc.u_Park_Transform.n709\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17158\,
            carryout => \foc.u_Park_Transform.n17159\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_16_lut_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34500\,
            in2 => \N__30304\,
            in3 => \N__30097\,
            lcout => \foc.u_Park_Transform.n766\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17159\,
            carryout => \foc.u_Park_Transform.n767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n767_THRU_LUT4_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30265\,
            lcout => \foc.u_Park_Transform.n767_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_2_lut_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32318\,
            in2 => \N__34272\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n75\,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \foc.u_Park_Transform.n17131\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_3_lut_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34227\,
            in2 => \N__30250\,
            in3 => \N__30229\,
            lcout => \foc.u_Park_Transform.n124\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17131\,
            carryout => \foc.u_Park_Transform.n17132\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_4_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34228\,
            in2 => \N__30226\,
            in3 => \N__30208\,
            lcout => \foc.u_Park_Transform.n173\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17132\,
            carryout => \foc.u_Park_Transform.n17133\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_5_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30205\,
            in2 => \N__34273\,
            in3 => \N__30187\,
            lcout => \foc.u_Park_Transform.n222\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17133\,
            carryout => \foc.u_Park_Transform.n17134\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_6_lut_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34232\,
            in2 => \N__30184\,
            in3 => \N__30166\,
            lcout => \foc.u_Park_Transform.n271\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17134\,
            carryout => \foc.u_Park_Transform.n17135\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_7_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30163\,
            in2 => \N__34274\,
            in3 => \N__30145\,
            lcout => \foc.u_Park_Transform.n320\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17135\,
            carryout => \foc.u_Park_Transform.n17136\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_8_lut_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34236\,
            in2 => \N__30142\,
            in3 => \N__30124\,
            lcout => \foc.u_Park_Transform.n369\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17136\,
            carryout => \foc.u_Park_Transform.n17137\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_9_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30418\,
            in2 => \N__34275\,
            in3 => \N__30406\,
            lcout => \foc.u_Park_Transform.n418_adj_2024\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17137\,
            carryout => \foc.u_Park_Transform.n17138\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_10_lut_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30403\,
            in2 => \N__34221\,
            in3 => \N__30385\,
            lcout => \foc.u_Park_Transform.n467_adj_2019\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \foc.u_Park_Transform.n17139\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_11_lut_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34165\,
            in2 => \N__30382\,
            in3 => \N__30364\,
            lcout => \foc.u_Park_Transform.n516_adj_2018\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17139\,
            carryout => \foc.u_Park_Transform.n17140\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_12_lut_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30361\,
            in2 => \N__34222\,
            in3 => \N__30343\,
            lcout => \foc.u_Park_Transform.n565\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17140\,
            carryout => \foc.u_Park_Transform.n17141\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_13_lut_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34169\,
            in2 => \N__30340\,
            in3 => \N__30322\,
            lcout => \foc.u_Park_Transform.n614_adj_2017\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17141\,
            carryout => \foc.u_Park_Transform.n17142\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_14_lut_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30281\,
            in2 => \N__34223\,
            in3 => \N__30307\,
            lcout => \foc.u_Park_Transform.n663_adj_2016\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17142\,
            carryout => \foc.u_Park_Transform.n17143\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_15_lut_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34173\,
            in2 => \N__30288\,
            in3 => \N__30292\,
            lcout => \foc.u_Park_Transform.n712_adj_2015\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17143\,
            carryout => \foc.u_Park_Transform.n17144\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_16_lut_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32619\,
            in2 => \N__30289\,
            in3 => \N__30268\,
            lcout => \foc.u_Park_Transform.n770_adj_2030\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17144\,
            carryout => \foc.u_Park_Transform.n771_adj_2032\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n771_adj_2032_THRU_LUT4_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30454\,
            lcout => \foc.u_Park_Transform.n771_adj_2032_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i20_2_lut_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32169\,
            lcout => \foc.u_Park_Transform.n616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i18_2_lut_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32181\,
            lcout => \foc.u_Park_Transform.n613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i525_2_lut_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__32170\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i522_2_lut_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__32182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_2_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44241\,
            in2 => \N__32134\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n87\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \foc.u_Park_Transform.n18160\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_3_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32124\,
            in2 => \N__32029\,
            in3 => \N__30430\,
            lcout => \foc.u_Park_Transform.n136\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n18160\,
            carryout => \foc.u_Park_Transform.n18161\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_4_lut_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32135\,
            in2 => \N__32047\,
            in3 => \N__30427\,
            lcout => \foc.u_Park_Transform.n185\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n18161\,
            carryout => \foc.u_Park_Transform.n18162\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_5_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32125\,
            in2 => \N__34317\,
            in3 => \N__30424\,
            lcout => \foc.u_Park_Transform.n234\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n18162\,
            carryout => \foc.u_Park_Transform.n18163\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_6_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32136\,
            in2 => \N__34360\,
            in3 => \N__30421\,
            lcout => \foc.u_Park_Transform.n283\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n18163\,
            carryout => \foc.u_Park_Transform.n18164\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_7_lut_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34349\,
            in2 => \N__32140\,
            in3 => \N__30508\,
            lcout => \foc.u_Park_Transform.n332\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n18164\,
            carryout => \foc.u_Park_Transform.n18165\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_573_8_lut_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32397\,
            in2 => \N__34361\,
            in3 => \N__30505\,
            lcout => \foc.u_Park_Transform.n786\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n18165\,
            carryout => \foc.u_Park_Transform.n787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n787_THRU_LUT4_0_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30502\,
            lcout => \foc.u_Park_Transform.n787_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_2_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32133\,
            in2 => \N__31788\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n84_adj_2118\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \foc.u_Park_Transform.n16915\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_3_lut_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31772\,
            in2 => \N__30499\,
            in3 => \N__30490\,
            lcout => \foc.u_Park_Transform.n133\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16915\,
            carryout => \foc.u_Park_Transform.n16916\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_4_lut_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31773\,
            in2 => \N__30487\,
            in3 => \N__30478\,
            lcout => \foc.u_Park_Transform.n182\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16916\,
            carryout => \foc.u_Park_Transform.n16917\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_5_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30475\,
            in2 => \N__31789\,
            in3 => \N__30469\,
            lcout => \foc.u_Park_Transform.n231\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16917\,
            carryout => \foc.u_Park_Transform.n16918\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_6_lut_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31777\,
            in2 => \N__30466\,
            in3 => \N__30457\,
            lcout => \foc.u_Park_Transform.n280\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16918\,
            carryout => \foc.u_Park_Transform.n16919\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_7_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30646\,
            in2 => \N__31790\,
            in3 => \N__30640\,
            lcout => \foc.u_Park_Transform.n329\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16919\,
            carryout => \foc.u_Park_Transform.n16920\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_8_lut_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31781\,
            in2 => \N__30627\,
            in3 => \N__30637\,
            lcout => \foc.u_Park_Transform.n378\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16920\,
            carryout => \foc.u_Park_Transform.n16921\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_9_lut_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30623\,
            in2 => \N__31791\,
            in3 => \N__30634\,
            lcout => \foc.u_Park_Transform.n427\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16921\,
            carryout => \foc.u_Park_Transform.n16922\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_572_10_lut_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32011\,
            in2 => \N__30631\,
            in3 => \N__30607\,
            lcout => \foc.u_Park_Transform.n782\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \foc.u_Park_Transform.n783_adj_2167\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n783_adj_2167_THRU_LUT4_0_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30604\,
            lcout => \foc.u_Park_Transform.n783_adj_2167_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_2_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31792\,
            in2 => \N__30845\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n81_adj_2120\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \foc.u_Park_Transform.n16924\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_3_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30820\,
            in2 => \N__30589\,
            in3 => \N__30562\,
            lcout => \foc.u_Park_Transform.n130_adj_2105\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16924\,
            carryout => \foc.u_Park_Transform.n16925\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_4_lut_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30821\,
            in2 => \N__30559\,
            in3 => \N__30535\,
            lcout => \foc.u_Park_Transform.n179_adj_2076\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16925\,
            carryout => \foc.u_Park_Transform.n16926\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_5_lut_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30532\,
            in2 => \N__30846\,
            in3 => \N__30511\,
            lcout => \foc.u_Park_Transform.n228\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16926\,
            carryout => \foc.u_Park_Transform.n16927\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_6_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30825\,
            in2 => \N__30967\,
            in3 => \N__30940\,
            lcout => \foc.u_Park_Transform.n277\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16927\,
            carryout => \foc.u_Park_Transform.n16928\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_7_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30937\,
            in2 => \N__30847\,
            in3 => \N__30916\,
            lcout => \foc.u_Park_Transform.n326\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16928\,
            carryout => \foc.u_Park_Transform.n16929\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_8_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30829\,
            in2 => \N__30913\,
            in3 => \N__30886\,
            lcout => \foc.u_Park_Transform.n375\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16929\,
            carryout => \foc.u_Park_Transform.n16930\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_9_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30883\,
            in2 => \N__30848\,
            in3 => \N__30868\,
            lcout => \foc.u_Park_Transform.n424\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16930\,
            carryout => \foc.u_Park_Transform.n16931\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_10_lut_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30833\,
            in2 => \N__30672\,
            in3 => \N__30853\,
            lcout => \foc.u_Park_Transform.n473\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \foc.u_Park_Transform.n16932\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_11_lut_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30668\,
            in2 => \N__30849\,
            in3 => \N__30694\,
            lcout => \foc.u_Park_Transform.n522\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16932\,
            carryout => \foc.u_Park_Transform.n16933\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_571_12_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30691\,
            in2 => \N__30673\,
            in3 => \N__30652\,
            lcout => \foc.u_Park_Transform.n778\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16933\,
            carryout => \foc.u_Park_Transform.n779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n779_THRU_LUT4_0_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30649\,
            lcout => \foc.u_Park_Transform.n779_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_2_lut_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31287\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2417\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_3_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34779\,
            in2 => \N__31129\,
            in3 => \N__30991\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2517\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_4_lut_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31114\,
            in2 => \N__34795\,
            in3 => \N__30988\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2617\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_5_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34783\,
            in2 => \N__31099\,
            in3 => \N__30985\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2717\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_6_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31081\,
            in2 => \N__34796\,
            in3 => \N__30982\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2817\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_7_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34787\,
            in2 => \N__31069\,
            in3 => \N__30979\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2917\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_8_lut_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31348\,
            in2 => \N__34797\,
            in3 => \N__30976\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3017\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_9_lut_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34791\,
            in2 => \N__31336\,
            in3 => \N__30973\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3117\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17392\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_10_lut_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31276\,
            in2 => \_gnd_net_\,
            in3 => \N__30970\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3223\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_LUT4_0_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31054\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_2_lut_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31173\,
            in2 => \N__32738\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2329\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_3_lut_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31051\,
            in2 => \_gnd_net_\,
            in3 => \N__31045\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2429\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_4_lut_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31174\,
            in2 => \N__31042\,
            in3 => \N__31033\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2529\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_5_lut_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31030\,
            in2 => \N__31191\,
            in3 => \N__31024\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2629\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_6_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31178\,
            in2 => \N__31021\,
            in3 => \N__31012\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2729\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_7_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31009\,
            in2 => \N__31192\,
            in3 => \N__31003\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2829\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_8_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31000\,
            in2 => \N__31194\,
            in3 => \N__30994\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2929\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_9_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31210\,
            in2 => \N__31193\,
            in3 => \N__31204\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3029\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17428\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_10_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31201\,
            in2 => \N__31195\,
            in3 => \N__31144\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3129\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_11_lut_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31141\,
            in2 => \_gnd_net_\,
            in3 => \N__31135\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3239\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_LUT4_0_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31132\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_2_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33495\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2420\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_3_lut_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31306\,
            in2 => \N__33295\,
            in3 => \N__31102\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2520\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_4_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33640\,
            in2 => \N__31319\,
            in3 => \N__31084\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2620\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_5_lut_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31310\,
            in2 => \N__33622\,
            in3 => \N__31072\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2720\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_6_lut_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33598\,
            in2 => \N__31320\,
            in3 => \N__31057\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2820\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_7_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31314\,
            in2 => \N__33580\,
            in3 => \N__31339\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2920\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_8_lut_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33556\,
            in2 => \N__31321\,
            in3 => \N__31324\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3020\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_9_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31318\,
            in2 => \N__33538\,
            in3 => \N__31267\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3120\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17401\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_10_lut_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33457\,
            in2 => \_gnd_net_\,
            in3 => \N__31264\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3227\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_LUT4_0_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31261\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_i1719_2_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31439\,
            in2 => \N__32805\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_3_lut_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31258\,
            in2 => \_gnd_net_\,
            in3 => \N__31237\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7472\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_4_lut_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31440\,
            in2 => \N__31234\,
            in3 => \N__31213\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7471\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_5_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31447\,
            in2 => \N__31681\,
            in3 => \N__31663\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7470\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_6_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31660\,
            in2 => \N__31493\,
            in3 => \N__31642\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7469\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_7_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31639\,
            in2 => \N__31491\,
            in3 => \N__31624\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7468\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_8_lut_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31621\,
            in2 => \N__31494\,
            in3 => \N__31603\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7467\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_9_lut_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31600\,
            in2 => \N__31492\,
            in3 => \N__31585\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7466\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17357\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_10_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__31457\,
            in2 => \_gnd_net_\,
            in3 => \N__31384\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_2_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32117\,
            in2 => \N__31733\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n84\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \foc.u_Park_Transform.n17098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_3_lut_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31714\,
            in2 => \N__31993\,
            in3 => \N__31351\,
            lcout => \foc.u_Park_Transform.n133_adj_2101\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17098\,
            carryout => \foc.u_Park_Transform.n17099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31715\,
            in2 => \N__31981\,
            in3 => \N__31888\,
            lcout => \foc.u_Park_Transform.n182_adj_2094\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17099\,
            carryout => \foc.u_Park_Transform.n17100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_5_lut_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31966\,
            in2 => \N__31734\,
            in3 => \N__31873\,
            lcout => \foc.u_Park_Transform.n231_adj_2089\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17100\,
            carryout => \foc.u_Park_Transform.n17101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_6_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31719\,
            in2 => \N__31954\,
            in3 => \N__31858\,
            lcout => \foc.u_Park_Transform.n280_adj_2087\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17101\,
            carryout => \foc.u_Park_Transform.n17102\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_7_lut_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31939\,
            in2 => \N__31735\,
            in3 => \N__31840\,
            lcout => \foc.u_Park_Transform.n329_adj_2080\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17102\,
            carryout => \foc.u_Park_Transform.n17103\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_8_lut_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31723\,
            in2 => \N__31927\,
            in3 => \N__31828\,
            lcout => \foc.u_Park_Transform.n378_adj_2078\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17103\,
            carryout => \foc.u_Park_Transform.n17104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_9_lut_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31926\,
            in2 => \N__31736\,
            in3 => \N__31801\,
            lcout => \foc.u_Park_Transform.n427_adj_2069\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17104\,
            carryout => \foc.u_Park_Transform.n17105\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_10_lut_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32004\,
            in2 => \N__31922\,
            in3 => \N__31798\,
            lcout => \foc.u_Park_Transform.n782_adj_2109\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \foc.u_Park_Transform.n783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n783_THRU_LUT4_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31795\,
            lcout => \foc.u_Park_Transform.n783_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i24_2_lut_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32445\,
            lcout => \foc.u_Park_Transform.n622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i531_2_lut_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__32446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_2_lut_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44254\,
            in2 => \N__32113\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n87_adj_2138\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \foc.u_Park_Transform.n17980\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_3_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32022\,
            in2 => \N__32115\,
            in3 => \N__31969\,
            lcout => \foc.u_Park_Transform.n136_adj_2127\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17980\,
            carryout => \foc.u_Park_Transform.n17981\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_4_lut_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32040\,
            in2 => \N__32114\,
            in3 => \N__31957\,
            lcout => \foc.u_Park_Transform.n185_adj_2126\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17981\,
            carryout => \foc.u_Park_Transform.n17982\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_5_lut_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32089\,
            in2 => \N__34321\,
            in3 => \N__31942\,
            lcout => \foc.u_Park_Transform.n234_adj_2125\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17982\,
            carryout => \foc.u_Park_Transform.n17983\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_6_lut_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32093\,
            in2 => \N__34362\,
            in3 => \N__31930\,
            lcout => \foc.u_Park_Transform.n283_adj_2122\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17983\,
            carryout => \foc.u_Park_Transform.n17984\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_7_lut_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34356\,
            in2 => \N__32116\,
            in3 => \N__31903\,
            lcout => \foc.u_Park_Transform.n332_adj_2110\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17984\,
            carryout => \foc.u_Park_Transform.n17985\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_8_lut_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32404\,
            in2 => \N__34363\,
            in3 => \N__31900\,
            lcout => \foc.u_Park_Transform.n786_adj_2152\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17985\,
            carryout => \foc.u_Park_Transform.n787_adj_2149\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n787_adj_2149_THRU_LUT4_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32143\,
            lcout => \foc.u_Park_Transform.n787_adj_2149_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i519_2_lut_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__32194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i26_2_lut_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32419\,
            lcout => \foc.u_Park_Transform.n625\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16567_2_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__40485\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44410\,
            lcout => OPEN,
            ltout => \n21486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100101101010"
        )
    port map (
            in0 => \N__44253\,
            in1 => \_gnd_net_\,
            in2 => \N__32050\,
            in3 => \N__40446\,
            lcout => n139,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i14_2_lut_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32205\,
            lcout => \foc.u_Park_Transform.n607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i516_2_lut_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__32206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i11560_3_lut_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__40484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44409\,
            lcout => \foc.u_Park_Transform.n90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i16_2_lut_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32193\,
            lcout => \foc.u_Park_Transform.n610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_2_lut_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32641\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.Look_Up_Table_out1_1_2\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_3_lut_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33043\,
            in2 => \_gnd_net_\,
            in3 => \N__32215\,
            lcout => \foc.Look_Up_Table_out1_1_3\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_4_lut_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33031\,
            in2 => \_gnd_net_\,
            in3 => \N__32212\,
            lcout => \foc.Look_Up_Table_out1_1_4\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_5_lut_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33013\,
            in2 => \_gnd_net_\,
            in3 => \N__32209\,
            lcout => \foc.Look_Up_Table_out1_1_5\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_6_lut_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32980\,
            in2 => \_gnd_net_\,
            in3 => \N__32197\,
            lcout => \foc.Look_Up_Table_out1_1_6\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_7_lut_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32950\,
            in2 => \_gnd_net_\,
            in3 => \N__32185\,
            lcout => \foc.Look_Up_Table_out1_1_7\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_8_lut_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32935\,
            in2 => \_gnd_net_\,
            in3 => \N__32173\,
            lcout => \foc.Look_Up_Table_out1_1_8\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_9_lut_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32914\,
            in2 => \_gnd_net_\,
            in3 => \N__32161\,
            lcout => \foc.Look_Up_Table_out1_1_9\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15951\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_10_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32878\,
            in2 => \_gnd_net_\,
            in3 => \N__32146\,
            lcout => \foc.Look_Up_Table_out1_1_10\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_11_lut_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33262\,
            in2 => \_gnd_net_\,
            in3 => \N__32434\,
            lcout => \foc.Look_Up_Table_out1_1_11\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_12_lut_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33226\,
            in2 => \_gnd_net_\,
            in3 => \N__32431\,
            lcout => \foc.Look_Up_Table_out1_1_12\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_13_lut_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33181\,
            in2 => \_gnd_net_\,
            in3 => \N__32428\,
            lcout => \Look_Up_Table_out1_1_13\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_14_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33136\,
            in2 => \N__44860\,
            in3 => \N__32425\,
            lcout => \Look_Up_Table_out1_1_14\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15956\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_15_lut_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33091\,
            in2 => \_gnd_net_\,
            in3 => \N__32422\,
            lcout => \Look_Up_Table_out1_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i534_2_lut_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32415\,
            lcout => \foc.u_Park_Transform.n785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_2_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32352\,
            in2 => \N__34276\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n75_adj_2123\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \foc.u_Park_Transform.n16948\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_3_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32242\,
            in2 => \N__34277\,
            in3 => \N__32233\,
            lcout => \foc.u_Park_Transform.n124_adj_2090\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16948\,
            carryout => \foc.u_Park_Transform.n16949\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_4_lut_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34249\,
            in2 => \N__32230\,
            in3 => \N__32218\,
            lcout => \foc.u_Park_Transform.n173_adj_2061\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16949\,
            carryout => \foc.u_Park_Transform.n16950\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_5_lut_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34243\,
            in2 => \N__32578\,
            in3 => \N__32566\,
            lcout => \foc.u_Park_Transform.n222_adj_2049\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16950\,
            carryout => \foc.u_Park_Transform.n16951\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_6_lut_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34250\,
            in2 => \N__32563\,
            in3 => \N__32551\,
            lcout => \foc.u_Park_Transform.n271_adj_2043\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16951\,
            carryout => \foc.u_Park_Transform.n16952\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_7_lut_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34244\,
            in2 => \N__32548\,
            in3 => \N__32536\,
            lcout => \foc.u_Park_Transform.n320_adj_2036\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16952\,
            carryout => \foc.u_Park_Transform.n16953\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_8_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34251\,
            in2 => \N__32533\,
            in3 => \N__32521\,
            lcout => \foc.u_Park_Transform.n369_adj_2026\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16953\,
            carryout => \foc.u_Park_Transform.n16954\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_9_lut_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34245\,
            in2 => \N__32518\,
            in3 => \N__32506\,
            lcout => \foc.u_Park_Transform.n418\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16954\,
            carryout => \foc.u_Park_Transform.n16955\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_10_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34280\,
            in2 => \N__32503\,
            in3 => \N__32488\,
            lcout => \foc.u_Park_Transform.n467\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \foc.u_Park_Transform.n16956\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_11_lut_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32485\,
            in2 => \N__34292\,
            in3 => \N__32476\,
            lcout => \foc.u_Park_Transform.n516\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16956\,
            carryout => \foc.u_Park_Transform.n16957\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_12_lut_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34284\,
            in2 => \N__32473\,
            in3 => \N__32461\,
            lcout => \foc.u_Park_Transform.n565_adj_2020\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16957\,
            carryout => \foc.u_Park_Transform.n16958\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_13_lut_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32458\,
            in2 => \N__34293\,
            in3 => \N__32449\,
            lcout => \foc.u_Park_Transform.n614\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16958\,
            carryout => \foc.u_Park_Transform.n16959\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_14_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32600\,
            in2 => \N__34294\,
            in3 => \N__32629\,
            lcout => \foc.u_Park_Transform.n663\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16959\,
            carryout => \foc.u_Park_Transform.n16960\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_15_lut_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34291\,
            in2 => \N__32607\,
            in3 => \N__32626\,
            lcout => \foc.u_Park_Transform.n712\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16960\,
            carryout => \foc.u_Park_Transform.n16961\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_569_16_lut_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32623\,
            in2 => \N__32608\,
            in3 => \N__32584\,
            lcout => \foc.u_Park_Transform.n770\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16961\,
            carryout => \foc.u_Park_Transform.n771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n771_THRU_LUT4_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32581\,
            lcout => \foc.u_Park_Transform.n771_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_2_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36660\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17358\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_3_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32848\,
            in2 => \N__36415\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17358\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17359\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_4_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36388\,
            in2 => \N__32861\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17359\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17360\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_5_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32852\,
            in2 => \N__36364\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17360\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17361\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_6_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36334\,
            in2 => \N__32862\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17361\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17362\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_7_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32856\,
            in2 => \N__36310\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17362\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_8_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36286\,
            in2 => \N__32863\,
            in3 => \N__32866\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3008\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_9_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32860\,
            in2 => \N__36265\,
            in3 => \N__32824\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3108\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17365\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_10_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36622\,
            in2 => \_gnd_net_\,
            in3 => \N__32821\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3211\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_LUT4_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32818\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_2_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32815\,
            in2 => \N__32804\,
            in3 => \_gnd_net_\,
            lcout => \foc.Look_Up_Table_out1_1_0\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_3_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32659\,
            in2 => \_gnd_net_\,
            in3 => \N__32650\,
            lcout => \foc.Look_Up_Table_out1_1_1\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_4_lut_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32647\,
            in2 => \_gnd_net_\,
            in3 => \N__32632\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_34\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_5_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36601\,
            in2 => \N__33052\,
            in3 => \N__33034\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_35\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_6_lut_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34837\,
            in2 => \N__36583\,
            in3 => \N__33022\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_36\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_7_lut_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33019\,
            in2 => \N__34825\,
            in3 => \N__33004\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_37\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_8_lut_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33001\,
            in2 => \N__32989\,
            in3 => \N__32968\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_38\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_9_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33439\,
            in2 => \N__32965\,
            in3 => \N__32938\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_39\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17497\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_10_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33376\,
            in2 => \N__33748\,
            in3 => \N__32926\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_40\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_11_lut_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32923\,
            in2 => \N__33361\,
            in3 => \N__32905\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_41\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_12_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32902\,
            in2 => \N__32890\,
            in3 => \N__32869\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_42\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_13_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33286\,
            in2 => \N__33277\,
            in3 => \N__33253\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_43\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_14_lut_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33250\,
            in2 => \N__33238\,
            in3 => \N__33214\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_44\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_15_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33211\,
            in2 => \N__33196\,
            in3 => \N__33169\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_45\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_16_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33166\,
            in2 => \N__33154\,
            in3 => \N__33124\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_46\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17504\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_17_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33121\,
            in1 => \N__33106\,
            in2 => \_gnd_net_\,
            in3 => \N__33094\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_2_lut_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33079\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2426\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_3_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33327\,
            in2 => \N__33073\,
            in3 => \N__33064\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2526\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_4_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33061\,
            in2 => \N__33345\,
            in3 => \N__33055\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2626\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_5_lut_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33331\,
            in2 => \N__33430\,
            in3 => \N__33421\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2726\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_6_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33418\,
            in2 => \N__33346\,
            in3 => \N__33412\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2826\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_7_lut_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33409\,
            in2 => \N__33348\,
            in3 => \N__33403\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2926\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_8_lut_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33400\,
            in2 => \N__33347\,
            in3 => \N__33394\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3026\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_9_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33391\,
            in2 => \N__33349\,
            in3 => \N__33385\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3126\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17419\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_10_lut_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33382\,
            in2 => \_gnd_net_\,
            in3 => \N__33367\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3235\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_LUT4_0_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33364\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_2_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33344\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2423\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_3_lut_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33496\,
            in2 => \N__33652\,
            in3 => \N__33634\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2523\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_4_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33631\,
            in2 => \N__33513\,
            in3 => \N__33613\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2623\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_5_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33500\,
            in2 => \N__33610\,
            in3 => \N__33592\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2723\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_6_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33589\,
            in2 => \N__33514\,
            in3 => \N__33568\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2823\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_7_lut_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33565\,
            in2 => \N__33516\,
            in3 => \N__33550\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2923\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_8_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33547\,
            in2 => \N__33515\,
            in3 => \N__33529\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3023\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_9_lut_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33526\,
            in2 => \N__33517\,
            in3 => \N__33451\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3123\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17410\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_10_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33448\,
            in2 => \_gnd_net_\,
            in3 => \N__33754\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3231\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_LUT4_0_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33751\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_2_lut_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35813\,
            in2 => \N__36133\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n69\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \foc.u_Park_Transform.n17161\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_3_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36124\,
            in2 => \N__33736\,
            in3 => \N__33724\,
            lcout => \foc.u_Park_Transform.n118\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17161\,
            carryout => \foc.u_Park_Transform.n17162\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_4_lut_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36029\,
            in2 => \N__33721\,
            in3 => \N__33709\,
            lcout => \foc.u_Park_Transform.n167\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17162\,
            carryout => \foc.u_Park_Transform.n17163\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_5_lut_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33706\,
            in2 => \N__36082\,
            in3 => \N__33697\,
            lcout => \foc.u_Park_Transform.n216\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17163\,
            carryout => \foc.u_Park_Transform.n17164\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_6_lut_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36033\,
            in2 => \N__33694\,
            in3 => \N__33682\,
            lcout => \foc.u_Park_Transform.n265\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17164\,
            carryout => \foc.u_Park_Transform.n17165\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_7_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33679\,
            in2 => \N__36083\,
            in3 => \N__33670\,
            lcout => \foc.u_Park_Transform.n314\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17165\,
            carryout => \foc.u_Park_Transform.n17166\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_8_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36037\,
            in2 => \N__33667\,
            in3 => \N__33655\,
            lcout => \foc.u_Park_Transform.n363\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17166\,
            carryout => \foc.u_Park_Transform.n17167\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_9_lut_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33862\,
            in2 => \N__36084\,
            in3 => \N__33853\,
            lcout => \foc.u_Park_Transform.n412\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17167\,
            carryout => \foc.u_Park_Transform.n17168\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_10_lut_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33850\,
            in2 => \N__36078\,
            in3 => \N__33838\,
            lcout => \foc.u_Park_Transform.n461\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \foc.u_Park_Transform.n17169\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_11_lut_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36018\,
            in2 => \N__33835\,
            in3 => \N__33823\,
            lcout => \foc.u_Park_Transform.n510_adj_2004\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17169\,
            carryout => \foc.u_Park_Transform.n17170\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_12_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33820\,
            in2 => \N__36079\,
            in3 => \N__33811\,
            lcout => \foc.u_Park_Transform.n559_adj_2001\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17170\,
            carryout => \foc.u_Park_Transform.n17171\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_13_lut_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36022\,
            in2 => \N__33808\,
            in3 => \N__33796\,
            lcout => \foc.u_Park_Transform.n608\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17171\,
            carryout => \foc.u_Park_Transform.n17172\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_14_lut_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33793\,
            in2 => \N__36080\,
            in3 => \N__33784\,
            lcout => \foc.u_Park_Transform.n657\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17172\,
            carryout => \foc.u_Park_Transform.n17173\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_15_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33781\,
            in2 => \N__36081\,
            in3 => \N__33772\,
            lcout => \foc.u_Park_Transform.n706\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17173\,
            carryout => \foc.u_Park_Transform.n17174\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_16_lut_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35934\,
            in2 => \N__33769\,
            in3 => \N__33757\,
            lcout => \foc.u_Park_Transform.n762\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17174\,
            carryout => \foc.u_Park_Transform.n763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n763_THRU_LUT4_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33961\,
            lcout => \foc.u_Park_Transform.n763_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_2_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35976\,
            in2 => \N__37759\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n66\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \foc.u_Park_Transform.n17176\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_3_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37736\,
            in2 => \N__33958\,
            in3 => \N__33946\,
            lcout => \foc.u_Park_Transform.n115\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17176\,
            carryout => \foc.u_Park_Transform.n17177\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_4_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37737\,
            in2 => \N__33943\,
            in3 => \N__33931\,
            lcout => \foc.u_Park_Transform.n164\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17177\,
            carryout => \foc.u_Park_Transform.n17178\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_5_lut_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33928\,
            in2 => \N__37760\,
            in3 => \N__33919\,
            lcout => \foc.u_Park_Transform.n213\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17178\,
            carryout => \foc.u_Park_Transform.n17179\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_6_lut_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37741\,
            in2 => \N__33916\,
            in3 => \N__33904\,
            lcout => \foc.u_Park_Transform.n262_adj_1996\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17179\,
            carryout => \foc.u_Park_Transform.n17180\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_7_lut_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33901\,
            in2 => \N__37761\,
            in3 => \N__33892\,
            lcout => \foc.u_Park_Transform.n311\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17180\,
            carryout => \foc.u_Park_Transform.n17181\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_8_lut_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37745\,
            in2 => \N__33889\,
            in3 => \N__33877\,
            lcout => \foc.u_Park_Transform.n360\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17181\,
            carryout => \foc.u_Park_Transform.n17182\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_9_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33874\,
            in2 => \N__37762\,
            in3 => \N__33865\,
            lcout => \foc.u_Park_Transform.n409\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17182\,
            carryout => \foc.u_Park_Transform.n17183\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_10_lut_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37643\,
            in2 => \N__34057\,
            in3 => \N__34045\,
            lcout => \foc.u_Park_Transform.n458\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \foc.u_Park_Transform.n17184\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_11_lut_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34042\,
            in2 => \N__37713\,
            in3 => \N__34033\,
            lcout => \foc.u_Park_Transform.n507_adj_2165\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17184\,
            carryout => \foc.u_Park_Transform.n17185\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_12_lut_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37647\,
            in2 => \N__34030\,
            in3 => \N__34018\,
            lcout => \foc.u_Park_Transform.n556_adj_2164\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17185\,
            carryout => \foc.u_Park_Transform.n17186\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_13_lut_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34015\,
            in2 => \N__37714\,
            in3 => \N__34006\,
            lcout => \foc.u_Park_Transform.n605_adj_2163\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17186\,
            carryout => \foc.u_Park_Transform.n17187\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_14_lut_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34003\,
            in2 => \N__37716\,
            in3 => \N__33994\,
            lcout => \foc.u_Park_Transform.n654_adj_2162\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17187\,
            carryout => \foc.u_Park_Transform.n17188\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_15_lut_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33991\,
            in2 => \N__37715\,
            in3 => \N__33982\,
            lcout => \foc.u_Park_Transform.n703_adj_2160\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17188\,
            carryout => \foc.u_Park_Transform.n17189\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_16_lut_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35541\,
            in2 => \N__33979\,
            in3 => \N__33967\,
            lcout => \foc.u_Park_Transform.n758_adj_2168\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17189\,
            carryout => \foc.u_Park_Transform.n759_adj_2166\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n759_adj_2166_THRU_LUT4_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33964\,
            lcout => \foc.u_Park_Transform.n759_adj_2166_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i8_2_lut_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34083\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i507_2_lut_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__34084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i510_2_lut_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__34066\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i504_2_lut_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__42714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i513_2_lut_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__34075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i12_2_lut_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34074\,
            lcout => \foc.u_Park_Transform.n604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.u_29__I_0_71_inv_0_i4_1_lut_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Amp25_out1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i10_2_lut_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34065\,
            lcout => \foc.u_Park_Transform.n601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i498_2_lut_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36568\,
            lcout => \foc.u_Park_Transform.n737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i2_4_lut_4_lut_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010110100"
        )
    port map (
            in0 => \N__44188\,
            in1 => \N__44317\,
            in2 => \_gnd_net_\,
            in3 => \N__44394\,
            lcout => \foc.u_Park_Transform.n790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11567_4_lut_4_lut_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__44395\,
            in1 => \N__44240\,
            in2 => \_gnd_net_\,
            in3 => \N__40475\,
            lcout => n4,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_3_lut_4_lut_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44315\,
            in2 => \N__34366\,
            in3 => \N__44392\,
            lcout => \foc.u_Park_Transform.n237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i2_2_lut_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36567\,
            lcout => \foc.u_Park_Transform.dCurrent_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i2_3_lut_4_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__42507\,
            in1 => \N__44316\,
            in2 => \_gnd_net_\,
            in3 => \N__44393\,
            lcout => \foc.u_Park_Transform.n188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_2_lut_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34279\,
            in2 => \N__35883\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n72_adj_2062\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \foc.u_Park_Transform.n16963\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_3_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34126\,
            in2 => \N__35884\,
            in3 => \N__34120\,
            lcout => \foc.u_Park_Transform.n121_adj_2051\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16963\,
            carryout => \foc.u_Park_Transform.n16964\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_4_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35838\,
            in2 => \N__34117\,
            in3 => \N__34108\,
            lcout => \foc.u_Park_Transform.n170_adj_2048\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16964\,
            carryout => \foc.u_Park_Transform.n16965\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_5_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34105\,
            in2 => \N__35885\,
            in3 => \N__34099\,
            lcout => \foc.u_Park_Transform.n219_adj_2040\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16965\,
            carryout => \foc.u_Park_Transform.n16966\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_6_lut_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35842\,
            in2 => \N__34096\,
            in3 => \N__34087\,
            lcout => \foc.u_Park_Transform.n268_adj_2027\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16966\,
            carryout => \foc.u_Park_Transform.n16967\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_7_lut_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34453\,
            in2 => \N__35886\,
            in3 => \N__34447\,
            lcout => \foc.u_Park_Transform.n317_adj_2021\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16967\,
            carryout => \foc.u_Park_Transform.n16968\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_8_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35846\,
            in2 => \N__34444\,
            in3 => \N__34435\,
            lcout => \foc.u_Park_Transform.n366_adj_2013\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16968\,
            carryout => \foc.u_Park_Transform.n16969\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_9_lut_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34432\,
            in2 => \N__35887\,
            in3 => \N__34426\,
            lcout => \foc.u_Park_Transform.n415\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16969\,
            carryout => \foc.u_Park_Transform.n16970\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_10_lut_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35850\,
            in2 => \N__34423\,
            in3 => \N__34414\,
            lcout => \foc.u_Park_Transform.n464\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \foc.u_Park_Transform.n16971\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_11_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34411\,
            in2 => \N__35888\,
            in3 => \N__34405\,
            lcout => \foc.u_Park_Transform.n513\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16971\,
            carryout => \foc.u_Park_Transform.n16972\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_12_lut_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35854\,
            in2 => \N__34402\,
            in3 => \N__34393\,
            lcout => \foc.u_Park_Transform.n562\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16972\,
            carryout => \foc.u_Park_Transform.n16973\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_13_lut_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34390\,
            in2 => \N__35889\,
            in3 => \N__34384\,
            lcout => \foc.u_Park_Transform.n611_adj_2107\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16973\,
            carryout => \foc.u_Park_Transform.n16974\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_14_lut_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34381\,
            in2 => \N__35891\,
            in3 => \N__34375\,
            lcout => \foc.u_Park_Transform.n660_adj_2091\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16974\,
            carryout => \foc.u_Park_Transform.n16975\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_15_lut_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34372\,
            in2 => \N__35890\,
            in3 => \N__34507\,
            lcout => \foc.u_Park_Transform.n709_adj_2066\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16975\,
            carryout => \foc.u_Park_Transform.n16976\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_568_16_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34504\,
            in2 => \N__34483\,
            in3 => \N__34474\,
            lcout => \foc.u_Park_Transform.n766_adj_2053\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16976\,
            carryout => \foc.u_Park_Transform.n767_adj_2041\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n767_adj_2041_THRU_LUT4_0_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34471\,
            lcout => \foc.u_Park_Transform.n767_adj_2041_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_1_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37989\,
            in2 => \N__37993\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \foc.u_Park_Transform.n16900\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_2_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40447\,
            in2 => \_gnd_net_\,
            in3 => \N__34468\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_15\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16900\,
            carryout => \foc.u_Park_Transform.n16901\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_3_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40141\,
            in2 => \N__37966\,
            in3 => \N__34465\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16901\,
            carryout => \foc.u_Park_Transform.n16902\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_4_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42763\,
            in2 => \N__40123\,
            in3 => \N__34462\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_17\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16902\,
            carryout => \foc.u_Park_Transform.n16903\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_5_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39931\,
            in2 => \N__42745\,
            in3 => \N__34459\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16903\,
            carryout => \foc.u_Park_Transform.n16904\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_6_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37813\,
            in2 => \N__40105\,
            in3 => \N__34456\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_19\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16904\,
            carryout => \foc.u_Park_Transform.n16905\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_7_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35530\,
            in2 => \N__37795\,
            in3 => \N__34678\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_20\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16905\,
            carryout => \foc.u_Park_Transform.n16906\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_8_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35515\,
            in2 => \N__35908\,
            in3 => \N__34675\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16906\,
            carryout => \foc.u_Park_Transform.n16907\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_9_lut_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34672\,
            in2 => \N__36487\,
            in3 => \N__34663\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_22\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \foc.u_Park_Transform.n16908\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_10_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34660\,
            in2 => \N__34651\,
            in3 => \N__34639\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16908\,
            carryout => \foc.u_Park_Transform.n16909\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_11_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34636\,
            in2 => \N__34624\,
            in3 => \N__34612\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16909\,
            carryout => \foc.u_Park_Transform.n16910\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_12_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34609\,
            in2 => \N__34600\,
            in3 => \N__34585\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_25\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16910\,
            carryout => \foc.u_Park_Transform.n16911\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_13_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34582\,
            in2 => \N__34570\,
            in3 => \N__34558\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16911\,
            carryout => \foc.u_Park_Transform.n16912\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_14_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34555\,
            in2 => \N__34543\,
            in3 => \N__34528\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_27\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16912\,
            carryout => \foc.u_Park_Transform.n16913\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_15_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35316\,
            in2 => \N__34525\,
            in3 => \N__34510\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_28\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16913\,
            carryout => \foc.u_Park_Transform.n16914\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1232_16_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36537\,
            in1 => \N__44467\,
            in2 => \_gnd_net_\,
            in3 => \N__34801\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_2_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34798\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2414\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_3_lut_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36447\,
            in2 => \N__34756\,
            in3 => \N__34744\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2514\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_4_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34741\,
            in2 => \N__36467\,
            in3 => \N__34732\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2614\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_5_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36451\,
            in2 => \N__34729\,
            in3 => \N__34717\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2714\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_6_lut_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34714\,
            in2 => \N__36468\,
            in3 => \N__34705\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2814\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_7_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34702\,
            in2 => \N__36470\,
            in3 => \N__34693\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2914\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_8_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34690\,
            in2 => \N__36469\,
            in3 => \N__34681\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3014\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_9_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34861\,
            in2 => \N__36471\,
            in3 => \N__34852\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3114\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17383\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_10_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34849\,
            in2 => \_gnd_net_\,
            in3 => \N__34831\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3219\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_LUT4_0_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34828\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66260\,
            in2 => \N__66515\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n78_adj_617\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36526\,
            in2 => \N__66517\,
            in3 => \N__34816\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n127_adj_615\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17656\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17657\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66464\,
            in2 => \N__36517\,
            in3 => \N__34813\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n176_adj_613\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17657\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17658\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36502\,
            in2 => \N__66518\,
            in3 => \N__34810\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n225_adj_611\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17658\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17659\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66468\,
            in2 => \N__36802\,
            in3 => \N__34807\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n274_adj_609\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17659\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17660\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36787\,
            in2 => \N__66519\,
            in3 => \N__34804\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n323_adj_607\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17660\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17661\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36772\,
            in2 => \N__66516\,
            in3 => \N__34885\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n372\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17661\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17662\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36760\,
            in2 => \N__66520\,
            in3 => \N__34882\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n421\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17662\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17663\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36745\,
            in2 => \N__66574\,
            in3 => \N__34879\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n470\,
            ltout => OPEN,
            carryin => \bfn_12_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17664\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36733\,
            in2 => \N__66575\,
            in3 => \N__34876\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n519\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17664\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17665\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66534\,
            in2 => \N__36720\,
            in3 => \N__34873\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n568\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17665\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17666\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36716\,
            in2 => \N__66576\,
            in3 => \N__34870\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n617\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17666\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17667\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45457\,
            in2 => \N__36721\,
            in3 => \N__34867\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n774\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17667\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_LUT4_0_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34864\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66538\,
            in2 => \N__66888\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n75_adj_618\,
            ltout => OPEN,
            carryin => \bfn_12_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18107\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34981\,
            in2 => \N__66923\,
            in3 => \N__34972\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n124_adj_616\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18107\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18108\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34969\,
            in2 => \N__66889\,
            in3 => \N__34960\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n173_adj_614\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18108\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18109\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34957\,
            in2 => \N__66924\,
            in3 => \N__34948\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n222_adj_612\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18109\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18110\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34945\,
            in2 => \N__66890\,
            in3 => \N__34936\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n271_adj_610\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18110\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18111\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34933\,
            in2 => \N__66925\,
            in3 => \N__34924\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n320_adj_608\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18111\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18112\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34921\,
            in2 => \N__66891\,
            in3 => \N__34912\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n369_adj_606\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18112\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18113\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34909\,
            in2 => \N__66926\,
            in3 => \N__34900\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n418_adj_605\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18113\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18114\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34897\,
            in2 => \N__66927\,
            in3 => \N__34888\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n467_adj_604\,
            ltout => OPEN,
            carryin => \bfn_12_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18115\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35053\,
            in2 => \N__66930\,
            in3 => \N__35044\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n516_adj_603\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18115\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18116\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35041\,
            in2 => \N__66928\,
            in3 => \N__35032\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n565_adj_602\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18116\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18117\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35029\,
            in2 => \N__66931\,
            in3 => \N__35020\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n614_adj_601\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18117\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18118\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35003\,
            in2 => \N__66929\,
            in3 => \N__35017\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n663_adj_600\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18118\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18119\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66913\,
            in2 => \N__35010\,
            in3 => \N__35014\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n712_adj_599\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18119\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18120\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45484\,
            in2 => \N__35011\,
            in3 => \N__34987\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n770_adj_597\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18120\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_LUT4_0_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34984\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i18_1_lut_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37354\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i20_1_lut_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37318\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n14_adj_517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i21_1_lut_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i22_1_lut_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37282\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n12_adj_516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i23_1_lut_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37264\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i24_1_lut_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37246\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i25_1_lut_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37228\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_1_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39645\,
            in2 => \N__39649\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \foc.u_Park_Transform.n17083\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_2_lut_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40462\,
            in2 => \_gnd_net_\,
            in3 => \N__35065\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_15\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17083\,
            carryout => \foc.u_Park_Transform.n17084\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_3_lut_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39907\,
            in2 => \N__39622\,
            in3 => \N__35062\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17084\,
            carryout => \foc.u_Park_Transform.n17085\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_4_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37483\,
            in2 => \N__39889\,
            in3 => \N__35059\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_17\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17085\,
            carryout => \foc.u_Park_Transform.n17086\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_5_lut_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42256\,
            in2 => \N__37777\,
            in3 => \N__35056\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17086\,
            carryout => \foc.u_Park_Transform.n17087\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_6_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35494\,
            in2 => \N__42238\,
            in3 => \N__35236\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_19\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17087\,
            carryout => \foc.u_Park_Transform.n17088\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_7_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35233\,
            in2 => \N__35479\,
            in3 => \N__35221\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_20\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17088\,
            carryout => \foc.u_Park_Transform.n17089\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_8_lut_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35218\,
            in2 => \N__35206\,
            in3 => \N__35197\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17089\,
            carryout => \foc.u_Park_Transform.n17090\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_9_lut_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35194\,
            in2 => \N__35185\,
            in3 => \N__35176\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_22\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \foc.u_Park_Transform.n17091\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_10_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35173\,
            in2 => \N__35161\,
            in3 => \N__35149\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17091\,
            carryout => \foc.u_Park_Transform.n17092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_11_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35146\,
            in2 => \N__35134\,
            in3 => \N__35119\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17092\,
            carryout => \foc.u_Park_Transform.n17093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_12_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35116\,
            in2 => \N__35107\,
            in3 => \N__35092\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_25\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17093\,
            carryout => \foc.u_Park_Transform.n17094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_13_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35089\,
            in2 => \N__35080\,
            in3 => \N__35068\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17094\,
            carryout => \foc.u_Park_Transform.n17095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_14_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35350\,
            in2 => \N__35338\,
            in3 => \N__35326\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_27\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17095\,
            carryout => \foc.u_Park_Transform.n17096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_15_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35323\,
            in2 => \N__35302\,
            in3 => \N__35287\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_28\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17096\,
            carryout => \foc.u_Park_Transform.n17097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_1234_16_lut_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44463\,
            in1 => \N__36544\,
            in2 => \_gnd_net_\,
            in3 => \N__35284\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_2_lut_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37754\,
            in2 => \N__41690\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n63_adj_2158\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \foc.u_Park_Transform.n17191\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_3_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35281\,
            in2 => \N__41691\,
            in3 => \N__35275\,
            lcout => \foc.u_Park_Transform.n112_adj_2157\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17191\,
            carryout => \foc.u_Park_Transform.n17192\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_4_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41666\,
            in2 => \N__35272\,
            in3 => \N__35263\,
            lcout => \foc.u_Park_Transform.n161_adj_2156\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17192\,
            carryout => \foc.u_Park_Transform.n17193\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_5_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41660\,
            in2 => \N__35260\,
            in3 => \N__35251\,
            lcout => \foc.u_Park_Transform.n210_adj_2155\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17193\,
            carryout => \foc.u_Park_Transform.n17194\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_6_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41667\,
            in2 => \N__35248\,
            in3 => \N__35239\,
            lcout => \foc.u_Park_Transform.n259_adj_2154\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17194\,
            carryout => \foc.u_Park_Transform.n17195\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_7_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41661\,
            in2 => \N__35449\,
            in3 => \N__35440\,
            lcout => \foc.u_Park_Transform.n308_adj_2153\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17195\,
            carryout => \foc.u_Park_Transform.n17196\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_8_lut_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41668\,
            in2 => \N__35437\,
            in3 => \N__35428\,
            lcout => \foc.u_Park_Transform.n357_adj_2151\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17196\,
            carryout => \foc.u_Park_Transform.n17197\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_9_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41662\,
            in2 => \N__35425\,
            in3 => \N__35416\,
            lcout => \foc.u_Park_Transform.n406_adj_2150\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17197\,
            carryout => \foc.u_Park_Transform.n17198\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_10_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35413\,
            in2 => \N__41651\,
            in3 => \N__35407\,
            lcout => \foc.u_Park_Transform.n455_adj_2148\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \foc.u_Park_Transform.n17199\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_11_lut_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41600\,
            in2 => \N__35404\,
            in3 => \N__35395\,
            lcout => \foc.u_Park_Transform.n504_adj_2147\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17199\,
            carryout => \foc.u_Park_Transform.n17200\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_12_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35392\,
            in2 => \N__41652\,
            in3 => \N__35386\,
            lcout => \foc.u_Park_Transform.n553_adj_2146\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17200\,
            carryout => \foc.u_Park_Transform.n17201\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_13_lut_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41604\,
            in2 => \N__35383\,
            in3 => \N__35374\,
            lcout => \foc.u_Park_Transform.n602_adj_2144\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17201\,
            carryout => \foc.u_Park_Transform.n17202\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_14_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35371\,
            in2 => \N__41653\,
            in3 => \N__35365\,
            lcout => \foc.u_Park_Transform.n651_adj_2143\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17202\,
            carryout => \foc.u_Park_Transform.n17203\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_15_lut_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41608\,
            in2 => \N__35362\,
            in3 => \N__35353\,
            lcout => \foc.u_Park_Transform.n700_adj_2141\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17203\,
            carryout => \foc.u_Park_Transform.n17204\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_16_lut_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37833\,
            in2 => \N__35503\,
            in3 => \N__35485\,
            lcout => \foc.u_Park_Transform.n754_adj_2159\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17204\,
            carryout => \foc.u_Park_Transform.n755_adj_2161\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n755_adj_2161_THRU_LUT4_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35482\,
            lcout => \foc.u_Park_Transform.n755_adj_2161_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_2_lut_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36085\,
            in2 => \N__37755\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n66_adj_2033\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \foc.u_Park_Transform.n16993\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_3_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37720\,
            in2 => \N__35707\,
            in3 => \N__35467\,
            lcout => \foc.u_Park_Transform.n115_adj_2028\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16993\,
            carryout => \foc.u_Park_Transform.n16994\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_4_lut_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37721\,
            in2 => \N__35689\,
            in3 => \N__35464\,
            lcout => \foc.u_Park_Transform.n164_adj_2014\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16994\,
            carryout => \foc.u_Park_Transform.n16995\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_5_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35665\,
            in2 => \N__37756\,
            in3 => \N__35461\,
            lcout => \foc.u_Park_Transform.n213_adj_1999\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16995\,
            carryout => \foc.u_Park_Transform.n16996\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_6_lut_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37725\,
            in2 => \N__35647\,
            in3 => \N__35458\,
            lcout => \foc.u_Park_Transform.n262\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16996\,
            carryout => \foc.u_Park_Transform.n16997\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_7_lut_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35623\,
            in2 => \N__37757\,
            in3 => \N__35455\,
            lcout => \foc.u_Park_Transform.n311_adj_2022\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16997\,
            carryout => \foc.u_Park_Transform.n16998\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_8_lut_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37729\,
            in2 => \N__35605\,
            in3 => \N__35452\,
            lcout => \foc.u_Park_Transform.n360_adj_2009\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16998\,
            carryout => \foc.u_Park_Transform.n16999\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_9_lut_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35581\,
            in2 => \N__37758\,
            in3 => \N__35563\,
            lcout => \foc.u_Park_Transform.n409_adj_1997\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16999\,
            carryout => \foc.u_Park_Transform.n17000\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_10_lut_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37696\,
            in2 => \N__36250\,
            in3 => \N__35560\,
            lcout => \foc.u_Park_Transform.n458_adj_2093\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \foc.u_Park_Transform.n17001\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_11_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36229\,
            in2 => \N__37750\,
            in3 => \N__35557\,
            lcout => \foc.u_Park_Transform.n507\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17001\,
            carryout => \foc.u_Park_Transform.n17002\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_12_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37700\,
            in2 => \N__36211\,
            in3 => \N__35554\,
            lcout => \foc.u_Park_Transform.n556\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17002\,
            carryout => \foc.u_Park_Transform.n17003\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_13_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36187\,
            in2 => \N__37751\,
            in3 => \N__35551\,
            lcout => \foc.u_Park_Transform.n605\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17003\,
            carryout => \foc.u_Park_Transform.n17004\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_14_lut_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36169\,
            in2 => \N__37753\,
            in3 => \N__35548\,
            lcout => \foc.u_Park_Transform.n654\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17004\,
            carryout => \foc.u_Park_Transform.n17005\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_15_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36151\,
            in2 => \N__37752\,
            in3 => \N__35545\,
            lcout => \foc.u_Park_Transform.n703\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17005\,
            carryout => \foc.u_Park_Transform.n17006\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_566_16_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35542\,
            in2 => \N__35956\,
            in3 => \N__35521\,
            lcout => \foc.u_Park_Transform.n758\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17006\,
            carryout => \foc.u_Park_Transform.n759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n759_THRU_LUT4_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35518\,
            lcout => \foc.u_Park_Transform.n759_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_2_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36091\,
            in2 => \N__35892\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n69_adj_2059\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \foc.u_Park_Transform.n16978\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_3_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35695\,
            in2 => \N__36125\,
            in3 => \N__35677\,
            lcout => \foc.u_Park_Transform.n118_adj_2037\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16978\,
            carryout => \foc.u_Park_Transform.n16979\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_4_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36095\,
            in2 => \N__35674\,
            in3 => \N__35656\,
            lcout => \foc.u_Park_Transform.n167_adj_2029\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16979\,
            carryout => \foc.u_Park_Transform.n16980\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_5_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35653\,
            in2 => \N__36126\,
            in3 => \N__35635\,
            lcout => \foc.u_Park_Transform.n216_adj_2025\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16980\,
            carryout => \foc.u_Park_Transform.n16981\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_6_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36099\,
            in2 => \N__35632\,
            in3 => \N__35614\,
            lcout => \foc.u_Park_Transform.n265_adj_2023\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16981\,
            carryout => \foc.u_Park_Transform.n16982\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_7_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35611\,
            in2 => \N__36127\,
            in3 => \N__35593\,
            lcout => \foc.u_Park_Transform.n314_adj_2010\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16982\,
            carryout => \foc.u_Park_Transform.n16983\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_8_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36103\,
            in2 => \N__35590\,
            in3 => \N__35572\,
            lcout => \foc.u_Park_Transform.n363_adj_1998\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16983\,
            carryout => \foc.u_Park_Transform.n16984\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_9_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35569\,
            in2 => \N__36128\,
            in3 => \N__36241\,
            lcout => \foc.u_Park_Transform.n412_adj_1995\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16984\,
            carryout => \foc.u_Park_Transform.n16985\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_10_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36107\,
            in2 => \N__36238\,
            in3 => \N__36220\,
            lcout => \foc.u_Park_Transform.n461_adj_2007\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \foc.u_Park_Transform.n16986\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_11_lut_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36217\,
            in2 => \N__36129\,
            in3 => \N__36199\,
            lcout => \foc.u_Park_Transform.n510\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16986\,
            carryout => \foc.u_Park_Transform.n16987\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_12_lut_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36111\,
            in2 => \N__36196\,
            in3 => \N__36178\,
            lcout => \foc.u_Park_Transform.n559\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16987\,
            carryout => \foc.u_Park_Transform.n16988\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_13_lut_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36175\,
            in2 => \N__36130\,
            in3 => \N__36160\,
            lcout => \foc.u_Park_Transform.n608_adj_2067\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16988\,
            carryout => \foc.u_Park_Transform.n16989\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_14_lut_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36157\,
            in2 => \N__36132\,
            in3 => \N__36142\,
            lcout => \foc.u_Park_Transform.n657_adj_2064\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16989\,
            carryout => \foc.u_Park_Transform.n16990\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_15_lut_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36139\,
            in2 => \N__36131\,
            in3 => \N__35944\,
            lcout => \foc.u_Park_Transform.n706_adj_2044\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16990\,
            carryout => \foc.u_Park_Transform.n16991\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_567_16_lut_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35941\,
            in2 => \N__35920\,
            in3 => \N__35899\,
            lcout => \foc.u_Park_Transform.n762_adj_2065\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n16991\,
            carryout => \foc.u_Park_Transform.n763_adj_2054\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n763_adj_2054_THRU_LUT4_0_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36490\,
            lcout => \foc.u_Park_Transform.n763_adj_2054_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_2_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36472\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2411\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36661\,
            in2 => \N__36400\,
            in3 => \N__36379\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2511\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36376\,
            in2 => \N__36678\,
            in3 => \N__36349\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2611\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_5_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36665\,
            in2 => \N__36346\,
            in3 => \N__36322\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2711\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_6_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36319\,
            in2 => \N__36679\,
            in3 => \N__36298\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2811\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_7_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36295\,
            in2 => \N__36681\,
            in3 => \N__36277\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2911\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_8_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36274\,
            in2 => \N__36680\,
            in3 => \N__36253\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3011\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_9_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36691\,
            in2 => \N__36682\,
            in3 => \N__36610\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3111\,
            ltout => OPEN,
            carryin => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17374\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_10_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36607\,
            in2 => \_gnd_net_\,
            in3 => \N__36589\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3215\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_LUT4_0_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36586\,
            lcout => \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i1_1_lut_2_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__36561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__44894\,
            in1 => \N__40458\,
            in2 => \_gnd_net_\,
            in3 => \N__40497\,
            lcout => n794,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66056\,
            in2 => \N__66217\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n81_adj_750\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17856\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66180\,
            in2 => \N__38416\,
            in3 => \N__36505\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n130_adj_748\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17856\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17857\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38407\,
            in2 => \N__66218\,
            in3 => \N__36493\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n179_adj_746\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17857\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17858\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66184\,
            in2 => \N__38398\,
            in3 => \N__36790\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n228_adj_742\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17858\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17859\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38386\,
            in2 => \N__66219\,
            in3 => \N__36775\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n277_adj_741\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17859\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17860\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66188\,
            in2 => \N__38536\,
            in3 => \N__36763\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n326\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17860\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17861\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38524\,
            in2 => \N__66220\,
            in3 => \N__36748\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n375\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17861\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17862\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66192\,
            in2 => \N__38515\,
            in3 => \N__36736\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n424\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17862\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17863\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38495\,
            in2 => \N__66293\,
            in3 => \N__36724\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n473\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17864\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66259\,
            in2 => \N__38502\,
            in3 => \N__36700\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n522\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17864\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17865\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45426\,
            in2 => \N__38503\,
            in3 => \N__36697\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n778_adj_737\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17865\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_LUT4_0_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36694\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_1_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43245\,
            in2 => \N__43249\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17957\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_2_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48968\,
            in2 => \_gnd_net_\,
            in3 => \N__36826\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17957\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17958\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_3_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43759\,
            in2 => \N__43222\,
            in3 => \N__36823\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17958\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17959\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_4_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43510\,
            in2 => \N__43741\,
            in3 => \N__36820\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17959\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17960\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_5_lut_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38794\,
            in2 => \N__43489\,
            in3 => \N__36817\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17960\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17961\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_6_lut_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38629\,
            in2 => \N__38776\,
            in3 => \N__36814\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17961\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17962\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_7_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41017\,
            in2 => \N__38614\,
            in3 => \N__36811\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17962\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17963\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_8_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41284\,
            in2 => \N__40999\,
            in3 => \N__36808\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17963\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17964\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_9_lut_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37009\,
            in2 => \N__41266\,
            in3 => \N__36805\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_22\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17965\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_10_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36994\,
            in2 => \N__36910\,
            in3 => \N__36898\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17965\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17966\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_11_lut_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36895\,
            in2 => \N__36889\,
            in3 => \N__36877\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17966\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17967\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_12_lut_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36874\,
            in2 => \N__36865\,
            in3 => \N__36856\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17967\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17968\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_13_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38479\,
            in2 => \N__36853\,
            in3 => \N__36841\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17968\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17969\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_14_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40651\,
            in2 => \N__38467\,
            in3 => \N__36838\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17969\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17970\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_15_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40633\,
            in2 => \N__40789\,
            in3 => \N__36835\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17970\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17971\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_16_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40774\,
            in2 => \N__40819\,
            in3 => \N__36832\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17971\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17972\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_17_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49011\,
            in2 => \_gnd_net_\,
            in3 => \N__36829\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66822\,
            in2 => \N__63111\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n72_adj_634\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36985\,
            in2 => \N__63132\,
            in3 => \N__36979\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n121_adj_633\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18092\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36976\,
            in2 => \N__63112\,
            in3 => \N__36970\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n170_adj_632\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18093\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36967\,
            in2 => \N__63133\,
            in3 => \N__36961\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n219_adj_631\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18094\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36958\,
            in2 => \N__63113\,
            in3 => \N__36952\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n268_adj_630\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18095\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36949\,
            in2 => \N__63134\,
            in3 => \N__36943\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n317_adj_629\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18096\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36940\,
            in2 => \N__63114\,
            in3 => \N__36934\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n366_adj_628\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18097\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36931\,
            in2 => \N__63135\,
            in3 => \N__36925\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n415_adj_627\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18098\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36922\,
            in2 => \N__63096\,
            in3 => \N__36913\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n464_adj_626\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63044\,
            in2 => \N__37072\,
            in3 => \N__37063\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n513_adj_625\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18100\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37060\,
            in2 => \N__63097\,
            in3 => \N__37054\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n562_adj_624\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18101\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18102\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63048\,
            in2 => \N__37051\,
            in3 => \N__37042\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n611_adj_623\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18102\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18103\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37039\,
            in2 => \N__63098\,
            in3 => \N__37033\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n660_adj_622\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18103\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63052\,
            in2 => \N__37030\,
            in3 => \N__37021\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n709_adj_621\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18104\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18105\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45169\,
            in2 => \N__37018\,
            in3 => \N__37000\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n766_adj_619\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18105\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_LUT4_0_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36997\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i9_1_lut_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37084\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i19_1_lut_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37336\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15_adj_518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i6_1_lut_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37120\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i26_1_lut_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37429\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i5_1_lut_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37129\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i8_1_lut_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37096\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i4_1_lut_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39151\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i7_1_lut_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37108\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i17_1_lut_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37141\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i14_1_lut_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37177\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i11_1_lut_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i16_1_lut_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37153\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i10_1_lut_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37216\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i13_1_lut_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i15_1_lut_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37165\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i12_1_lut_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37198\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_2_lut_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39139\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.dCurrent_4\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \foc.u_Park_Transform.n17277\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_3_lut_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39127\,
            in2 => \_gnd_net_\,
            in3 => \N__37111\,
            lcout => \foc.dCurrent_5\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17277\,
            carryout => \foc.u_Park_Transform.n17278\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_4_lut_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39115\,
            in2 => \_gnd_net_\,
            in3 => \N__37099\,
            lcout => \foc.dCurrent_6\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17278\,
            carryout => \foc.u_Park_Transform.n17279\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_5_lut_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39103\,
            in2 => \_gnd_net_\,
            in3 => \N__37087\,
            lcout => \foc.dCurrent_7\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17279\,
            carryout => \foc.u_Park_Transform.n17280\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_6_lut_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39091\,
            in2 => \_gnd_net_\,
            in3 => \N__37075\,
            lcout => \foc.dCurrent_8\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17280\,
            carryout => \foc.u_Park_Transform.n17281\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_7_lut_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39484\,
            in2 => \_gnd_net_\,
            in3 => \N__37210\,
            lcout => \foc.dCurrent_9\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17281\,
            carryout => \foc.u_Park_Transform.n17282\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_8_lut_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39472\,
            in2 => \_gnd_net_\,
            in3 => \N__37201\,
            lcout => \foc.dCurrent_10\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17282\,
            carryout => \foc.u_Park_Transform.n17283\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_9_lut_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39457\,
            in2 => \_gnd_net_\,
            in3 => \N__37192\,
            lcout => \foc.dCurrent_11\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17283\,
            carryout => \foc.u_Park_Transform.n17284\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_10_lut_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39442\,
            in2 => \_gnd_net_\,
            in3 => \N__37180\,
            lcout => \foc.dCurrent_12\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \foc.u_Park_Transform.n17285\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_11_lut_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39427\,
            in2 => \_gnd_net_\,
            in3 => \N__37168\,
            lcout => \foc.dCurrent_13\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17285\,
            carryout => \foc.u_Park_Transform.n17286\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_12_lut_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39415\,
            in2 => \_gnd_net_\,
            in3 => \N__37156\,
            lcout => \foc.dCurrent_14\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17286\,
            carryout => \foc.u_Park_Transform.n17287\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_13_lut_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39403\,
            in2 => \_gnd_net_\,
            in3 => \N__37144\,
            lcout => \foc.dCurrent_15\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17287\,
            carryout => \foc.u_Park_Transform.n17288\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_14_lut_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39211\,
            in2 => \_gnd_net_\,
            in3 => \N__37132\,
            lcout => \foc.dCurrent_16\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17288\,
            carryout => \foc.u_Park_Transform.n17289\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_15_lut_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37360\,
            in2 => \_gnd_net_\,
            in3 => \N__37345\,
            lcout => \foc.dCurrent_17\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17289\,
            carryout => \foc.u_Park_Transform.n17290\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_16_lut_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37342\,
            in2 => \_gnd_net_\,
            in3 => \N__37327\,
            lcout => \foc.dCurrent_18\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17290\,
            carryout => \foc.u_Park_Transform.n17291\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_17_lut_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37324\,
            in2 => \_gnd_net_\,
            in3 => \N__37309\,
            lcout => \foc.dCurrent_19\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17291\,
            carryout => \foc.u_Park_Transform.n17292\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_18_lut_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37306\,
            in2 => \_gnd_net_\,
            in3 => \N__37291\,
            lcout => \foc.dCurrent_20\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \foc.u_Park_Transform.n17293\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_19_lut_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37288\,
            in2 => \_gnd_net_\,
            in3 => \N__37273\,
            lcout => \foc.dCurrent_21\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17293\,
            carryout => \foc.u_Park_Transform.n17294\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_20_lut_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37270\,
            in2 => \_gnd_net_\,
            in3 => \N__37255\,
            lcout => \foc.dCurrent_22\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17294\,
            carryout => \foc.u_Park_Transform.n17295\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_21_lut_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37252\,
            in2 => \_gnd_net_\,
            in3 => \N__37237\,
            lcout => \foc.dCurrent_23\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17295\,
            carryout => \foc.u_Park_Transform.n17296\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_22_lut_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37234\,
            in2 => \_gnd_net_\,
            in3 => \N__37219\,
            lcout => \foc.dCurrent_24\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17296\,
            carryout => \foc.u_Park_Transform.n17297\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_23_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37435\,
            in2 => \_gnd_net_\,
            in3 => \N__37420\,
            lcout => \foc.dCurrent_25\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17297\,
            carryout => \foc.u_Park_Transform.n17298\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_24_lut_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37417\,
            in2 => \_gnd_net_\,
            in3 => \N__37411\,
            lcout => \foc.dCurrent_26\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17298\,
            carryout => \foc.u_Park_Transform.n17299\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_25_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37408\,
            in2 => \_gnd_net_\,
            in3 => \N__37402\,
            lcout => \foc.dCurrent_27\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17299\,
            carryout => \foc.u_Park_Transform.n17300\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_26_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37399\,
            in2 => \_gnd_net_\,
            in3 => \N__37393\,
            lcout => \foc.dCurrent_28\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \foc.u_Park_Transform.n17301\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_27_lut_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37390\,
            in2 => \_gnd_net_\,
            in3 => \N__37384\,
            lcout => \foc.dCurrent_29\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17301\,
            carryout => \foc.u_Park_Transform.n17302\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_28_lut_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37381\,
            in2 => \_gnd_net_\,
            in3 => \N__37375\,
            lcout => \foc.dCurrent_30\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17302\,
            carryout => \foc.u_Park_Transform.n17303\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.add_8094_29_lut_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37372\,
            in2 => \_gnd_net_\,
            in3 => \N__37366\,
            lcout => OPEN,
            ltout => \foc.dCurrent_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i32_1_lut_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37363\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i30_1_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n4_adj_515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i29_1_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37462\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i31_1_lut_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37456\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_2_lut_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42182\,
            in2 => \N__42700\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n57_adj_2116\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \foc.u_Park_Transform.n17221\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_3_lut_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42683\,
            in2 => \N__41542\,
            in3 => \N__37450\,
            lcout => \foc.u_Park_Transform.n106_adj_2115\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17221\,
            carryout => \foc.u_Park_Transform.n17222\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_4_lut_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42684\,
            in2 => \N__41521\,
            in3 => \N__37447\,
            lcout => \foc.u_Park_Transform.n155_adj_2114\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17222\,
            carryout => \foc.u_Park_Transform.n17223\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_5_lut_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41494\,
            in2 => \N__42701\,
            in3 => \N__37444\,
            lcout => \foc.u_Park_Transform.n204_adj_2113\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17223\,
            carryout => \foc.u_Park_Transform.n17224\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_6_lut_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42688\,
            in2 => \N__41473\,
            in3 => \N__37441\,
            lcout => \foc.u_Park_Transform.n253_adj_2112\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17224\,
            carryout => \foc.u_Park_Transform.n17225\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_7_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41446\,
            in2 => \N__42702\,
            in3 => \N__37438\,
            lcout => \foc.u_Park_Transform.n302_adj_2111\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17225\,
            carryout => \foc.u_Park_Transform.n17226\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_8_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42692\,
            in2 => \N__41422\,
            in3 => \N__37507\,
            lcout => \foc.u_Park_Transform.n351_adj_2108\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17226\,
            carryout => \foc.u_Park_Transform.n17227\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_9_lut_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41917\,
            in2 => \N__42703\,
            in3 => \N__37504\,
            lcout => \foc.u_Park_Transform.n400_adj_2106\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17227\,
            carryout => \foc.u_Park_Transform.n17228\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_10_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42666\,
            in2 => \N__41896\,
            in3 => \N__37501\,
            lcout => \foc.u_Park_Transform.n449_adj_2103\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \foc.u_Park_Transform.n17229\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_11_lut_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41863\,
            in2 => \N__42696\,
            in3 => \N__37498\,
            lcout => \foc.u_Park_Transform.n498_adj_2102\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17229\,
            carryout => \foc.u_Park_Transform.n17230\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_12_lut_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42670\,
            in2 => \N__41842\,
            in3 => \N__37495\,
            lcout => \foc.u_Park_Transform.n547_adj_2100\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17230\,
            carryout => \foc.u_Park_Transform.n17231\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_13_lut_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41815\,
            in2 => \N__42697\,
            in3 => \N__37492\,
            lcout => \foc.u_Park_Transform.n596_adj_2099\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17231\,
            carryout => \foc.u_Park_Transform.n17232\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_14_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41791\,
            in2 => \N__42699\,
            in3 => \N__37489\,
            lcout => \foc.u_Park_Transform.n645_adj_2098\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17232\,
            carryout => \foc.u_Park_Transform.n17233\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_15_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41770\,
            in2 => \N__42698\,
            in3 => \N__37486\,
            lcout => \foc.u_Park_Transform.n694_adj_2097\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17233\,
            carryout => \foc.u_Park_Transform.n17234\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_16_lut_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42789\,
            in2 => \N__41749\,
            in3 => \N__37471\,
            lcout => \foc.u_Park_Transform.n746\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17234\,
            carryout => \foc.u_Park_Transform.n747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n747_THRU_LUT4_0_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37780\,
            lcout => \foc.u_Park_Transform.n747_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_2_lut_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37749\,
            in2 => \N__41685\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n63\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \foc.u_Park_Transform.n17008\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_3_lut_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41638\,
            in2 => \N__37582\,
            in3 => \N__37573\,
            lcout => \foc.u_Park_Transform.n112\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17008\,
            carryout => \foc.u_Park_Transform.n17009\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_4_lut_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41639\,
            in2 => \N__37570\,
            in3 => \N__37561\,
            lcout => \foc.u_Park_Transform.n161\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17009\,
            carryout => \foc.u_Park_Transform.n17010\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_5_lut_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37558\,
            in2 => \N__41686\,
            in3 => \N__37552\,
            lcout => \foc.u_Park_Transform.n210\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17010\,
            carryout => \foc.u_Park_Transform.n17011\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_6_lut_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41643\,
            in2 => \N__37549\,
            in3 => \N__37540\,
            lcout => \foc.u_Park_Transform.n259\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17011\,
            carryout => \foc.u_Park_Transform.n17012\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_7_lut_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37537\,
            in2 => \N__41687\,
            in3 => \N__37531\,
            lcout => \foc.u_Park_Transform.n308\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17012\,
            carryout => \foc.u_Park_Transform.n17013\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_8_lut_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41647\,
            in2 => \N__37528\,
            in3 => \N__37519\,
            lcout => \foc.u_Park_Transform.n357\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17013\,
            carryout => \foc.u_Park_Transform.n17014\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_9_lut_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37516\,
            in2 => \N__41688\,
            in3 => \N__37510\,
            lcout => \foc.u_Park_Transform.n406\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17014\,
            carryout => \foc.u_Park_Transform.n17015\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_10_lut_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41692\,
            in2 => \N__37903\,
            in3 => \N__37894\,
            lcout => \foc.u_Park_Transform.n455\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \foc.u_Park_Transform.n17016\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_11_lut_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37891\,
            in2 => \N__41707\,
            in3 => \N__37885\,
            lcout => \foc.u_Park_Transform.n504\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17016\,
            carryout => \foc.u_Park_Transform.n17017\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_12_lut_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41696\,
            in2 => \N__37882\,
            in3 => \N__37873\,
            lcout => \foc.u_Park_Transform.n553\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17017\,
            carryout => \foc.u_Park_Transform.n17018\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_13_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37870\,
            in2 => \N__41708\,
            in3 => \N__37864\,
            lcout => \foc.u_Park_Transform.n602\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17018\,
            carryout => \foc.u_Park_Transform.n17019\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_14_lut_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41700\,
            in2 => \N__37861\,
            in3 => \N__37852\,
            lcout => \foc.u_Park_Transform.n651\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17019\,
            carryout => \foc.u_Park_Transform.n17020\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_15_lut_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37849\,
            in2 => \N__41709\,
            in3 => \N__37843\,
            lcout => \foc.u_Park_Transform.n700\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17020\,
            carryout => \foc.u_Park_Transform.n17021\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_565_16_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37840\,
            in2 => \N__37822\,
            in3 => \N__37801\,
            lcout => \foc.u_Park_Transform.n754\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17021\,
            carryout => \foc.u_Park_Transform.n755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n755_THRU_LUT4_0_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37798\,
            lcout => \foc.u_Park_Transform.n755_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_2_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40313\,
            in2 => \N__39313\,
            in3 => \_gnd_net_\,
            lcout => \foc.qCurrent_3\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \foc.u_Park_Transform.n17068\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_3_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39274\,
            in2 => \N__40090\,
            in3 => \N__37927\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_2\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17068\,
            carryout => \foc.u_Park_Transform.n17069\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40081\,
            in2 => \N__39314\,
            in3 => \N__37924\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_3\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17069\,
            carryout => \foc.u_Park_Transform.n17070\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_5_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39278\,
            in2 => \N__40072\,
            in3 => \N__37921\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_4\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17070\,
            carryout => \foc.u_Park_Transform.n17071\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_6_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40060\,
            in2 => \N__39315\,
            in3 => \N__37918\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_5\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17071\,
            carryout => \foc.u_Park_Transform.n17072\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_7_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39282\,
            in2 => \N__40051\,
            in3 => \N__37915\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_6\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17072\,
            carryout => \foc.u_Park_Transform.n17073\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_8_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40039\,
            in2 => \N__39316\,
            in3 => \N__37912\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_7\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17073\,
            carryout => \foc.u_Park_Transform.n17074\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_9_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39286\,
            in2 => \N__40030\,
            in3 => \N__37909\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_8\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17074\,
            carryout => \foc.u_Park_Transform.n17075\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_10_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40018\,
            in2 => \N__39348\,
            in3 => \N__37906\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_9\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \foc.u_Park_Transform.n17076\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_11_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40198\,
            in2 => \N__39351\,
            in3 => \N__38008\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_10\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17076\,
            carryout => \foc.u_Park_Transform.n17077\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_12_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40189\,
            in2 => \N__39349\,
            in3 => \N__38005\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_11\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17077\,
            carryout => \foc.u_Park_Transform.n17078\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_13_lut_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40180\,
            in2 => \N__39352\,
            in3 => \N__38002\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_12\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17078\,
            carryout => \foc.u_Park_Transform.n17079\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_14_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40171\,
            in2 => \N__39350\,
            in3 => \N__37999\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_13\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17079\,
            carryout => \foc.u_Park_Transform.n17080\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_15_lut_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40162\,
            in2 => \N__39353\,
            in3 => \N__37996\,
            lcout => \foc.u_Park_Transform.Product4_mul_temp_14\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17080\,
            carryout => \foc.u_Park_Transform.n17081\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_561_16_lut_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39195\,
            in2 => \N__40153\,
            in3 => \N__37972\,
            lcout => \foc.u_Park_Transform.n738_adj_2003\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17081\,
            carryout => \foc.u_Park_Transform.n739_adj_2006\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n739_adj_2006_THRU_LUT4_0_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37969\,
            lcout => \foc.u_Park_Transform.n739_adj_2006_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_2_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37951\,
            in2 => \N__44893\,
            in3 => \N__37942\,
            lcout => \foc.qCurrent_4\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \foc.u_Park_Transform.n15748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_3_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37939\,
            in2 => \N__68390\,
            in3 => \N__37930\,
            lcout => \foc.qCurrent_5\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15748\,
            carryout => \foc.u_Park_Transform.n15749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_4_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38107\,
            in2 => \N__68393\,
            in3 => \N__38098\,
            lcout => \foc.qCurrent_6\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15749\,
            carryout => \foc.u_Park_Transform.n15750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_5_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38095\,
            in2 => \N__68391\,
            in3 => \N__38086\,
            lcout => \foc.qCurrent_7\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15750\,
            carryout => \foc.u_Park_Transform.n15751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_6_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38083\,
            in2 => \N__68394\,
            in3 => \N__38074\,
            lcout => \foc.qCurrent_8\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15751\,
            carryout => \foc.u_Park_Transform.n15752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_7_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38071\,
            in2 => \N__68392\,
            in3 => \N__38062\,
            lcout => \foc.qCurrent_9\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15752\,
            carryout => \foc.u_Park_Transform.n15753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_8_lut_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38059\,
            in2 => \N__68395\,
            in3 => \N__38050\,
            lcout => \foc.qCurrent_10\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15753\,
            carryout => \foc.u_Park_Transform.n15754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_9_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68332\,
            in2 => \N__38047\,
            in3 => \N__38038\,
            lcout => \foc.qCurrent_11\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15754\,
            carryout => \foc.u_Park_Transform.n15755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_10_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38035\,
            in2 => \N__68396\,
            in3 => \N__38026\,
            lcout => \foc.qCurrent_12\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \foc.u_Park_Transform.n15756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_11_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68336\,
            in2 => \N__38023\,
            in3 => \N__38011\,
            lcout => \foc.qCurrent_13\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15756\,
            carryout => \foc.u_Park_Transform.n15757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_12_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38245\,
            in2 => \N__68397\,
            in3 => \N__38236\,
            lcout => \foc.qCurrent_14\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15757\,
            carryout => \foc.u_Park_Transform.n15758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_13_lut_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68340\,
            in2 => \N__38233\,
            in3 => \N__38221\,
            lcout => \foc.qCurrent_15\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15758\,
            carryout => \foc.u_Park_Transform.n15759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_14_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38218\,
            in2 => \N__68398\,
            in3 => \N__38209\,
            lcout => \foc.qCurrent_16\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15759\,
            carryout => \foc.u_Park_Transform.n15760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_15_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68344\,
            in2 => \N__38206\,
            in3 => \N__38191\,
            lcout => \foc.qCurrent_17\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15760\,
            carryout => \foc.u_Park_Transform.n15761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_16_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38188\,
            in2 => \N__68399\,
            in3 => \N__38176\,
            lcout => \foc.qCurrent_18\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15761\,
            carryout => \foc.u_Park_Transform.n15762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_17_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68348\,
            in2 => \N__38173\,
            in3 => \N__38158\,
            lcout => \foc.qCurrent_19\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15762\,
            carryout => \foc.u_Park_Transform.n15763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_18_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38155\,
            in2 => \N__68400\,
            in3 => \N__38143\,
            lcout => \foc.qCurrent_20\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \foc.u_Park_Transform.n15764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_19_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68352\,
            in2 => \N__38140\,
            in3 => \N__38125\,
            lcout => \foc.qCurrent_21\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15764\,
            carryout => \foc.u_Park_Transform.n15765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_20_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38122\,
            in2 => \N__68401\,
            in3 => \N__38110\,
            lcout => \foc.qCurrent_22\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15765\,
            carryout => \foc.u_Park_Transform.n15766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_21_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68356\,
            in2 => \N__38377\,
            in3 => \N__38362\,
            lcout => \foc.qCurrent_23\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15766\,
            carryout => \foc.u_Park_Transform.n15767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_22_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38359\,
            in2 => \N__68402\,
            in3 => \N__38347\,
            lcout => \foc.qCurrent_24\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15767\,
            carryout => \foc.u_Park_Transform.n15768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_23_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68360\,
            in2 => \N__38344\,
            in3 => \N__38329\,
            lcout => \foc.qCurrent_25\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15768\,
            carryout => \foc.u_Park_Transform.n15769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_24_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38326\,
            in2 => \N__68403\,
            in3 => \N__38314\,
            lcout => \foc.qCurrent_26\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15769\,
            carryout => \foc.u_Park_Transform.n15770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_25_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68364\,
            in2 => \N__38311\,
            in3 => \N__38296\,
            lcout => \foc.qCurrent_27\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15770\,
            carryout => \foc.u_Park_Transform.n15771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_26_lut_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38293\,
            in2 => \N__68426\,
            in3 => \N__38281\,
            lcout => \foc.qCurrent_28\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \foc.u_Park_Transform.n15772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_27_lut_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68407\,
            in2 => \N__38278\,
            in3 => \N__38263\,
            lcout => \foc.qCurrent_29\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15772\,
            carryout => \foc.u_Park_Transform.n15773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_28_lut_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38260\,
            in2 => \N__68427\,
            in3 => \N__38248\,
            lcout => \foc.qCurrent_30\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n15773\,
            carryout => \foc.u_Park_Transform.n15774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.sub_65_add_2_29_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38455\,
            in1 => \N__68411\,
            in2 => \_gnd_net_\,
            in3 => \N__38443\,
            lcout => \foc.qCurrent_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i20_1_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38440\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i28_1_lut_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i22_1_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38428\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i29_1_lut_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38422\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65739\,
            in2 => \N__66028\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n84_adj_749\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40723\,
            in2 => \N__66031\,
            in3 => \N__38401\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n133_adj_747\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17727\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17728\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40717\,
            in2 => \N__66029\,
            in3 => \N__38389\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n182_adj_745\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17728\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17729\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65975\,
            in2 => \N__40708\,
            in3 => \N__38380\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n231_adj_744\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17729\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17730\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40696\,
            in2 => \N__66030\,
            in3 => \N__38527\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n280_adj_743\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17730\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17731\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65979\,
            in2 => \N__40687\,
            in3 => \N__38518\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n329_adj_740\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17731\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17732\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65983\,
            in2 => \N__40674\,
            in3 => \N__38506\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n378_adj_739\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17732\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17733\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40670\,
            in2 => \N__66032\,
            in3 => \N__38482\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17733\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45399\,
            in2 => \N__40675\,
            in3 => \N__38473\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n782_adj_735\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_LUT4_0_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38470\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__48967\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63607\,
            in2 => \N__63889\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n63_adj_682\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18047\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40762\,
            in2 => \N__63893\,
            in3 => \N__38458\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n112_adj_681\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18047\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18048\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40756\,
            in2 => \N__63890\,
            in3 => \N__38563\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n161_adj_680\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18048\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18049\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40747\,
            in2 => \N__63894\,
            in3 => \N__38560\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n210_adj_679\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18049\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18050\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40738\,
            in2 => \N__63891\,
            in3 => \N__38557\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n259_adj_678\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18050\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18051\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40900\,
            in2 => \N__63895\,
            in3 => \N__38554\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n308_adj_677\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18051\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18052\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40891\,
            in2 => \N__63892\,
            in3 => \N__38551\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n357_adj_676\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18052\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18053\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40882\,
            in2 => \N__63896\,
            in3 => \N__38548\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n406_adj_675\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18053\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18054\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40873\,
            in2 => \N__63946\,
            in3 => \N__38545\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n455_adj_674\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18055\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40864\,
            in2 => \N__63949\,
            in3 => \N__38542\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n504_adj_673\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18055\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18056\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40855\,
            in2 => \N__63947\,
            in3 => \N__38539\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n553_adj_672\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18056\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18057\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40846\,
            in2 => \N__63950\,
            in3 => \N__38638\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n602_adj_671\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18057\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18058\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40837\,
            in2 => \N__63948\,
            in3 => \N__38635\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n651_adj_670\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18058\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18059\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41038\,
            in2 => \N__63951\,
            in3 => \N__38632\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n700_adj_669\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18059\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18060\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45241\,
            in2 => \N__41029\,
            in3 => \N__38620\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n754_adj_667\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18060\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_LUT4_0_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38617\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63875\,
            in2 => \N__64237\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n60_adj_698\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18032\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64207\,
            in2 => \N__38602\,
            in3 => \N__38590\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n109_adj_697\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18032\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18033\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38587\,
            in2 => \N__64238\,
            in3 => \N__38578\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n158_adj_696\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18033\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18034\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64211\,
            in2 => \N__38575\,
            in3 => \N__38749\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n207_adj_695\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18034\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18035\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38746\,
            in2 => \N__64239\,
            in3 => \N__38737\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n256_adj_694\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18035\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18036\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64215\,
            in2 => \N__38734\,
            in3 => \N__38722\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n305_adj_693\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18036\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18037\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38719\,
            in2 => \N__64240\,
            in3 => \N__38710\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n354_adj_692\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18037\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18038\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64219\,
            in2 => \N__38707\,
            in3 => \N__38695\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n403_adj_691\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18038\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18039\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38692\,
            in2 => \N__64233\,
            in3 => \N__38683\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n452_adj_690\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18040\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64192\,
            in2 => \N__38680\,
            in3 => \N__38668\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n501_adj_689\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18040\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18041\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38665\,
            in2 => \N__64234\,
            in3 => \N__38656\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n550_adj_688\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18041\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18042\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64196\,
            in2 => \N__38653\,
            in3 => \N__38641\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n599_adj_687\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18042\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18043\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38833\,
            in2 => \N__64235\,
            in3 => \N__38824\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n648_adj_686\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18043\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18044\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64200\,
            in2 => \N__38821\,
            in3 => \N__38809\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n697_adj_685\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18044\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18045\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45268\,
            in2 => \N__38806\,
            in3 => \N__38782\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n750_adj_683\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18045\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_LUT4_0_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38779\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_2_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68435\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_3_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42856\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15775\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_4_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38761\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15776\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_5_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38755\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15777\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_6_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38887\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15778\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_7_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38881\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15779\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_8_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38875\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15780\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_9_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38869\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15781\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_10_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38863\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_11_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38857\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15783\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_12_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38851\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15784\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_13_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38845\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15785\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_14_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38839\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15786\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_15_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38980\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15787\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_16_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38974\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15788\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_17_lut_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38968\,
            in2 => \_gnd_net_\,
            in3 => \N__38962\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15789\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_18_lut_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38959\,
            in2 => \_gnd_net_\,
            in3 => \N__38947\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_19_lut_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38944\,
            in2 => \_gnd_net_\,
            in3 => \N__38935\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15791\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_20_lut_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38932\,
            in2 => \_gnd_net_\,
            in3 => \N__38920\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15792\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_21_lut_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38917\,
            in2 => \_gnd_net_\,
            in3 => \N__38905\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15793\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_22_lut_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38902\,
            in2 => \_gnd_net_\,
            in3 => \N__38890\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15794\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_23_lut_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39079\,
            in2 => \_gnd_net_\,
            in3 => \N__39067\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_22\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15795\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_24_lut_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39064\,
            in2 => \_gnd_net_\,
            in3 => \N__39052\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15796\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_25_lut_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39049\,
            in2 => \_gnd_net_\,
            in3 => \N__39037\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15797\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_26_lut_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39034\,
            in2 => \_gnd_net_\,
            in3 => \N__39025\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_25\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_27_lut_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39157\,
            in2 => \_gnd_net_\,
            in3 => \N__39022\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15799\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_28_lut_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41722\,
            in2 => \_gnd_net_\,
            in3 => \N__39019\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15800\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_29_lut_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39016\,
            in2 => \_gnd_net_\,
            in3 => \N__39007\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15801\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_30_lut_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39004\,
            in2 => \_gnd_net_\,
            in3 => \N__38995\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15802\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_31_lut_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38992\,
            in2 => \_gnd_net_\,
            in3 => \N__38983\,
            lcout => \Error_sub_temp_30\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15803\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_32_lut_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__39175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39166\,
            lcout => \Error_sub_temp_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i27_1_lut_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39163\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_2_lut_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40390\,
            in2 => \N__39387\,
            in3 => \_gnd_net_\,
            lcout => \foc.dCurrent_3\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \foc.u_Park_Transform.n17251\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_3_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39607\,
            in2 => \N__39391\,
            in3 => \N__39130\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_2\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17251\,
            carryout => \foc.u_Park_Transform.n17252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_4_lut_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39589\,
            in2 => \N__39388\,
            in3 => \N__39118\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_3\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17252\,
            carryout => \foc.u_Park_Transform.n17253\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_5_lut_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39372\,
            in2 => \N__39568\,
            in3 => \N__39106\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_4\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17253\,
            carryout => \foc.u_Park_Transform.n17254\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_6_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39547\,
            in2 => \N__39389\,
            in3 => \N__39094\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_5\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17254\,
            carryout => \foc.u_Park_Transform.n17255\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_7_lut_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39376\,
            in2 => \N__39526\,
            in3 => \N__39082\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_6\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17255\,
            carryout => \foc.u_Park_Transform.n17256\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_8_lut_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39505\,
            in2 => \N__39390\,
            in3 => \N__39475\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_7\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17256\,
            carryout => \foc.u_Park_Transform.n17257\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_9_lut_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39380\,
            in2 => \N__39808\,
            in3 => \N__39460\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_8\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17257\,
            carryout => \foc.u_Park_Transform.n17258\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_10_lut_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39787\,
            in2 => \N__39384\,
            in3 => \N__39445\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_9\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \foc.u_Park_Transform.n17259\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_11_lut_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39357\,
            in2 => \N__39769\,
            in3 => \N__39430\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_10\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17259\,
            carryout => \foc.u_Park_Transform.n17260\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_12_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39748\,
            in2 => \N__39385\,
            in3 => \N__39418\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_11\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17260\,
            carryout => \foc.u_Park_Transform.n17261\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_13_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39361\,
            in2 => \N__39727\,
            in3 => \N__39406\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_12\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17261\,
            carryout => \foc.u_Park_Transform.n17262\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_14_lut_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39706\,
            in2 => \N__39386\,
            in3 => \N__39394\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_13\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17262\,
            carryout => \foc.u_Park_Transform.n17263\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_15_lut_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39365\,
            in2 => \N__39685\,
            in3 => \N__39202\,
            lcout => \foc.u_Park_Transform.Product1_mul_temp_14\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17263\,
            carryout => \foc.u_Park_Transform.n17264\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_16_lut_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39199\,
            in2 => \N__39664\,
            in3 => \N__39628\,
            lcout => \foc.u_Park_Transform.n738\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17264\,
            carryout => \foc.u_Park_Transform.n739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n739_THRU_LUT4_0_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39625\,
            lcout => \foc.u_Park_Transform.n739_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_2_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42633\,
            in2 => \N__40386\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n54_adj_2095\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \foc.u_Park_Transform.n17236\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_3_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40367\,
            in2 => \N__39598\,
            in3 => \N__39580\,
            lcout => \foc.u_Park_Transform.n103_adj_2092\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17236\,
            carryout => \foc.u_Park_Transform.n17237\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_4_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40368\,
            in2 => \N__39577\,
            in3 => \N__39556\,
            lcout => \foc.u_Park_Transform.n152_adj_2088\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17237\,
            carryout => \foc.u_Park_Transform.n17238\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_5_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39553\,
            in2 => \N__40387\,
            in3 => \N__39538\,
            lcout => \foc.u_Park_Transform.n201_adj_2085\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17238\,
            carryout => \foc.u_Park_Transform.n17239\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_6_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40372\,
            in2 => \N__39535\,
            in3 => \N__39514\,
            lcout => \foc.u_Park_Transform.n250_adj_2084\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17239\,
            carryout => \foc.u_Park_Transform.n17240\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_7_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39511\,
            in2 => \N__40388\,
            in3 => \N__39496\,
            lcout => \foc.u_Park_Transform.n299_adj_2083\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17240\,
            carryout => \foc.u_Park_Transform.n17241\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_8_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40376\,
            in2 => \N__39493\,
            in3 => \N__39796\,
            lcout => \foc.u_Park_Transform.n348_adj_2082\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17241\,
            carryout => \foc.u_Park_Transform.n17242\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_9_lut_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39793\,
            in2 => \N__40389\,
            in3 => \N__39781\,
            lcout => \foc.u_Park_Transform.n397_adj_2081\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17242\,
            carryout => \foc.u_Park_Transform.n17243\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_10_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40352\,
            in2 => \N__39778\,
            in3 => \N__39757\,
            lcout => \foc.u_Park_Transform.n446_adj_2079\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \foc.u_Park_Transform.n17244\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_11_lut_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39754\,
            in2 => \N__40383\,
            in3 => \N__39739\,
            lcout => \foc.u_Park_Transform.n495_adj_2077\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17244\,
            carryout => \foc.u_Park_Transform.n17245\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_12_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40356\,
            in2 => \N__39736\,
            in3 => \N__39715\,
            lcout => \foc.u_Park_Transform.n544_adj_2074\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17245\,
            carryout => \foc.u_Park_Transform.n17246\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_13_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39712\,
            in2 => \N__40384\,
            in3 => \N__39697\,
            lcout => \foc.u_Park_Transform.n593_adj_2073\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17246\,
            carryout => \foc.u_Park_Transform.n17247\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_14_lut_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40360\,
            in2 => \N__39694\,
            in3 => \N__39673\,
            lcout => \foc.u_Park_Transform.n642_adj_2072\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17247\,
            carryout => \foc.u_Park_Transform.n17248\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_15_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39670\,
            in2 => \N__40385\,
            in3 => \N__39652\,
            lcout => \foc.u_Park_Transform.n691_adj_2071\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17248\,
            carryout => \foc.u_Park_Transform.n17249\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_16_lut_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40516\,
            in2 => \N__39916\,
            in3 => \N__39895\,
            lcout => \foc.u_Park_Transform.n742\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17249\,
            carryout => \foc.u_Park_Transform.n743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n743_THRU_LUT4_0_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39892\,
            lcout => \foc.u_Park_Transform.n743_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_2_lut_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42091\,
            in2 => \N__41689\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n60\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \foc.u_Park_Transform.n17023\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_3_lut_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39874\,
            in2 => \N__42134\,
            in3 => \N__39868\,
            lcout => \foc.u_Park_Transform.n109\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17023\,
            carryout => \foc.u_Park_Transform.n17024\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_4_lut_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42095\,
            in2 => \N__39865\,
            in3 => \N__39856\,
            lcout => \foc.u_Park_Transform.n158\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17024\,
            carryout => \foc.u_Park_Transform.n17025\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_5_lut_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39853\,
            in2 => \N__42135\,
            in3 => \N__39847\,
            lcout => \foc.u_Park_Transform.n207\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17025\,
            carryout => \foc.u_Park_Transform.n17026\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_6_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42099\,
            in2 => \N__39844\,
            in3 => \N__39835\,
            lcout => \foc.u_Park_Transform.n256\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17026\,
            carryout => \foc.u_Park_Transform.n17027\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_7_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39832\,
            in2 => \N__42136\,
            in3 => \N__39826\,
            lcout => \foc.u_Park_Transform.n305\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17027\,
            carryout => \foc.u_Park_Transform.n17028\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_8_lut_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42103\,
            in2 => \N__39823\,
            in3 => \N__39811\,
            lcout => \foc.u_Park_Transform.n354\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17028\,
            carryout => \foc.u_Park_Transform.n17029\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_9_lut_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40012\,
            in2 => \N__42137\,
            in3 => \N__40006\,
            lcout => \foc.u_Park_Transform.n403\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17029\,
            carryout => \foc.u_Park_Transform.n17030\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_10_lut_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42138\,
            in2 => \N__40003\,
            in3 => \N__39994\,
            lcout => \foc.u_Park_Transform.n452\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \foc.u_Park_Transform.n17031\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_11_lut_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39991\,
            in2 => \N__42183\,
            in3 => \N__39985\,
            lcout => \foc.u_Park_Transform.n501\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17031\,
            carryout => \foc.u_Park_Transform.n17032\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_12_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42142\,
            in2 => \N__39982\,
            in3 => \N__39973\,
            lcout => \foc.u_Park_Transform.n550\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17032\,
            carryout => \foc.u_Park_Transform.n17033\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_13_lut_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39970\,
            in2 => \N__42184\,
            in3 => \N__39964\,
            lcout => \foc.u_Park_Transform.n599\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17033\,
            carryout => \foc.u_Park_Transform.n17034\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_14_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42146\,
            in2 => \N__39961\,
            in3 => \N__39952\,
            lcout => \foc.u_Park_Transform.n648\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17034\,
            carryout => \foc.u_Park_Transform.n17035\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_15_lut_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39949\,
            in2 => \N__42185\,
            in3 => \N__39943\,
            lcout => \foc.u_Park_Transform.n697\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17035\,
            carryout => \foc.u_Park_Transform.n17036\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_564_16_lut_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42291\,
            in2 => \N__39940\,
            in3 => \N__39919\,
            lcout => \foc.u_Park_Transform.n750_adj_2117\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17036\,
            carryout => \foc.u_Park_Transform.n751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n751_THRU_LUT4_0_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40108\,
            lcout => \foc.u_Park_Transform.n751_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_2_lut_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40303\,
            in2 => \N__42593\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n54\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \foc.u_Park_Transform.n17053\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_3_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42040\,
            in2 => \N__40350\,
            in3 => \N__40075\,
            lcout => \foc.u_Park_Transform.n103\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17053\,
            carryout => \foc.u_Park_Transform.n17054\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_4_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40307\,
            in2 => \N__42025\,
            in3 => \N__40063\,
            lcout => \foc.u_Park_Transform.n152\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17054\,
            carryout => \foc.u_Park_Transform.n17055\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_5_lut_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41998\,
            in2 => \N__40351\,
            in3 => \N__40054\,
            lcout => \foc.u_Park_Transform.n201\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17055\,
            carryout => \foc.u_Park_Transform.n17056\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_6_lut_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40311\,
            in2 => \N__41980\,
            in3 => \N__40042\,
            lcout => \foc.u_Park_Transform.n250\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17056\,
            carryout => \foc.u_Park_Transform.n17057\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_7_lut_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40348\,
            in2 => \N__41956\,
            in3 => \N__40033\,
            lcout => \foc.u_Park_Transform.n299\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17057\,
            carryout => \foc.u_Park_Transform.n17058\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_8_lut_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40312\,
            in2 => \N__41935\,
            in3 => \N__40021\,
            lcout => \foc.u_Park_Transform.n348\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17058\,
            carryout => \foc.u_Park_Transform.n17059\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_9_lut_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40349\,
            in2 => \N__42469\,
            in3 => \N__40201\,
            lcout => \foc.u_Park_Transform.n397\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17059\,
            carryout => \foc.u_Park_Transform.n17060\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_10_lut_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40261\,
            in2 => \N__42448\,
            in3 => \N__40192\,
            lcout => \foc.u_Park_Transform.n446\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \foc.u_Park_Transform.n17061\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_11_lut_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42421\,
            in2 => \N__40301\,
            in3 => \N__40183\,
            lcout => \foc.u_Park_Transform.n495\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17061\,
            carryout => \foc.u_Park_Transform.n17062\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_12_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40265\,
            in2 => \N__42403\,
            in3 => \N__40174\,
            lcout => \foc.u_Park_Transform.n544\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17062\,
            carryout => \foc.u_Park_Transform.n17063\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_13_lut_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42376\,
            in2 => \N__40302\,
            in3 => \N__40165\,
            lcout => \foc.u_Park_Transform.n593\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17063\,
            carryout => \foc.u_Park_Transform.n17064\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_14_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40269\,
            in2 => \N__42358\,
            in3 => \N__40156\,
            lcout => \foc.u_Park_Transform.n642\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17064\,
            carryout => \foc.u_Park_Transform.n17065\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_15_lut_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40270\,
            in2 => \N__42334\,
            in3 => \N__40144\,
            lcout => \foc.u_Park_Transform.n691\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17065\,
            carryout => \foc.u_Park_Transform.n17066\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_562_16_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40512\,
            in2 => \N__42313\,
            in3 => \N__40129\,
            lcout => \foc.u_Park_Transform.n742_adj_2086\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17066\,
            carryout => \foc.u_Park_Transform.n743_adj_2096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n743_adj_2096_THRU_LUT4_0_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40126\,
            lcout => \foc.u_Park_Transform.n743_adj_2096_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i5_1_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n27_adj_753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_i501_2_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40405\,
            lcout => \foc.u_Park_Transform.n741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__40501\,
            in1 => \N__40457\,
            in2 => \_gnd_net_\,
            in3 => \N__44912\,
            lcout => n142,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i7_1_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40411\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i4_2_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40404\,
            lcout => \foc.u_Park_Transform.n592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i2_1_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40228\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i17_1_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40219\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i18_1_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i12_1_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i15_1_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40576\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i13_1_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40570\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i3_1_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40564\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i10_1_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40558\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i14_1_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i21_1_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40546\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i16_1_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40540\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i23_1_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40534\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i26_1_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i25_1_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40621\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i11_1_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40615\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_adj_752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_272_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011100000"
        )
    port map (
            in0 => \N__65508\,
            in1 => \N__44687\,
            in2 => \N__44832\,
            in3 => \N__44668\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i27_1_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i19_1_lut_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40603\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_271_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011000000"
        )
    port map (
            in0 => \N__44667\,
            in1 => \N__65507\,
            in2 => \N__44689\,
            in3 => \N__44823\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_757_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__65510\,
            in1 => \N__44688\,
            in2 => \N__40597\,
            in3 => \N__44828\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19841_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_273_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011000000"
        )
    port map (
            in0 => \N__40594\,
            in1 => \N__65509\,
            in2 => \N__40585\,
            in3 => \N__44827\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n26_adj_759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i30_1_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i24_1_lut_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40729\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65467\,
            in2 => \N__65734\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n87_adj_730\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17973\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40828\,
            in2 => \N__65737\,
            in3 => \N__40711\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n136_adj_728\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17973\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17974\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44779\,
            in2 => \N__65735\,
            in3 => \N__40699\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n185_adj_726\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17974\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17975\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43048\,
            in2 => \N__65738\,
            in3 => \N__40690\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n234_adj_724\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17975\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17976\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43034\,
            in2 => \N__65736\,
            in3 => \N__40678\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n283_adj_723\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17976\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17977\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65697\,
            in2 => \N__43041\,
            in3 => \N__40654\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17977\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17978\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45375\,
            in2 => \N__43042\,
            in3 => \N__40639\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n786_adj_719\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17978\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_LUT4_0_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40636\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i12078_3_lut_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__45049\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45124\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n90_adj_729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_291_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001000"
        )
    port map (
            in0 => \N__40802\,
            in1 => \N__65118\,
            in2 => \_gnd_net_\,
            in3 => \N__65284\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n7_adj_760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_274_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__45125\,
            in1 => \N__40803\,
            in2 => \N__40822\,
            in3 => \N__65511\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_adj_732\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_4_lut_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010110100"
        )
    port map (
            in0 => \N__40804\,
            in1 => \N__44833\,
            in2 => \_gnd_net_\,
            in3 => \N__45126\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n790_adj_733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12680_3_lut_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__45050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65119\,
            lcout => n794_adj_2425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63180\,
            in2 => \N__63632\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n66_adj_666\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18062\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63587\,
            in2 => \N__40984\,
            in3 => \N__40750\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n115_adj_665\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18062\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18063\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40960\,
            in2 => \N__63633\,
            in3 => \N__40741\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n164_adj_664\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18063\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18064\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63591\,
            in2 => \N__40939\,
            in3 => \N__40732\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n213_adj_663\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18064\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18065\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40912\,
            in2 => \N__63634\,
            in3 => \N__40894\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n262_adj_662\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18065\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18066\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63595\,
            in2 => \N__41221\,
            in3 => \N__40885\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n311_adj_661\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18066\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18067\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41194\,
            in2 => \N__63635\,
            in3 => \N__40876\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n360_adj_660\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18067\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18068\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63599\,
            in2 => \N__41170\,
            in3 => \N__40867\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n409_adj_659\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18068\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18069\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41146\,
            in2 => \N__63622\,
            in3 => \N__40858\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n458_adj_658\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18070\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63561\,
            in2 => \N__41125\,
            in3 => \N__40849\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n507_adj_657\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18070\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18071\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41098\,
            in2 => \N__63623\,
            in3 => \N__40840\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n556_adj_656\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18071\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18072\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63565\,
            in2 => \N__41077\,
            in3 => \N__40831\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n605_adj_655\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18072\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18073\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41050\,
            in2 => \N__63624\,
            in3 => \N__41032\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n654_adj_654\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18073\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18074\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41335\,
            in2 => \N__63625\,
            in3 => \N__41020\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n703_adj_653\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18074\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18075\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45217\,
            in2 => \N__41311\,
            in3 => \N__41005\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n758_adj_651\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18075\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_LUT4_0_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41002\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62999\,
            in2 => \N__63284\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n69_adj_650\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18077\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63229\,
            in2 => \N__40972\,
            in3 => \N__40951\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n118_adj_649\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18077\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18078\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40948\,
            in2 => \N__63285\,
            in3 => \N__40927\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n167_adj_648\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18078\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18079\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63233\,
            in2 => \N__40924\,
            in3 => \N__40903\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n216_adj_647\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18079\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18080\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41230\,
            in2 => \N__63286\,
            in3 => \N__41209\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n265_adj_646\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18080\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18081\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63237\,
            in2 => \N__41206\,
            in3 => \N__41185\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n314_adj_645\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18081\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18082\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63280\,
            in2 => \N__41182\,
            in3 => \N__41158\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n363_adj_644\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18082\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18083\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41155\,
            in2 => \N__63336\,
            in3 => \N__41140\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n412_adj_643\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18083\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18084\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41137\,
            in2 => \N__63358\,
            in3 => \N__41113\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n461_adj_642\,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18085\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63311\,
            in2 => \N__41110\,
            in3 => \N__41089\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n510_adj_641\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18085\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18086\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41086\,
            in2 => \N__63359\,
            in3 => \N__41065\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n559_adj_640\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18086\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18087\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63315\,
            in2 => \N__41062\,
            in3 => \N__41041\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n608_adj_639\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18087\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18088\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41344\,
            in2 => \N__63360\,
            in3 => \N__41326\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n657_adj_638\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18088\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18089\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63319\,
            in2 => \N__41323\,
            in3 => \N__41299\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n706_adj_637\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18089\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18090\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45193\,
            in2 => \N__41296\,
            in3 => \N__41272\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n762_adj_635\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18090\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_LUT4_0_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41269\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__41241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41391\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__41251\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41250\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41242\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41380\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__41367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i11954_3_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__50342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44114\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__41392\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41379\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50343\,
            lcout => n141,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__41356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__41371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__41355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_128_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__44115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i28_1_lut_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41734\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_2_lut_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41710\,
            in2 => \N__42215\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n60_adj_2140\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \foc.u_Park_Transform.n17206\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_3_lut_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41530\,
            in2 => \N__42220\,
            in3 => \N__41509\,
            lcout => \foc.u_Park_Transform.n109_adj_2139\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17206\,
            carryout => \foc.u_Park_Transform.n17207\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_4_lut_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42203\,
            in2 => \N__41506\,
            in3 => \N__41485\,
            lcout => \foc.u_Park_Transform.n158_adj_2137\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17207\,
            carryout => \foc.u_Park_Transform.n17208\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_5_lut_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41482\,
            in2 => \N__42221\,
            in3 => \N__41461\,
            lcout => \foc.u_Park_Transform.n207_adj_2136\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17208\,
            carryout => \foc.u_Park_Transform.n17209\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_6_lut_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42207\,
            in2 => \N__41458\,
            in3 => \N__41434\,
            lcout => \foc.u_Park_Transform.n256_adj_2135\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17209\,
            carryout => \foc.u_Park_Transform.n17210\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_7_lut_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41431\,
            in2 => \N__42222\,
            in3 => \N__41407\,
            lcout => \foc.u_Park_Transform.n305_adj_2134\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17210\,
            carryout => \foc.u_Park_Transform.n17211\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_8_lut_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42211\,
            in2 => \N__41404\,
            in3 => \N__41908\,
            lcout => \foc.u_Park_Transform.n354_adj_2133\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17211\,
            carryout => \foc.u_Park_Transform.n17212\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_9_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41905\,
            in2 => \N__42223\,
            in3 => \N__41881\,
            lcout => \foc.u_Park_Transform.n403_adj_2132\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17212\,
            carryout => \foc.u_Park_Transform.n17213\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_10_lut_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42186\,
            in2 => \N__41878\,
            in3 => \N__41854\,
            lcout => \foc.u_Park_Transform.n452_adj_2131\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \foc.u_Park_Transform.n17214\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_11_lut_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41851\,
            in2 => \N__42216\,
            in3 => \N__41830\,
            lcout => \foc.u_Park_Transform.n501_adj_2130\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17214\,
            carryout => \foc.u_Park_Transform.n17215\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_12_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42190\,
            in2 => \N__41827\,
            in3 => \N__41803\,
            lcout => \foc.u_Park_Transform.n550_adj_2129\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17215\,
            carryout => \foc.u_Park_Transform.n17216\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_13_lut_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41800\,
            in2 => \N__42217\,
            in3 => \N__41782\,
            lcout => \foc.u_Park_Transform.n599_adj_2128\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17216\,
            carryout => \foc.u_Park_Transform.n17217\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_14_lut_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41779\,
            in2 => \N__42219\,
            in3 => \N__41761\,
            lcout => \foc.u_Park_Transform.n648_adj_2124\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17217\,
            carryout => \foc.u_Park_Transform.n17218\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_15_lut_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41758\,
            in2 => \N__42218\,
            in3 => \N__41737\,
            lcout => \foc.u_Park_Transform.n697_adj_2121\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17218\,
            carryout => \foc.u_Park_Transform.n17219\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_16_lut_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42295\,
            in2 => \N__42268\,
            in3 => \N__42244\,
            lcout => \foc.u_Park_Transform.n750\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17219\,
            carryout => \foc.u_Park_Transform.n751_adj_2142\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n751_adj_2142_THRU_LUT4_0_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42241\,
            lcout => \foc.u_Park_Transform.n751_adj_2142_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_2_lut_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42130\,
            in2 => \N__42628\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_Park_Transform.n57\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \foc.u_Park_Transform.n17038\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_3_lut_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42031\,
            in2 => \N__42629\,
            in3 => \N__42010\,
            lcout => \foc.u_Park_Transform.n106\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17038\,
            carryout => \foc.u_Park_Transform.n17039\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_4_lut_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42603\,
            in2 => \N__42007\,
            in3 => \N__41989\,
            lcout => \foc.u_Park_Transform.n155\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17039\,
            carryout => \foc.u_Park_Transform.n17040\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_5_lut_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41986\,
            in2 => \N__42630\,
            in3 => \N__41968\,
            lcout => \foc.u_Park_Transform.n204\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17040\,
            carryout => \foc.u_Park_Transform.n17041\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_6_lut_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42607\,
            in2 => \N__41965\,
            in3 => \N__41944\,
            lcout => \foc.u_Park_Transform.n253\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17041\,
            carryout => \foc.u_Park_Transform.n17042\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_7_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41941\,
            in2 => \N__42631\,
            in3 => \N__41920\,
            lcout => \foc.u_Park_Transform.n302\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17042\,
            carryout => \foc.u_Park_Transform.n17043\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_8_lut_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42611\,
            in2 => \N__42478\,
            in3 => \N__42457\,
            lcout => \foc.u_Park_Transform.n351\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17043\,
            carryout => \foc.u_Park_Transform.n17044\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_9_lut_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42454\,
            in2 => \N__42632\,
            in3 => \N__42433\,
            lcout => \foc.u_Park_Transform.n400\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17044\,
            carryout => \foc.u_Park_Transform.n17045\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_10_lut_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42555\,
            in2 => \N__42430\,
            in3 => \N__42412\,
            lcout => \foc.u_Park_Transform.n449\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \foc.u_Park_Transform.n17046\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_11_lut_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42409\,
            in2 => \N__42594\,
            in3 => \N__42388\,
            lcout => \foc.u_Park_Transform.n498\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17046\,
            carryout => \foc.u_Park_Transform.n17047\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_12_lut_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42559\,
            in2 => \N__42385\,
            in3 => \N__42367\,
            lcout => \foc.u_Park_Transform.n547\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17047\,
            carryout => \foc.u_Park_Transform.n17048\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_13_lut_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42364\,
            in2 => \N__42595\,
            in3 => \N__42346\,
            lcout => \foc.u_Park_Transform.n596\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17048\,
            carryout => \foc.u_Park_Transform.n17049\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_14_lut_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42563\,
            in2 => \N__42343\,
            in3 => \N__42322\,
            lcout => \foc.u_Park_Transform.n645\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17049\,
            carryout => \foc.u_Park_Transform.n17050\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_15_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42319\,
            in2 => \N__42596\,
            in3 => \N__42298\,
            lcout => \foc.u_Park_Transform.n694\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17050\,
            carryout => \foc.u_Park_Transform.n17051\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Beta_15__I_0_add_563_16_lut_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42796\,
            in2 => \N__42772\,
            in3 => \N__42751\,
            lcout => \foc.u_Park_Transform.n746_adj_2011\,
            ltout => OPEN,
            carryin => \foc.u_Park_Transform.n17051\,
            carryout => \foc.u_Park_Transform.n747_adj_2012\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.n747_adj_2012_THRU_LUT4_0_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42748\,
            lcout => \foc.u_Park_Transform.n747_adj_2012_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_3_lut_3_lut_4_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__44292\,
            in1 => \N__44436\,
            in2 => \_gnd_net_\,
            in3 => \N__42517\,
            lcout => OPEN,
            ltout => \foc.u_Park_Transform.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_3_lut_4_lut_adj_308_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44339\,
            in2 => \N__42727\,
            in3 => \N__44435\,
            lcout => \foc.u_Park_Transform.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i6_2_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42724\,
            lcout => \foc.u_Park_Transform.n595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_2_lut_4_lut_4_lut_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010001000"
        )
    port map (
            in0 => \N__42516\,
            in1 => \N__44291\,
            in2 => \_gnd_net_\,
            in3 => \N__44434\,
            lcout => \foc.u_Park_Transform.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i9_1_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42496\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i6_1_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42487\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i4_1_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42880\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i8_1_lut_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42871\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_2_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42862\,
            in2 => \N__42849\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15720\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_3_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42826\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15720\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15721\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_4_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42820\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15721\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15722\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_5_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42814\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15722\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15723\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_6_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42808\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15723\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15724\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_7_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42802\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15724\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15725\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_8_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42940\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15725\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15726\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_9_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42934\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15726\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_10_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42928\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15728\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_11_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42922\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15728\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15729\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_12_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42916\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15729\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15730\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_13_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42910\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15730\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15731\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_14_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42904\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15731\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15732\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_15_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42898\,
            in2 => \_gnd_net_\,
            in3 => \N__42892\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15732\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15733\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_16_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42889\,
            in2 => \_gnd_net_\,
            in3 => \N__42883\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15733\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_17_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43021\,
            in2 => \_gnd_net_\,
            in3 => \N__43015\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15734\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15735\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_18_lut_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43012\,
            in2 => \_gnd_net_\,
            in3 => \N__43003\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_19_lut_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43000\,
            in2 => \_gnd_net_\,
            in3 => \N__42994\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15736\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15737\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_20_lut_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42991\,
            in2 => \_gnd_net_\,
            in3 => \N__42982\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15737\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15738\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_21_lut_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42979\,
            in2 => \_gnd_net_\,
            in3 => \N__42973\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_22\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15738\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_22_lut_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42970\,
            in2 => \_gnd_net_\,
            in3 => \N__42961\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15739\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_23_lut_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42958\,
            in2 => \_gnd_net_\,
            in3 => \N__42952\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15740\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_24_lut_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42949\,
            in2 => \_gnd_net_\,
            in3 => \N__42943\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15741\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_25_lut_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43120\,
            in2 => \_gnd_net_\,
            in3 => \N__43114\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15742\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_26_lut_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43111\,
            in2 => \_gnd_net_\,
            in3 => \N__43099\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_27\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_27_lut_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43096\,
            in2 => \_gnd_net_\,
            in3 => \N__43090\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15744\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_28_lut_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43087\,
            in2 => \_gnd_net_\,
            in3 => \N__43075\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15745\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_29_lut_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43072\,
            in2 => \_gnd_net_\,
            in3 => \N__43060\,
            lcout => \Error_sub_temp_30_adj_2385\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15746\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_30_lut_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43057\,
            in2 => \_gnd_net_\,
            in3 => \N__43051\,
            lcout => \Error_sub_temp_31_adj_2384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_3_lut_4_lut_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__44822\,
            in1 => \N__44767\,
            in2 => \_gnd_net_\,
            in3 => \N__45120\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n188_adj_725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000100010"
        )
    port map (
            in0 => \N__44821\,
            in1 => \N__44766\,
            in2 => \_gnd_net_\,
            in3 => \N__45119\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__43144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__43152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43153\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45072\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43131\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43143\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__46554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__43132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64947\,
            in2 => \N__64638\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_1\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17987\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64588\,
            in2 => \N__43471\,
            in3 => \N__43180\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_2\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17987\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17988\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43444\,
            in2 => \N__64639\,
            in3 => \N__43177\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_3\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17988\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17989\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64592\,
            in2 => \N__43423\,
            in3 => \N__43174\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_4\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17989\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17990\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43399\,
            in2 => \N__64640\,
            in3 => \N__43171\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_5\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17990\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17991\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43708\,
            in2 => \N__64641\,
            in3 => \N__43168\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_6\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17991\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17992\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64599\,
            in2 => \N__43687\,
            in3 => \N__43165\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_7\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17992\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17993\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43663\,
            in2 => \N__64642\,
            in3 => \N__43162\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_8\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17993\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17994\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43642\,
            in2 => \N__64643\,
            in3 => \N__43159\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_9\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17995\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43621\,
            in2 => \N__64646\,
            in3 => \N__43156\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_10\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17995\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17996\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43600\,
            in2 => \N__64644\,
            in3 => \N__43261\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_11\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17996\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17997\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43579\,
            in2 => \N__64647\,
            in3 => \N__43258\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_12\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17997\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17998\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43558\,
            in2 => \N__64645\,
            in3 => \N__43255\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17998\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17999\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64612\,
            in2 => \N__43810\,
            in3 => \N__43252\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_14\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n17999\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18000\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43786\,
            in2 => \N__45325\,
            in3 => \N__43228\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n738_adj_718\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18000\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_LUT4_0_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43225\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64091\,
            in2 => \N__64381\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n57_adj_714\,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18017\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64323\,
            in2 => \N__43207\,
            in3 => \N__43195\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n106_adj_713\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18017\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18018\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43192\,
            in2 => \N__64382\,
            in3 => \N__43183\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n155_adj_712\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18018\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18019\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64327\,
            in2 => \N__43387\,
            in3 => \N__43375\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n204_adj_711\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18019\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18020\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43372\,
            in2 => \N__64383\,
            in3 => \N__43363\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n253_adj_710\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18020\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18021\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64331\,
            in2 => \N__43360\,
            in3 => \N__43348\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n302_adj_709\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18021\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18022\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43345\,
            in2 => \N__64384\,
            in3 => \N__43336\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n351_adj_708\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18022\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18023\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64335\,
            in2 => \N__43333\,
            in3 => \N__43321\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n400_adj_707\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18023\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18024\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43318\,
            in2 => \N__64437\,
            in3 => \N__43306\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n449_adj_706\,
            ltout => OPEN,
            carryin => \bfn_16_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18025\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64388\,
            in2 => \N__43303\,
            in3 => \N__43291\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n498_adj_705\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18025\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18026\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43288\,
            in2 => \N__64438\,
            in3 => \N__43279\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n547_adj_704\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18026\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18027\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64392\,
            in2 => \N__43276\,
            in3 => \N__43264\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n596_adj_703\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18027\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18028\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43546\,
            in2 => \N__64439\,
            in3 => \N__43537\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n645_adj_702\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18028\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18029\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64396\,
            in2 => \N__43534\,
            in3 => \N__43522\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n694_adj_701\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18029\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18030\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43519\,
            in2 => \N__45289\,
            in3 => \N__43495\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n746_adj_699\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18030\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_LUT4_0_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43492\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64453\,
            in2 => \N__65004\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n54\,
            ltout => OPEN,
            carryin => \bfn_16_27_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18002\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64964\,
            in2 => \N__43456\,
            in3 => \N__43435\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n103\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18002\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18003\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43432\,
            in2 => \N__65005\,
            in3 => \N__43411\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n152\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18003\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18004\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43408\,
            in2 => \N__65014\,
            in3 => \N__43390\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n201\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18004\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18005\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43717\,
            in2 => \N__65006\,
            in3 => \N__43699\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n250\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18005\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18006\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43696\,
            in2 => \N__65015\,
            in3 => \N__43675\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n299\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18006\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18007\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43672\,
            in2 => \N__65007\,
            in3 => \N__43654\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n348\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18007\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18008\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43651\,
            in2 => \N__65016\,
            in3 => \N__43633\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n397\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18008\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18009\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43630\,
            in2 => \N__65008\,
            in3 => \N__43612\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n446\,
            ltout => OPEN,
            carryin => \bfn_16_28_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18010\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43609\,
            in2 => \N__65011\,
            in3 => \N__43591\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n495\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18010\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18011\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43588\,
            in2 => \N__65009\,
            in3 => \N__43570\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n544\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18011\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18012\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43567\,
            in2 => \N__65012\,
            in3 => \N__43549\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n593\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18012\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18013\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43819\,
            in2 => \N__65010\,
            in3 => \N__43798\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n642\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18013\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18014\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43795\,
            in2 => \N__65013\,
            in3 => \N__43774\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n691_adj_717\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18014\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18015\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45310\,
            in2 => \N__43771\,
            in3 => \N__43747\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n742_adj_715\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18015\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_LUT4_0_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43744\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55663\,
            in2 => \N__55872\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n84\,
            ltout => OPEN,
            carryin => \bfn_17_5_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18135\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55823\,
            in2 => \N__43912\,
            in3 => \N__43726\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n133\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18135\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18136\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43891\,
            in2 => \N__55873\,
            in3 => \N__43723\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n182\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18136\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18137\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55827\,
            in2 => \N__43879\,
            in3 => \N__43720\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n231\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18137\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18138\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43864\,
            in2 => \N__55874\,
            in3 => \N__43852\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n280\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18138\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18139\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55831\,
            in2 => \N__44023\,
            in3 => \N__43849\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n329\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18139\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18140\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44003\,
            in2 => \N__55875\,
            in3 => \N__43846\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n378\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18140\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18141\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55835\,
            in2 => \N__44008\,
            in3 => \N__43843\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n427\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18141\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18142\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45654\,
            in2 => \N__44007\,
            in3 => \N__43840\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n782_adj_351\,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_LUT4_0_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43837\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__43834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43938\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__43833\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45582\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43923\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43939\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43924\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55233\,
            in2 => \N__55616\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n87_adj_400\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18167\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43897\,
            in2 => \N__55619\,
            in3 => \N__43882\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n136_adj_399\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18167\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18168\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43966\,
            in2 => \N__55617\,
            in3 => \N__43867\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n185_adj_398\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18168\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18169\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43975\,
            in2 => \N__55620\,
            in3 => \N__43855\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n234_adj_397\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18169\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18170\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43952\,
            in2 => \N__55618\,
            in3 => \N__44011\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n283\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18170\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18171\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55582\,
            in2 => \N__43959\,
            in3 => \N__43984\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n332\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18171\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18172\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45774\,
            in2 => \N__43960\,
            in3 => \N__43981\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n786_adj_348\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18172\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_LUT4_0_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43978\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i2_3_lut_4_lut_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__44152\,
            in1 => \N__44141\,
            in2 => \_gnd_net_\,
            in3 => \N__44058\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44140\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n138\,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__44139\,
            in1 => \N__55073\,
            in2 => \N__43969\,
            in3 => \N__54969\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_315_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50362\,
            lcout => n793,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__44166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_4_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000100010"
        )
    port map (
            in0 => \N__44057\,
            in1 => \N__44151\,
            in2 => \_gnd_net_\,
            in3 => \N__44138\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__44167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__51127\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50364\,
            lcout => n142_adj_2419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i11961_4_lut_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__55089\,
            in1 => \N__44142\,
            in2 => \N__55266\,
            in3 => \N__50363\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n4\,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_4_lut_4_lut_4_lut_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__44143\,
            in1 => \_gnd_net_\,
            in2 => \N__44098\,
            in3 => \N__44056\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_3_lut_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__44059\,
            in1 => \N__55267\,
            in2 => \N__44091\,
            in3 => \N__44087\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19269\,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_adj_135_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100111100"
        )
    port map (
            in0 => \N__44068\,
            in1 => \N__45756\,
            in2 => \N__44095\,
            in3 => \N__44062\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__55268\,
            in1 => \N__44060\,
            in2 => \N__44092\,
            in3 => \N__44086\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19273\,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_129_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010101000"
        )
    port map (
            in0 => \N__44061\,
            in1 => \N__45755\,
            in2 => \N__44032\,
            in3 => \N__44029\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51128\,
            lcout => n146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_3_lut_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__44323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44186\,
            lcout => OPEN,
            ltout => \foc.u_Park_Transform.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_4_lut_adj_307_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__44187\,
            in1 => \N__44239\,
            in2 => \N__44470\,
            in3 => \N__44437\,
            lcout => \foc.u_Park_Transform.n791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_4_lut_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010001000"
        )
    port map (
            in0 => \N__44318\,
            in1 => \N__44368\,
            in2 => \N__44350\,
            in3 => \N__44225\,
            lcout => OPEN,
            ltout => \foc.u_Park_Transform.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i2_4_lut_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__44226\,
            in1 => \N__44349\,
            in2 => \N__44440\,
            in3 => \N__44319\,
            lcout => \foc.u_Park_Transform.n19845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.Alpha_15__I_0_11_i28_2_lut_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__44422\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n628,
            ltout => \n628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_4_lut_adj_305_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011100000"
        )
    port map (
            in0 => \N__44364\,
            in1 => \N__44313\,
            in2 => \N__44353\,
            in3 => \N__44340\,
            lcout => OPEN,
            ltout => \foc.u_Park_Transform.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_Park_Transform.i1_4_lut_adj_306_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010101000"
        )
    port map (
            in0 => \N__44314\,
            in1 => \N__44224\,
            in2 => \N__44197\,
            in3 => \N__44194\,
            lcout => \foc.u_Park_Transform.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60856\,
            in2 => \N__67442\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n66_adj_433\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44503\,
            in2 => \N__58905\,
            in3 => \N__44497\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n112\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17781\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48322\,
            in2 => \N__54806\,
            in3 => \N__44494\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n161\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17782\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48301\,
            in2 => \N__54516\,
            in3 => \N__44491\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n210\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17783\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48277\,
            in2 => \N__54248\,
            in3 => \N__44488\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n259\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17784\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48256\,
            in2 => \N__53990\,
            in3 => \N__44485\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n308_adj_368\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17785\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53680\,
            in2 => \N__48235\,
            in3 => \N__44482\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n357_adj_366\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17786\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53316\,
            in2 => \N__48211\,
            in3 => \N__44479\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n406_adj_363\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17787\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48187\,
            in2 => \N__53140\,
            in3 => \N__44476\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n455_adj_350\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48472\,
            in2 => \N__56182\,
            in3 => \N__44473\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n504\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17789\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48451\,
            in2 => \N__55944\,
            in3 => \N__44542\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n553\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17790\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48430\,
            in2 => \N__55723\,
            in3 => \N__44539\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n602\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17791\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48409\,
            in2 => \N__55348\,
            in3 => \N__44536\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n651_adj_474\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17792\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55181\,
            in2 => \N__48388\,
            in3 => \N__44533\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n700_adj_455\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17793\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54946\,
            in2 => \N__48361\,
            in3 => \N__44530\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n754\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17794\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_LUT4_0_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44527\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60966\,
            in2 => \N__67397\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n63_adj_384\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44524\,
            in2 => \N__58907\,
            in3 => \N__44518\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n109_adj_383\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17766\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44515\,
            in2 => \N__54813\,
            in3 => \N__44506\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n158_adj_375\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17767\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44656\,
            in2 => \N__54530\,
            in3 => \N__44647\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n207\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17768\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44644\,
            in2 => \N__54250\,
            in3 => \N__44635\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n256\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17769\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44632\,
            in2 => \N__54000\,
            in3 => \N__44623\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n305\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17770\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44620\,
            in2 => \N__53722\,
            in3 => \N__44611\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n354_adj_367\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17771\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53426\,
            in2 => \N__44608\,
            in3 => \N__44596\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n403_adj_365\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17772\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44593\,
            in2 => \N__53210\,
            in3 => \N__44584\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n452_adj_362\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44581\,
            in2 => \N__56204\,
            in3 => \N__44572\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n501\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17774\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55960\,
            in2 => \N__44569\,
            in3 => \N__44557\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n550\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17775\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44554\,
            in2 => \N__55738\,
            in3 => \N__44545\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n599\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17776\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44737\,
            in2 => \N__55337\,
            in3 => \N__44728\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n648_adj_347\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17777\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55182\,
            in2 => \N__44725\,
            in3 => \N__44713\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n697\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17778\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54958\,
            in2 => \N__44710\,
            in3 => \N__44698\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n750\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17779\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_LUT4_0_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44695\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44748\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__48940\,
            in1 => \_gnd_net_\,
            in2 => \N__44956\,
            in3 => \N__45051\,
            lcout => n142_adj_2422,
            ltout => \n142_adj_2422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_3_lut_4_lut_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__44765\,
            in1 => \_gnd_net_\,
            in2 => \N__44692\,
            in3 => \N__45129\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755\,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_292_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44785\,
            in2 => \N__44671\,
            in3 => \N__45128\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n14_adj_756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44997\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48939\,
            in2 => \_gnd_net_\,
            in3 => \N__44942\,
            lcout => n146_adj_2423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_3_lut_4_lut_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__44807\,
            in1 => \N__44764\,
            in2 => \_gnd_net_\,
            in3 => \N__45127\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n6_adj_763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_adj_275_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__45122\,
            in1 => \N__65438\,
            in2 => \N__65264\,
            in3 => \N__65061\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n139_adj_727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45123\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_312_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45048\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n141_adj_2421,
            ltout => \n141_adj_2421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i12085_4_lut_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__65437\,
            in1 => \N__45121\,
            in2 => \N__44770\,
            in3 => \N__45047\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_220_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__50922\,
            in1 => \N__52785\,
            in2 => \N__50708\,
            in3 => \N__44983\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44749\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__46785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_218_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__44971\,
            in1 => \N__59181\,
            in2 => \N__51009\,
            in3 => \N__51042\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_219_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__51190\,
            in1 => \N__59466\,
            in2 => \N__44986\,
            in3 => \N__52641\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_216_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46621\,
            in1 => \N__46651\,
            in2 => \N__46687\,
            in3 => \N__46747\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_217_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46716\,
            in1 => \N__46591\,
            in2 => \N__44977\,
            in3 => \N__46774\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1213_4_lut_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__48840\,
            in1 => \N__48819\,
            in2 => \N__44974\,
            in3 => \N__48867\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_211_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__44962\,
            in1 => \N__59465\,
            in2 => \N__51197\,
            in3 => \N__52640\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19827_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_212_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__50915\,
            in1 => \N__52772\,
            in2 => \N__44965\,
            in3 => \N__50693\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_210_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__48839\,
            in1 => \N__51041\,
            in2 => \N__51008\,
            in3 => \N__59180\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45148\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46573\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46518\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i537_2_lut_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45133\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45076\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_313_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__45055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n793_adj_2424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45022\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i31_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58367\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45004\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51082\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45321\,
            in2 => \N__65017\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n93\,
            ltout => OPEN,
            carryin => \bfn_17_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18369\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45303\,
            in2 => \N__64452\,
            in3 => \N__45292\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n142\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18369\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18370\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45282\,
            in2 => \N__64090\,
            in3 => \N__45271\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n191\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18370\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18371\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45258\,
            in2 => \N__63929\,
            in3 => \N__45244\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n240\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18371\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18372\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45237\,
            in2 => \N__63626\,
            in3 => \N__45220\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n289\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18372\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18373\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45213\,
            in2 => \N__63279\,
            in3 => \N__45196\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n338\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18373\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18374\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45189\,
            in2 => \N__62959\,
            in3 => \N__45172\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n387\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18374\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18375\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45162\,
            in2 => \N__66876\,
            in3 => \N__45151\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n436\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18375\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18376\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45477\,
            in2 => \N__66604\,
            in3 => \N__45460\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n485\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18377\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45456\,
            in2 => \N__66345\,
            in3 => \N__45433\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n534\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18377\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18378\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45430\,
            in2 => \N__66063\,
            in3 => \N__45406\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n583\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18378\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18379\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45403\,
            in2 => \N__65808\,
            in3 => \N__45382\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n632\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18379\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18380\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65492\,
            in2 => \N__45379\,
            in3 => \N__45358\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n681\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18380\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18381\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65313\,
            in2 => \N__45355\,
            in3 => \N__45343\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n730\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18381\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18382\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45340\,
            in2 => \N__65152\,
            in3 => \N__45331\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n794\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18382\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_LUT4_0_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45328\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55839\,
            in2 => \N__56145\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n81\,
            ltout => OPEN,
            carryin => \bfn_18_5_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17266\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_18_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56094\,
            in2 => \N__45562\,
            in3 => \N__45553\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n130\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17266\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17267\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_18_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45550\,
            in2 => \N__56146\,
            in3 => \N__45544\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n179\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17267\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17268\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56098\,
            in2 => \N__45541\,
            in3 => \N__45532\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n228\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17268\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17269\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45529\,
            in2 => \N__56147\,
            in3 => \N__45523\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n277\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17269\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17270\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56102\,
            in2 => \N__45520\,
            in3 => \N__45511\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n326\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17270\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17271\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45508\,
            in2 => \N__56148\,
            in3 => \N__45502\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n375\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17271\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17272\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_18_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56106\,
            in2 => \N__45499\,
            in3 => \N__45490\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n424\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17272\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17273\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45632\,
            in2 => \N__56038\,
            in3 => \N__45487\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n473\,
            ltout => OPEN,
            carryin => \bfn_18_6_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17274\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56013\,
            in2 => \N__45639\,
            in3 => \N__45643\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n522\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17274\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17275\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45672\,
            in2 => \N__45640\,
            in3 => \N__45619\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n778_adj_356\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17275\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_LUT4_0_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45616\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__45595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45613\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__45594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45583\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61236\,
            in2 => \N__60862\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n93\,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17942\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58983\,
            in2 => \N__58810\,
            in3 => \N__45568\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n142_adj_414\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17942\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17943\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52572\,
            in2 => \N__54625\,
            in3 => \N__45565\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n191\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17943\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17944\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52344\,
            in2 => \N__54386\,
            in3 => \N__45697\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n240\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17944\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17945\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50154\,
            in2 => \N__54080\,
            in3 => \N__45694\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n289\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17945\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17946\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52062\,
            in2 => \N__53819\,
            in3 => \N__45691\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n338\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17946\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17947\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49956\,
            in2 => \N__53585\,
            in3 => \N__45688\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n387\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17947\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17948\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47679\,
            in2 => \N__53427\,
            in3 => \N__45685\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n436\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17948\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17949\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47472\,
            in2 => \N__53075\,
            in3 => \N__45682\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n485\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17950\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49794\,
            in2 => \N__56090\,
            in3 => \N__45679\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n534\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17950\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17951\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45676\,
            in2 => \N__55915\,
            in3 => \N__45661\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n583\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17951\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17952\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45658\,
            in2 => \N__55615\,
            in3 => \N__45778\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n632\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17952\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17953\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55229\,
            in2 => \N__45775\,
            in3 => \N__45760\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n681\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17953\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17954\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55093\,
            in2 => \N__45757\,
            in3 => \N__45730\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n730\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17954\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17955\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45727\,
            in2 => \N__55005\,
            in3 => \N__45721\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n794_adj_413\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17955\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_LUT4_0_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45718\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60839\,
            in2 => \N__67296\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n84_adj_389\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17882\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58755\,
            in2 => \N__45715\,
            in3 => \N__45706\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n130_adj_453\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17882\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17883\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50125\,
            in2 => \N__54680\,
            in3 => \N__45703\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n179_adj_452\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17883\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17884\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50104\,
            in2 => \N__54480\,
            in3 => \N__45700\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n228_adj_450\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17884\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17885\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50083\,
            in2 => \N__54156\,
            in3 => \N__45805\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n277_adj_448\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17885\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17886\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50062\,
            in2 => \N__53937\,
            in3 => \N__45802\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n326_adj_443\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17886\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17887\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50038\,
            in2 => \N__53636\,
            in3 => \N__45799\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n375_adj_438\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17887\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17888\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50311\,
            in2 => \N__53373\,
            in3 => \N__45796\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n424_adj_435\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17888\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17889\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50290\,
            in2 => \N__53088\,
            in3 => \N__45793\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n473_adj_431\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17890\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50272\,
            in2 => \N__56149\,
            in3 => \N__45790\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n522_adj_430\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17890\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17891\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50251\,
            in2 => \N__55916\,
            in3 => \N__45787\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n571\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17891\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17892\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50230\,
            in2 => \N__55659\,
            in3 => \N__45784\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n620\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17892\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17893\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50209\,
            in2 => \N__55306\,
            in3 => \N__45781\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n669\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17893\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17894\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55122\,
            in2 => \N__50188\,
            in3 => \N__45871\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n718\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17894\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17895\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54914\,
            in2 => \N__50434\,
            in3 => \N__45868\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n778\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17895\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_LUT4_0_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45865\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60903\,
            in2 => \N__67351\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n81_adj_457\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17867\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45862\,
            in2 => \N__58870\,
            in3 => \N__45856\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n127_adj_479\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17867\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17868\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45853\,
            in2 => \N__54771\,
            in3 => \N__45844\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n176_adj_478\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17868\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17869\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45841\,
            in2 => \N__54481\,
            in3 => \N__45832\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n225_adj_477\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17869\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17870\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45829\,
            in2 => \N__54207\,
            in3 => \N__45820\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n274_adj_476\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17870\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17871\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45817\,
            in2 => \N__53970\,
            in3 => \N__45808\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n323_adj_475\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17871\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17872\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53637\,
            in2 => \N__45985\,
            in3 => \N__45973\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n372_adj_473\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17872\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17873\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45970\,
            in2 => \N__53408\,
            in3 => \N__45961\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n421_adj_465\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17873\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17874\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45958\,
            in2 => \N__53189\,
            in3 => \N__45949\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n470_adj_463\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17875\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45946\,
            in2 => \N__56150\,
            in3 => \N__45937\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n519_adj_461\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17875\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17876\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45934\,
            in2 => \N__55918\,
            in3 => \N__45925\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n568_adj_460\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17876\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17877\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45922\,
            in2 => \N__55698\,
            in3 => \N__45913\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n617_adj_459\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17877\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17878\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45910\,
            in2 => \N__55341\,
            in3 => \N__45901\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n666\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17878\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17879\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55125\,
            in2 => \N__45898\,
            in3 => \N__45883\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n715\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17879\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17880\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45880\,
            in2 => \N__54945\,
            in3 => \N__46063\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n774\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17880\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_LUT4_0_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46060\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60958\,
            in2 => \N__67396\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n78_adj_480\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17841\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46057\,
            in2 => \N__58874\,
            in3 => \N__46051\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n124_adj_507\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17841\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17842\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46048\,
            in2 => \N__54773\,
            in3 => \N__46039\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n173_adj_506\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17842\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17843\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46036\,
            in2 => \N__54526\,
            in3 => \N__46027\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n222_adj_505\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17843\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17844\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46024\,
            in2 => \N__54220\,
            in3 => \N__46015\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n271_adj_503\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17844\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17845\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46012\,
            in2 => \N__53991\,
            in3 => \N__46003\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n320_adj_502\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17845\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17846\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53650\,
            in2 => \N__46000\,
            in3 => \N__45988\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n369_adj_501\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17846\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17847\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46171\,
            in2 => \N__53469\,
            in3 => \N__46162\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n418_adj_500\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17847\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17848\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46159\,
            in2 => \N__53211\,
            in3 => \N__46150\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n467_adj_499\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17849\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46147\,
            in2 => \N__56190\,
            in3 => \N__46138\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n516_adj_498\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17849\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17850\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46135\,
            in2 => \N__55945\,
            in3 => \N__46126\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n565_adj_497\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17850\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17851\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46123\,
            in2 => \N__55724\,
            in3 => \N__46114\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n614_adj_496\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17851\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17852\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46111\,
            in2 => \N__55349\,
            in3 => \N__46102\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n663_adj_494\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17852\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17853\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55150\,
            in2 => \N__46099\,
            in3 => \N__46084\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n712_adj_493\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17853\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17854\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54959\,
            in2 => \N__46081\,
            in3 => \N__46069\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n770\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17854\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_LUT4_0_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46066\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60959\,
            in2 => \N__67465\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n75\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17826\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46255\,
            in2 => \N__58906\,
            in3 => \N__46249\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n121\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17826\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17827\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46246\,
            in2 => \N__54802\,
            in3 => \N__46237\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n170\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17827\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17828\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46234\,
            in2 => \N__54517\,
            in3 => \N__46225\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n219\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17828\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17829\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46222\,
            in2 => \N__54249\,
            in3 => \N__46213\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n268_adj_437\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17829\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17830\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46210\,
            in2 => \N__53992\,
            in3 => \N__46201\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n317_adj_428\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17830\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17831\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46198\,
            in2 => \N__53707\,
            in3 => \N__46189\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n366_adj_426\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17831\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17832\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53474\,
            in2 => \N__46186\,
            in3 => \N__46174\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n415\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17832\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17833\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46345\,
            in2 => \N__53190\,
            in3 => \N__46336\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n464_adj_423\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17834\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46333\,
            in2 => \N__56207\,
            in3 => \N__46324\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n513_adj_412\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17834\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17835\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46321\,
            in2 => \N__55946\,
            in3 => \N__46312\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n562_adj_378\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17835\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17836\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46309\,
            in2 => \N__55725\,
            in3 => \N__46300\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n611_adj_373\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17836\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17837\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46297\,
            in2 => \N__55378\,
            in3 => \N__46288\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n660_adj_372\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17837\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17838\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46285\,
            in2 => \N__55180\,
            in3 => \N__46276\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n709\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17838\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17839\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54987\,
            in2 => \N__46273\,
            in3 => \N__46261\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n766\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17839\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_LUT4_0_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46258\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60967\,
            in2 => \N__67466\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n60\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46423\,
            in2 => \N__58908\,
            in3 => \N__46417\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n106\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17751\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46414\,
            in2 => \N__54804\,
            in3 => \N__46408\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n155_adj_369\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17752\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54521\,
            in2 => \N__46405\,
            in3 => \N__46396\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n204_adj_361\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17753\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46393\,
            in2 => \N__54251\,
            in3 => \N__46387\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n253\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17754\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46384\,
            in2 => \N__54001\,
            in3 => \N__46378\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n302_adj_364\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17755\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46375\,
            in2 => \N__53711\,
            in3 => \N__46369\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n351\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17756\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53479\,
            in2 => \N__46366\,
            in3 => \N__46357\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n400_adj_511\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17757\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46354\,
            in2 => \N__53215\,
            in3 => \N__46348\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n449_adj_492\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46495\,
            in2 => \N__56205\,
            in3 => \N__46489\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n498_adj_469\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17759\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46486\,
            in2 => \N__55966\,
            in3 => \N__46480\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n547_adj_454\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17760\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46477\,
            in2 => \N__55736\,
            in3 => \N__46471\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n596_adj_434\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17761\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46468\,
            in2 => \N__55363\,
            in3 => \N__46462\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n645_adj_429\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17762\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55186\,
            in2 => \N__46459\,
            in3 => \N__46450\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n694_adj_427\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17763\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54988\,
            in2 => \N__46447\,
            in3 => \N__46438\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n746\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17764\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_LUT4_0_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46435\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_221_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__59351\,
            in1 => \N__59151\,
            in2 => \N__50655\,
            in3 => \N__46432\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_222_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__52929\,
            in1 => \N__52704\,
            in2 => \N__46426\,
            in3 => \N__52746\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_223_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50976\,
            in1 => \N__50873\,
            in2 => \N__46576\,
            in3 => \N__50949\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_215_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__50948\,
            in1 => \N__46525\,
            in2 => \N__50877\,
            in3 => \N__50975\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46572\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46555\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_213_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__59350\,
            in1 => \N__59150\,
            in2 => \N__50654\,
            in3 => \N__46537\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_214_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__52928\,
            in1 => \N__52703\,
            in2 => \N__46528\,
            in3 => \N__52745\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46519\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i15877_4_lut_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46683\,
            in1 => \N__46746\,
            in2 => \N__46717\,
            in3 => \N__46773\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i15889_4_lut_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46620\,
            in1 => \N__46590\,
            in2 => \N__46498\,
            in3 => \N__46650\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20870\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46789\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_2_lut_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__56913\,
            in1 => \N__57384\,
            in2 => \N__64693\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20174\,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15883\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_3_lut_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57333\,
            in2 => \N__46762\,
            in3 => \N__46735\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15883\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15884\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_4_lut_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57297\,
            in2 => \N__46732\,
            in3 => \N__46702\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15884\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15885\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_5_lut_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46699\,
            in2 => \N__57276\,
            in3 => \N__46672\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15885\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15886\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_6_lut_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57219\,
            in2 => \N__46669\,
            in3 => \N__46639\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15886\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15887\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_7_lut_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57195\,
            in2 => \N__46636\,
            in3 => \N__46609\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15887\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15888\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_8_lut_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57153\,
            in2 => \N__46606\,
            in3 => \N__46579\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15888\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15889\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_9_lut_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57114\,
            in2 => \N__46927\,
            in3 => \N__46912\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15889\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15890\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_10_lut_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57852\,
            in2 => \N__46909\,
            in3 => \N__46897\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9\,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15891\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_11_lut_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57813\,
            in2 => \N__46894\,
            in3 => \N__46879\,
            lcout => \foc.preSatVoltage_10\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15891\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15892\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_12_lut_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57744\,
            in2 => \N__46876\,
            in3 => \N__46861\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15892\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15893\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_13_lut_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57684\,
            in2 => \N__46858\,
            in3 => \N__46843\,
            lcout => \foc.preSatVoltage_12\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15893\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15894\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_14_lut_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57600\,
            in2 => \N__46840\,
            in3 => \N__46825\,
            lcout => \foc.preSatVoltage_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15894\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15895\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_15_lut_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57525\,
            in2 => \N__46822\,
            in3 => \N__46807\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15895\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15896\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_16_lut_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46804\,
            in2 => \N__57463\,
            in3 => \N__46792\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15896\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15897\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_17_lut_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58278\,
            in2 => \N__47104\,
            in3 => \N__47089\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15897\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15898\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_18_lut_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47086\,
            in2 => \N__58213\,
            in3 => \N__47074\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17\,
            ltout => OPEN,
            carryin => \bfn_18_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15899\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_19_lut_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58147\,
            in2 => \N__47071\,
            in3 => \N__47053\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15899\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15900\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_20_lut_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58080\,
            in2 => \N__47050\,
            in3 => \N__47032\,
            lcout => \foc.preSatVoltage_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15900\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15901\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_21_lut_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47029\,
            in2 => \N__58011\,
            in3 => \N__47014\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15901\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15902\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_22_lut_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57964\,
            in2 => \N__47011\,
            in3 => \N__46993\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15902\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15903\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_23_lut_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57909\,
            in2 => \N__46990\,
            in3 => \N__46972\,
            lcout => \foc.preSatVoltage_22\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15903\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15904\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_24_lut_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58512\,
            in2 => \N__46969\,
            in3 => \N__46951\,
            lcout => \foc.preSatVoltage_23\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15904\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15905\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_25_lut_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58433\,
            in2 => \N__46948\,
            in3 => \N__46930\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15905\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15906\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_26_lut_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58434\,
            in2 => \N__47233\,
            in3 => \N__47218\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_25\,
            ltout => OPEN,
            carryin => \bfn_18_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15907\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_27_lut_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47215\,
            in2 => \N__58450\,
            in3 => \N__47203\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15907\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15908\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_28_lut_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58438\,
            in2 => \N__47200\,
            in3 => \N__47182\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15908\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15909\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_29_lut_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47179\,
            in2 => \N__58451\,
            in3 => \N__47164\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15909\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15910\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_30_lut_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58442\,
            in2 => \N__47161\,
            in3 => \N__47143\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15910\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15911\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_31_lut_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47140\,
            in2 => \N__58452\,
            in3 => \N__47125\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_30\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15911\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15912\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_32_lut_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47122\,
            in1 => \N__58446\,
            in2 => \_gnd_net_\,
            in3 => \N__47107\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Voltage_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64921\,
            in2 => \N__64726\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18354\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64440\,
            in2 => \N__47326\,
            in3 => \N__47317\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n139\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18354\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18355\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64132\,
            in2 => \N__47314\,
            in3 => \N__47305\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n188\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18355\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18356\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63862\,
            in2 => \N__47302\,
            in3 => \N__47293\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n237\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18356\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18357\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47290\,
            in2 => \N__63608\,
            in3 => \N__47284\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n286\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18357\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18358\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47281\,
            in2 => \N__63361\,
            in3 => \N__47275\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n335\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18358\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18359\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47272\,
            in2 => \N__62974\,
            in3 => \N__47266\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n384\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18359\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18360\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_18_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47263\,
            in2 => \N__66824\,
            in3 => \N__47257\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n433\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18360\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18361\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_18_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47254\,
            in2 => \N__66629\,
            in3 => \N__47245\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n482\,
            ltout => OPEN,
            carryin => \bfn_18_27_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18362\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47242\,
            in2 => \N__66327\,
            in3 => \N__47236\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n531\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18362\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18363\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47380\,
            in2 => \N__66090\,
            in3 => \N__47374\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n580\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18363\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18364\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_18_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47371\,
            in2 => \N__65807\,
            in3 => \N__47365\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n629\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18364\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18365\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_18_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47362\,
            in2 => \N__65580\,
            in3 => \N__47356\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n678\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18365\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18366\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65341\,
            in2 => \N__47353\,
            in3 => \N__47344\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n727\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18366\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18367\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_18_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47341\,
            in2 => \N__65188\,
            in3 => \N__47335\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n790\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18367\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_LUT4_0_LC_18_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47332\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53147\,
            in2 => \N__53464\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n75_adj_510\,
            ltout => OPEN,
            carryin => \bfn_19_5_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17641\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53434\,
            in2 => \N__49441\,
            in3 => \N__47329\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n124\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17641\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17642\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49708\,
            in2 => \N__53465\,
            in3 => \N__47407\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n173\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17642\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17643\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53438\,
            in2 => \N__49690\,
            in3 => \N__47404\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n222\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17643\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17644\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_19_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49666\,
            in2 => \N__53466\,
            in3 => \N__47401\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n271\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17644\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17645\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_19_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49648\,
            in2 => \N__53468\,
            in3 => \N__47398\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n320\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17645\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17646\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_19_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49627\,
            in2 => \N__53467\,
            in3 => \N__47395\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n369\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17646\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17647\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53445\,
            in2 => \N__49606\,
            in3 => \N__47392\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n418\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17647\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17648\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53378\,
            in2 => \N__49585\,
            in3 => \N__47389\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n467\,
            ltout => OPEN,
            carryin => \bfn_19_6_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17649\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49561\,
            in2 => \N__53428\,
            in3 => \N__47386\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n516\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17649\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17650\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53382\,
            in2 => \N__49837\,
            in3 => \N__47383\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n565\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17650\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17651\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49825\,
            in2 => \N__53429\,
            in3 => \N__47488\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n614\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17651\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17652\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53386\,
            in2 => \N__49816\,
            in3 => \N__47485\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n663\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17652\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17653\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49814\,
            in2 => \N__53430\,
            in3 => \N__47482\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n712\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17653\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17654\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_19_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49815\,
            in2 => \N__47479\,
            in3 => \N__47455\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n770_adj_381\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17654\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_LUT4_0_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47452\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53377\,
            in2 => \N__53607\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n72_adj_508\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17626\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53559\,
            in2 => \N__47449\,
            in3 => \N__47437\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n121_adj_504\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17626\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17627\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47434\,
            in2 => \N__53608\,
            in3 => \N__47425\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n170_adj_490\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17627\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17628\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53563\,
            in2 => \N__47422\,
            in3 => \N__47410\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n219_adj_472\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17628\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17629\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47608\,
            in2 => \N__53609\,
            in3 => \N__47599\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n268\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17629\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17630\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53567\,
            in2 => \N__47596\,
            in3 => \N__47584\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n317\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17630\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17631\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53568\,
            in2 => \N__47581\,
            in3 => \N__47569\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n366\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17631\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17632\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47566\,
            in2 => \N__53610\,
            in3 => \N__47557\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n415_adj_449\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17632\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17633\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47554\,
            in2 => \N__53693\,
            in3 => \N__47545\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n464\,
            ltout => OPEN,
            carryin => \bfn_19_8_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17634\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53657\,
            in2 => \N__47542\,
            in3 => \N__47530\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n513\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17634\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17635\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47527\,
            in2 => \N__53694\,
            in3 => \N__47518\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n562\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17635\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17636\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53661\,
            in2 => \N__47515\,
            in3 => \N__47503\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n611\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17636\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17637\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47500\,
            in2 => \N__53695\,
            in3 => \N__47491\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n660\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17637\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17638\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53665\,
            in2 => \N__47695\,
            in3 => \N__47683\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n709_adj_512\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17638\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17639\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47680\,
            in2 => \N__47668\,
            in3 => \N__47656\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n766_adj_385\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17639\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_LUT4_0_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47653\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60796\,
            in2 => \N__67404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_9_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17927\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47650\,
            in2 => \N__58845\,
            in3 => \N__47644\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n139_adj_419\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17927\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17928\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47641\,
            in2 => \N__54714\,
            in3 => \N__47635\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n188_adj_418\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17928\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17929\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54433\,
            in2 => \N__47632\,
            in3 => \N__47623\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n237_adj_417\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17929\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17930\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54175\,
            in2 => \N__47620\,
            in3 => \N__47611\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n286\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17930\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17931\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47785\,
            in2 => \N__53938\,
            in3 => \N__47779\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n335\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17931\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17932\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47776\,
            in2 => \N__53706\,
            in3 => \N__47770\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n384\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17932\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17933\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47767\,
            in2 => \N__53284\,
            in3 => \N__47761\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n433\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17933\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17934\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53089\,
            in2 => \N__47758\,
            in3 => \N__47746\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n482\,
            ltout => OPEN,
            carryin => \bfn_19_10_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17935\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47743\,
            in2 => \N__56160\,
            in3 => \N__47737\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n531\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17935\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17936\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47734\,
            in2 => \N__55917\,
            in3 => \N__47728\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n580\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17936\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17937\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47725\,
            in2 => \N__55697\,
            in3 => \N__47719\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n629\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17937\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17938\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47716\,
            in2 => \N__55356\,
            in3 => \N__47710\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n678\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17938\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17939\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55123\,
            in2 => \N__47707\,
            in3 => \N__47698\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n727\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17939\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17940\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54996\,
            in2 => \N__47860\,
            in3 => \N__47851\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n790_adj_415\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17940\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_LUT4_0_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47848\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60828\,
            in2 => \N__67405\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n90_adj_420\,
            ltout => OPEN,
            carryin => \bfn_19_11_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17912\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58780\,
            in2 => \N__47845\,
            in3 => \N__47836\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n136\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17912\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17913\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47833\,
            in2 => \N__54772\,
            in3 => \N__47824\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n185\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17913\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17914\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47821\,
            in2 => \N__54501\,
            in3 => \N__47812\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n234\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17914\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17915\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47809\,
            in2 => \N__54256\,
            in3 => \N__47800\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n283_adj_514\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17915\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17916\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47797\,
            in2 => \N__53942\,
            in3 => \N__47788\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n332_adj_513\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17916\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17917\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47977\,
            in2 => \N__53715\,
            in3 => \N__47968\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n381\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17917\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17918\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47965\,
            in2 => \N__53409\,
            in3 => \N__47956\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n430\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17918\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17919\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47953\,
            in2 => \N__53201\,
            in3 => \N__47944\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n479\,
            ltout => OPEN,
            carryin => \bfn_19_12_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17920\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47941\,
            in2 => \N__56197\,
            in3 => \N__47932\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n528\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17920\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17921\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47929\,
            in2 => \N__55939\,
            in3 => \N__47920\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n577\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17921\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17922\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47917\,
            in2 => \N__55717\,
            in3 => \N__47908\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n626\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17922\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17923\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47905\,
            in2 => \N__55364\,
            in3 => \N__47896\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n675\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17923\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17924\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55124\,
            in2 => \N__47893\,
            in3 => \N__47878\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n724\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17924\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17925\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54940\,
            in2 => \N__47875\,
            in3 => \N__47863\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n786\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17925\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_LUT4_0_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48055\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60857\,
            in2 => \N__67395\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n72\,
            ltout => OPEN,
            carryin => \bfn_19_13_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58866\,
            in2 => \N__48052\,
            in3 => \N__48043\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n118\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17811\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48040\,
            in2 => \N__54774\,
            in3 => \N__48031\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n167\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17812\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48028\,
            in2 => \N__54525\,
            in3 => \N__48019\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n216\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17813\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17814\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48016\,
            in2 => \N__54255\,
            in3 => \N__48007\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n265\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17814\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17815\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48004\,
            in2 => \N__53969\,
            in3 => \N__47995\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n314_adj_401\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17815\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53705\,
            in2 => \N__47992\,
            in3 => \N__47980\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n363_adj_380\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17816\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17817\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48172\,
            in2 => \N__53410\,
            in3 => \N__48160\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n412\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17817\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17818\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53130\,
            in2 => \N__48157\,
            in3 => \N__48145\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n461\,
            ltout => OPEN,
            carryin => \bfn_19_14_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17819\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48142\,
            in2 => \N__56189\,
            in3 => \N__48130\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n510\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17819\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17820\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48127\,
            in2 => \N__55956\,
            in3 => \N__48118\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n559_adj_358\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17820\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17821\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48115\,
            in2 => \N__55729\,
            in3 => \N__48106\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n608_adj_377\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17821\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17822\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55370\,
            in2 => \N__48103\,
            in3 => \N__48091\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n657_adj_360\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17822\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17823\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48088\,
            in2 => \N__55166\,
            in3 => \N__48076\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n706_adj_371\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17823\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17824\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54989\,
            in2 => \N__48073\,
            in3 => \N__48061\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n762\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17824\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_LUT4_0_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48058\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60858\,
            in2 => \N__67455\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n69\,
            ltout => OPEN,
            carryin => \bfn_19_15_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48328\,
            in2 => \N__58904\,
            in3 => \N__48313\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n115\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17796\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48310\,
            in2 => \N__54803\,
            in3 => \N__48292\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n164\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17797\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54508\,
            in2 => \N__48289\,
            in3 => \N__48268\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n213\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17798\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48265\,
            in2 => \N__54264\,
            in3 => \N__48247\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n262_adj_425\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17799\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48244\,
            in2 => \N__53986\,
            in3 => \N__48223\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n311_adj_422\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17800\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48220\,
            in2 => \N__53728\,
            in3 => \N__48199\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n360\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17801\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48196\,
            in2 => \N__53470\,
            in3 => \N__48175\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n409\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17802\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53206\,
            in2 => \N__48484\,
            in3 => \N__48463\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n458\,
            ltout => OPEN,
            carryin => \bfn_19_16_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48460\,
            in2 => \N__56206\,
            in3 => \N__48442\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n507\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17804\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48439\,
            in2 => \N__55965\,
            in3 => \N__48421\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n556_adj_370\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17805\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17806\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48418\,
            in2 => \N__55722\,
            in3 => \N__48400\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n605_adj_462\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17806\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17807\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48397\,
            in2 => \N__55366\,
            in3 => \N__48376\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n654_adj_456\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17807\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17808\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55151\,
            in2 => \N__48373\,
            in3 => \N__48349\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n703_adj_359\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17808\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54997\,
            in2 => \N__48346\,
            in3 => \N__48334\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n758\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17809\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_LUT4_0_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48331\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_1_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51093\,
            in2 => \N__51097\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17711\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_2_lut_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55486\,
            in1 => \_gnd_net_\,
            in2 => \N__51158\,
            in3 => \N__48610\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17711\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17712\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_3_lut_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55490\,
            in1 => \N__50896\,
            in2 => \N__54862\,
            in3 => \N__48607\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17712\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17713\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_4_lut_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55487\,
            in1 => \N__48604\,
            in2 => \N__54841\,
            in3 => \N__48595\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17713\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17714\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_5_lut_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55491\,
            in1 => \N__48592\,
            in2 => \N__48580\,
            in3 => \N__48565\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17714\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17715\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_6_lut_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55488\,
            in1 => \N__48562\,
            in2 => \N__48547\,
            in3 => \N__48532\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17715\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_7_lut_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55492\,
            in1 => \N__48529\,
            in2 => \N__48523\,
            in3 => \N__48508\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17716\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17717\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_8_lut_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55489\,
            in1 => \N__48505\,
            in2 => \N__48496\,
            in3 => \N__48487\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_22\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17717\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17718\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_9_lut_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55512\,
            in1 => \N__48808\,
            in2 => \N__48799\,
            in3 => \N__48790\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_23\,
            ltout => OPEN,
            carryin => \bfn_19_18_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17719\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_10_lut_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55493\,
            in1 => \N__48787\,
            in2 => \N__48778\,
            in3 => \N__48769\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17719\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17720\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_11_lut_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55509\,
            in1 => \N__48766\,
            in2 => \N__48754\,
            in3 => \N__48739\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17720\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17721\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_12_lut_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55494\,
            in1 => \N__48736\,
            in2 => \N__48721\,
            in3 => \N__48706\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17721\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17722\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_13_lut_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55510\,
            in1 => \N__50404\,
            in2 => \N__48703\,
            in3 => \N__48688\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17722\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17723\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_14_lut_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55495\,
            in1 => \N__48685\,
            in2 => \N__50386\,
            in3 => \N__48676\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17723\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17724\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_15_lut_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55511\,
            in1 => \N__48673\,
            in2 => \N__48661\,
            in3 => \N__48646\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17724\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17725\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_16_lut_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55496\,
            in1 => \N__48643\,
            in2 => \N__48628\,
            in3 => \N__48613\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_30\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17725\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17726\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_17_lut_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__48889\,
            in1 => \N__50734\,
            in2 => \N__55519\,
            in3 => \N__48874\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i6663_2_lut_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__56677\,
            in1 => \_gnd_net_\,
            in2 => \N__48973\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n8356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i6661_2_lut_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48969\,
            in2 => \_gnd_net_\,
            in3 => \N__56676\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i7_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__56455\,
            in1 => \_gnd_net_\,
            in2 => \N__56365\,
            in3 => \N__62725\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i9_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__60358\,
            in1 => \N__56456\,
            in2 => \_gnd_net_\,
            in3 => \N__56352\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i15_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__56454\,
            in1 => \_gnd_net_\,
            in2 => \N__56364\,
            in3 => \N__60229\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i14_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__56345\,
            in1 => \_gnd_net_\,
            in2 => \N__56480\,
            in3 => \N__60196\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i11_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__60289\,
            in1 => \N__56450\,
            in2 => \_gnd_net_\,
            in3 => \N__56344\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__48871\,
            in1 => \N__48856\,
            in2 => \N__48850\,
            in3 => \N__48823\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i10_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__60412\,
            in1 => \N__56343\,
            in2 => \_gnd_net_\,
            in3 => \N__56449\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_1_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48987\,
            in2 => \N__48991\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18144\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_2_lut_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56817\,
            in1 => \N__48952\,
            in2 => \_gnd_net_\,
            in3 => \N__48919\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18144\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18145\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_3_lut_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56821\,
            in1 => \N__48916\,
            in2 => \N__56647\,
            in3 => \N__48907\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18145\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18146\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_4_lut_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56818\,
            in1 => \N__49132\,
            in2 => \N__56626\,
            in3 => \N__48904\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18146\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18147\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_5_lut_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56822\,
            in1 => \N__51394\,
            in2 => \N__49234\,
            in3 => \N__48901\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18147\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18148\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_6_lut_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56819\,
            in1 => \N__51586\,
            in2 => \N__51376\,
            in3 => \N__48898\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18148\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18149\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_7_lut_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56823\,
            in1 => \N__60595\,
            in2 => \N__51568\,
            in3 => \N__48895\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18149\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18150\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_8_lut_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56820\,
            in1 => \N__62770\,
            in2 => \N__60574\,
            in3 => \N__48892\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_22\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18150\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18151\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_9_lut_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56813\,
            in1 => \N__65029\,
            in2 => \N__62749\,
            in3 => \N__49099\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_23\,
            ltout => OPEN,
            carryin => \bfn_19_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18152\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_10_lut_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56806\,
            in1 => \N__61006\,
            in2 => \N__66994\,
            in3 => \N__49096\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18152\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18153\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_11_lut_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56810\,
            in1 => \N__58534\,
            in2 => \N__60985\,
            in3 => \N__49093\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18153\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18154\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_12_lut_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56807\,
            in1 => \N__51811\,
            in2 => \N__58933\,
            in3 => \N__49090\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18154\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18155\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_13_lut_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56811\,
            in1 => \N__49474\,
            in2 => \N__51790\,
            in3 => \N__49087\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18155\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18156\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_14_lut_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56808\,
            in1 => \N__49267\,
            in2 => \N__49456\,
            in3 => \N__49084\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18156\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18157\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_15_lut_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56812\,
            in1 => \N__49081\,
            in2 => \N__49252\,
            in3 => \N__49069\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18157\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18158\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_16_lut_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56809\,
            in1 => \N__49066\,
            in2 => \N__49051\,
            in3 => \N__49036\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_30\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18158\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18159\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_17_lut_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56824\,
            in1 => \N__49033\,
            in2 => \N__49021\,
            in3 => \N__48994\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i17_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__56493\,
            in1 => \N__56367\,
            in2 => \_gnd_net_\,
            in3 => \N__57785\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i18_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__56494\,
            in1 => \N__56368\,
            in2 => \_gnd_net_\,
            in3 => \N__57716\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i16_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56492\,
            in1 => \N__56366\,
            in2 => \_gnd_net_\,
            in3 => \N__60259\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64862\,
            in2 => \N__64734\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n60\,
            ltout => OPEN,
            carryin => \bfn_19_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18189\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49120\,
            in2 => \N__64466\,
            in3 => \N__49114\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n106\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18189\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18190\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64111\,
            in2 => \N__51352\,
            in3 => \N__49111\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n155\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18190\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18191\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51340\,
            in2 => \N__63955\,
            in3 => \N__49108\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n204\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18191\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18192\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51331\,
            in2 => \N__63648\,
            in3 => \N__49105\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n253\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18192\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18193\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51322\,
            in2 => \N__63377\,
            in3 => \N__49102\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n302\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18193\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18194\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51313\,
            in2 => \N__63031\,
            in3 => \N__49156\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n351\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18194\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18195\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51304\,
            in2 => \N__66823\,
            in3 => \N__49153\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n400\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18195\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18196\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51295\,
            in2 => \N__66608\,
            in3 => \N__49150\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n449\,
            ltout => OPEN,
            carryin => \bfn_19_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18197\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51454\,
            in2 => \N__66294\,
            in3 => \N__49147\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n498\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18197\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18198\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51445\,
            in2 => \N__66036\,
            in3 => \N__49144\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n547\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18198\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18199\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51436\,
            in2 => \N__65776\,
            in3 => \N__49141\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n596\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18199\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18200\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51427\,
            in2 => \N__65546\,
            in3 => \N__49138\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n645\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18200\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18201\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65320\,
            in2 => \N__51418\,
            in3 => \N__49135\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n694\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18201\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18202\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65135\,
            in2 => \N__51406\,
            in3 => \N__49123\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n746\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18202\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_LUT4_0_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49237\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64863\,
            in2 => \N__64727\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n90\,
            ltout => OPEN,
            carryin => \bfn_19_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18339\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49222\,
            in2 => \N__64470\,
            in3 => \N__49216\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n136\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18339\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18340\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64182\,
            in2 => \N__49213\,
            in3 => \N__49204\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n185\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18340\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18341\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49201\,
            in2 => \N__63962\,
            in3 => \N__49195\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n234\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18341\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18342\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49192\,
            in2 => \N__63682\,
            in3 => \N__49186\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n283\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18342\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18343\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49183\,
            in2 => \N__63400\,
            in3 => \N__49177\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n332\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18343\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18344\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49174\,
            in2 => \N__63099\,
            in3 => \N__49168\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n381\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18344\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18345\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49165\,
            in2 => \N__66828\,
            in3 => \N__49159\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n430\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18345\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18346\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66612\,
            in2 => \N__49336\,
            in3 => \N__49327\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n479\,
            ltout => OPEN,
            carryin => \bfn_19_27_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18347\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49324\,
            in2 => \N__66343\,
            in3 => \N__49318\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n528\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18347\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18348\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66040\,
            in2 => \N__49315\,
            in3 => \N__49306\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n577\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18348\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18349\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49303\,
            in2 => \N__65809\,
            in3 => \N__49297\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n626\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18349\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18350\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49294\,
            in2 => \N__65581\,
            in3 => \N__49288\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n675\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18350\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18351\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49285\,
            in2 => \N__65386\,
            in3 => \N__49279\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n724\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18351\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18352\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65171\,
            in2 => \N__49276\,
            in3 => \N__49258\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n786\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18352\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_LUT4_0_LC_19_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49255\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_19_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64747\,
            in2 => \N__64955\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n87\,
            ltout => OPEN,
            carryin => \bfn_19_28_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18324\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_19_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64471\,
            in2 => \N__49432\,
            in3 => \N__49423\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n133\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18324\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18325\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_19_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49420\,
            in2 => \N__64231\,
            in3 => \N__49411\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n182\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18325\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18326\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_19_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63975\,
            in2 => \N__49408\,
            in3 => \N__49396\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n231\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18326\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18327\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_19_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49393\,
            in2 => \N__63688\,
            in3 => \N__49384\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n280\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18327\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18328\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_19_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49381\,
            in2 => \N__63389\,
            in3 => \N__49372\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n329\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18328\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18329\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_19_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49369\,
            in2 => \N__63127\,
            in3 => \N__49360\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n378\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18329\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18330\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_19_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49357\,
            in2 => \N__66880\,
            in3 => \N__49348\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n427\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18330\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18331\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_19_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49345\,
            in2 => \N__66630\,
            in3 => \N__49552\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n476\,
            ltout => OPEN,
            carryin => \bfn_19_29_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18332\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_19_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49549\,
            in2 => \N__66344\,
            in3 => \N__49540\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n525\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18332\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18333\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_19_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49537\,
            in2 => \N__66092\,
            in3 => \N__49528\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n574\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18333\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18334\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_19_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49525\,
            in2 => \N__65845\,
            in3 => \N__49516\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n623\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18334\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18335\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_19_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49513\,
            in2 => \N__65582\,
            in3 => \N__49504\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n672\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18335\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18336\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_19_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65374\,
            in2 => \N__49501\,
            in3 => \N__49486\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n721\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18336\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18337\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_19_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49483\,
            in2 => \N__65169\,
            in3 => \N__49462\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n782\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18337\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_LUT4_0_LC_19_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49459\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_20_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56121\,
            in2 => \N__53197\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n78\,
            ltout => OPEN,
            carryin => \bfn_20_5_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18122\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_20_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53161\,
            in2 => \N__49720\,
            in3 => \N__49702\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n127\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18122\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18123\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_20_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49699\,
            in2 => \N__53198\,
            in3 => \N__49681\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n176\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18123\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18124\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_20_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53165\,
            in2 => \N__49678\,
            in3 => \N__49660\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n225\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18124\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18125\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_20_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49657\,
            in2 => \N__53199\,
            in3 => \N__49642\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n274\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18125\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18126\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_20_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53169\,
            in2 => \N__49639\,
            in3 => \N__49621\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n323\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18126\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18127\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_20_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53170\,
            in2 => \N__49618\,
            in3 => \N__49597\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n372\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18127\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18128\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_20_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49594\,
            in2 => \N__53200\,
            in3 => \N__49576\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n421\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18128\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18129\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_20_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49573\,
            in2 => \N__53194\,
            in3 => \N__49555\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n470\,
            ltout => OPEN,
            carryin => \bfn_20_6_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18130\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_20_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49846\,
            in2 => \N__53196\,
            in3 => \N__49828\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n519\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18130\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18131\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_20_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49763\,
            in2 => \N__53195\,
            in3 => \N__49819\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n568\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18131\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18132\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53154\,
            in2 => \N__49770\,
            in3 => \N__49798\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n617\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18132\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n18133\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_20_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49795\,
            in2 => \N__49771\,
            in3 => \N__49747\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n774_adj_374\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n18133\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_LUT4_0_LC_20_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49744\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53611\,
            in2 => \N__53881\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n69_adj_489\,
            ltout => OPEN,
            carryin => \bfn_20_7_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17611\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49741\,
            in2 => \N__53884\,
            in3 => \N__49735\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n118_adj_487\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17611\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17612\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_20_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53832\,
            in2 => \N__49732\,
            in3 => \N__49723\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n167_adj_486\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17612\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17613\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49930\,
            in2 => \N__53885\,
            in3 => \N__49924\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n216_adj_485\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17613\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17614\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_20_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49921\,
            in2 => \N__53882\,
            in3 => \N__49915\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n265_adj_471\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17614\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17615\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49912\,
            in2 => \N__53886\,
            in3 => \N__49906\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n314\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17615\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17616\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49903\,
            in2 => \N__53883\,
            in3 => \N__49897\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n363\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17616\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17617\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49894\,
            in2 => \N__53887\,
            in3 => \N__49888\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n412_adj_482\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17617\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17618\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49885\,
            in2 => \N__53939\,
            in3 => \N__49879\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n461_adj_470\,
            ltout => OPEN,
            carryin => \bfn_20_8_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17619\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53903\,
            in2 => \N__49876\,
            in3 => \N__49867\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n510_adj_458\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17619\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17620\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49864\,
            in2 => \N__53940\,
            in3 => \N__49858\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n559\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17620\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17621\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53907\,
            in2 => \N__49855\,
            in3 => \N__49996\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n608\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17621\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17622\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49993\,
            in2 => \N__53941\,
            in3 => \N__49987\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n657\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17622\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17623\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53911\,
            in2 => \N__49984\,
            in3 => \N__49975\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n706\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17623\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17624\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49972\,
            in2 => \N__49966\,
            in3 => \N__49945\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n762_adj_402\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17624\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_LUT4_0_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49942\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54176\,
            in2 => \N__54497\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n63\,
            ltout => OPEN,
            carryin => \bfn_20_9_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17581\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51772\,
            in2 => \N__54499\,
            in3 => \N__49939\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n112_adj_442\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17581\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17582\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54445\,
            in2 => \N__51754\,
            in3 => \N__49936\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n161_adj_395\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17582\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51997\,
            in2 => \N__54500\,
            in3 => \N__49933\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n210_adj_393\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17583\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54449\,
            in2 => \N__51979\,
            in3 => \N__50023\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n259_adj_391\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17584\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54437\,
            in2 => \N__51958\,
            in3 => \N__50020\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n308\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17585\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51937\,
            in2 => \N__54498\,
            in3 => \N__50017\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n357\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17586\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17587\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54441\,
            in2 => \N__51919\,
            in3 => \N__50014\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n406\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17587\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17588\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51898\,
            in2 => \N__54509\,
            in3 => \N__50011\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n455\,
            ltout => OPEN,
            carryin => \bfn_20_10_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51880\,
            in2 => \N__54510\,
            in3 => \N__50008\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n504_adj_467\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17589\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54469\,
            in2 => \N__52174\,
            in3 => \N__50005\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n553_adj_446\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17590\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52153\,
            in2 => \N__54511\,
            in3 => \N__50002\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n602_adj_355\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17591\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54473\,
            in2 => \N__52132\,
            in3 => \N__49999\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n651\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17592\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52111\,
            in2 => \N__54512\,
            in3 => \N__50161\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n700\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17593\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50158\,
            in2 => \N__52087\,
            in3 => \N__50137\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n754_adj_405\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17594\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_LUT4_0_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50134\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60829\,
            in2 => \N__67409\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n87\,
            ltout => OPEN,
            carryin => \bfn_20_11_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17897\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50131\,
            in2 => \N__58899\,
            in3 => \N__50113\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n133_adj_388\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17897\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17898\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50110\,
            in2 => \N__54805\,
            in3 => \N__50092\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n182_adj_451\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17898\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17899\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50089\,
            in2 => \N__54534\,
            in3 => \N__50071\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n231_adj_387\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17899\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17900\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50068\,
            in2 => \N__54257\,
            in3 => \N__50050\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n280_adj_379\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17900\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17901\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53915\,
            in2 => \N__50047\,
            in3 => \N__50026\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n329_adj_439\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17901\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17902\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50317\,
            in2 => \N__53724\,
            in3 => \N__50299\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n378_adj_436\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17902\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17903\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50296\,
            in2 => \N__53369\,
            in3 => \N__50281\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n427_adj_432\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17903\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17904\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50278\,
            in2 => \N__53202\,
            in3 => \N__50260\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n476\,
            ltout => OPEN,
            carryin => \bfn_20_12_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17905\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50257\,
            in2 => \N__56214\,
            in3 => \N__50239\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n525\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17905\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17906\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50236\,
            in2 => \N__55940\,
            in3 => \N__50218\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n574\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17906\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17907\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50215\,
            in2 => \N__55718\,
            in3 => \N__50197\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n623\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17907\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17908\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50194\,
            in2 => \N__55365\,
            in3 => \N__50173\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n672\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17908\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17909\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55155\,
            in2 => \N__50170\,
            in3 => \N__50416\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n721\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17909\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17910\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54941\,
            in2 => \N__50413\,
            in3 => \N__50392\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n782\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17910\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_LUT4_0_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50389\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12703_3_lut_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55001\,
            in2 => \_gnd_net_\,
            in3 => \N__50371\,
            lcout => n794_adj_2420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51139\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_1_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61200\,
            in2 => \N__61204\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_14_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17505\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_2_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51149\,
            in2 => \_gnd_net_\,
            in3 => \N__50326\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17505\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17506\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_3_lut_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58966\,
            in2 => \N__61177\,
            in3 => \N__50323\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17506\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17507\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_4_lut_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58948\,
            in2 => \N__52546\,
            in3 => \N__50320\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17507\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17508\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_5_lut_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52324\,
            in2 => \N__52528\,
            in3 => \N__50620\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17508\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17509\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_6_lut_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50617\,
            in2 => \N__52306\,
            in3 => \N__50608\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17509\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17510\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_7_lut_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52042\,
            in2 => \N__50605\,
            in3 => \N__50593\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17510\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17511\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_8_lut_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50590\,
            in2 => \N__52024\,
            in3 => \N__50581\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17511\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17512\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_9_lut_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50578\,
            in2 => \N__50566\,
            in3 => \N__50554\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_22\,
            ltout => OPEN,
            carryin => \bfn_20_15_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17513\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_10_lut_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50551\,
            in2 => \N__50536\,
            in3 => \N__50521\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17513\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17514\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_11_lut_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50518\,
            in2 => \N__50506\,
            in3 => \N__50491\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17514\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17515\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_12_lut_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50488\,
            in2 => \N__50470\,
            in3 => \N__50455\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17515\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17516\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_13_lut_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50452\,
            in2 => \N__50851\,
            in3 => \N__50830\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17516\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17517\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_14_lut_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50827\,
            in2 => \N__50812\,
            in3 => \N__50797\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17517\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17518\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_15_lut_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50794\,
            in2 => \N__50782\,
            in3 => \N__50764\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17518\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17519\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_16_lut_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50761\,
            in2 => \N__50752\,
            in3 => \N__50737\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17519\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17520\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_17_lut_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50730\,
            in2 => \_gnd_net_\,
            in3 => \N__50716\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_269_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__50671\,
            in1 => \N__50664\,
            in2 => \N__50713\,
            in3 => \N__50626\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13205_2_lut_3_lut_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__59418\,
            in1 => \N__59295\,
            in2 => \_gnd_net_\,
            in3 => \N__51022\,
            lcout => \foc.qVoltage_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13212_2_lut_3_lut_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__59419\,
            in1 => \N__50712\,
            in2 => \_gnd_net_\,
            in3 => \N__59296\,
            lcout => \foc.qVoltage_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13215_2_lut_3_lut_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__50665\,
            in1 => \_gnd_net_\,
            in2 => \N__59440\,
            in3 => \N__59297\,
            lcout => \foc.qVoltage_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13206_2_lut_3_lut_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__51055\,
            in1 => \_gnd_net_\,
            in2 => \N__59315\,
            in3 => \N__59426\,
            lcout => OPEN,
            ltout => \foc.qVoltage_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_266_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__51061\,
            in1 => \N__51054\,
            in2 => \N__51025\,
            in3 => \N__51021\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13209_2_lut_3_lut_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__59304\,
            in1 => \N__51208\,
            in2 => \_gnd_net_\,
            in3 => \N__59427\,
            lcout => \foc.qVoltage_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i27_3_lut_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__59299\,
            in1 => \N__50983\,
            in2 => \_gnd_net_\,
            in3 => \N__59424\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_260_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011100100"
        )
    port map (
            in0 => \N__59425\,
            in1 => \N__59300\,
            in2 => \N__50959\,
            in3 => \N__52842\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13210_2_lut_3_lut_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__59305\,
            in1 => \N__50932\,
            in2 => \_gnd_net_\,
            in3 => \N__59428\,
            lcout => OPEN,
            ltout => \foc.qVoltage_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i18_2_lut_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__50931\,
            in1 => \_gnd_net_\,
            in2 => \N__50899\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i6572_2_lut_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55033\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51160\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n8265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_261_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101001110010"
        )
    port map (
            in0 => \N__59442\,
            in1 => \N__50890\,
            in2 => \N__59326\,
            in3 => \N__50881\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20586_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_265_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51235\,
            in1 => \N__51229\,
            in2 => \N__51223\,
            in3 => \N__51220\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_270_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__51214\,
            in1 => \N__51204\,
            in2 => \N__51169\,
            in3 => \N__51166\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i6570_2_lut_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__55032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51159\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i20_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56463\,
            in1 => \N__56342\,
            in2 => \_gnd_net_\,
            in3 => \N__57561\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51078\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i27_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56441\,
            in1 => \N__56308\,
            in2 => \_gnd_net_\,
            in3 => \N__57987\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i24_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__56306\,
            in1 => \N__56440\,
            in2 => \_gnd_net_\,
            in3 => \N__58170\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i29_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56442\,
            in1 => \N__56309\,
            in2 => \_gnd_net_\,
            in3 => \N__57887\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_289_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__57562\,
            in1 => \N__51274\,
            in2 => \N__57424\,
            in3 => \N__57492\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20664_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_290_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__58171\,
            in1 => \N__58240\,
            in2 => \N__51265\,
            in3 => \N__58111\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i790_4_lut_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__57988\,
            in1 => \N__57940\,
            in2 => \N__51262\,
            in3 => \N__58042\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_293_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__58487\,
            in1 => \N__57888\,
            in2 => \N__51259\,
            in3 => \N__58369\,
            lcout => \Saturate_out1_31__N_266_adj_2417\,
            ltout => \Saturate_out1_31__N_266_adj_2417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i26_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__56307\,
            in1 => \_gnd_net_\,
            in2 => \N__51256\,
            in3 => \N__58041\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i21_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__56458\,
            in1 => \N__56298\,
            in2 => \_gnd_net_\,
            in3 => \N__57493\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i19_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__57640\,
            in1 => \N__56297\,
            in2 => \_gnd_net_\,
            in3 => \N__56457\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i2_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__56460\,
            in1 => \N__60076\,
            in2 => \_gnd_net_\,
            in3 => \N__56300\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i62_4_lut_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51253\,
            in1 => \N__59122\,
            in2 => \N__52957\,
            in3 => \N__51244\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_283_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__58368\,
            in1 => \N__58489\,
            in2 => \N__57889\,
            in3 => \N__56608\,
            lcout => \Saturate_out1_31__N_267_adj_2418\,
            ltout => \Saturate_out1_31__N_267_adj_2418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i6_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__62671\,
            in1 => \_gnd_net_\,
            in2 => \N__51286\,
            in3 => \N__56462\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i30_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56461\,
            in1 => \N__56301\,
            in2 => \_gnd_net_\,
            in3 => \N__58488\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i23_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__56299\,
            in1 => \N__58239\,
            in2 => \_gnd_net_\,
            in3 => \N__56459\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i12_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__56481\,
            in1 => \N__56302\,
            in2 => \_gnd_net_\,
            in3 => \N__60327\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i4_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__56304\,
            in1 => \N__60112\,
            in2 => \_gnd_net_\,
            in3 => \N__56483\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i772_4_lut_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__62647\,
            in1 => \N__60411\,
            in2 => \N__60354\,
            in3 => \N__60382\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n22_adj_762_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_286_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__60328\,
            in1 => \N__60310\,
            in2 => \N__51283\,
            in3 => \N__60285\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20694_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_287_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__60222\,
            in1 => \N__60189\,
            in2 => \N__51280\,
            in3 => \N__60258\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_288_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__57786\,
            in1 => \N__57639\,
            in2 => \N__51277\,
            in3 => \N__57717\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i8_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56484\,
            in1 => \N__56305\,
            in2 => \_gnd_net_\,
            in3 => \N__60381\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i13_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__56303\,
            in1 => \N__60309\,
            in2 => \_gnd_net_\,
            in3 => \N__56482\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64712\,
            in2 => \N__64887\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n63\,
            ltout => OPEN,
            carryin => \bfn_20_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18204\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64454\,
            in2 => \N__51361\,
            in3 => \N__51343\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n109\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18204\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18205\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51544\,
            in2 => \N__64178\,
            in3 => \N__51334\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n158\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18205\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18206\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51532\,
            in2 => \N__63888\,
            in3 => \N__51325\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n207\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18206\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18207\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51520\,
            in2 => \N__63631\,
            in3 => \N__51316\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n256\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18207\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18208\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51508\,
            in2 => \N__63378\,
            in3 => \N__51307\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n305\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18208\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18209\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62938\,
            in2 => \N__51496\,
            in3 => \N__51298\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n354\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18209\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18210\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66760\,
            in2 => \N__51481\,
            in3 => \N__51457\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n403\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18210\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18211\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51466\,
            in2 => \N__66599\,
            in3 => \N__51448\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n452\,
            ltout => OPEN,
            carryin => \bfn_20_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18212\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51670\,
            in2 => \N__66286\,
            in3 => \N__51439\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n501\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18212\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18213\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51658\,
            in2 => \N__66091\,
            in3 => \N__51430\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n550\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18213\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18214\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51646\,
            in2 => \N__65830\,
            in3 => \N__51421\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n599\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18214\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18215\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65595\,
            in2 => \N__51634\,
            in3 => \N__51409\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n648\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18215\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18216\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65348\,
            in2 => \N__51619\,
            in3 => \N__51397\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n697\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18216\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18217\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65139\,
            in2 => \N__51601\,
            in3 => \N__51382\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n750\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18217\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_LUT4_0_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51379\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64713\,
            in2 => \N__64900\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n66\,
            ltout => OPEN,
            carryin => \bfn_20_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18219\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64478\,
            in2 => \N__51553\,
            in3 => \N__51535\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n112\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18219\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18220\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60544\,
            in2 => \N__64230\,
            in3 => \N__51523\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n161\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18220\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18221\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60532\,
            in2 => \N__63963\,
            in3 => \N__51511\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n210\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18221\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18222\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60520\,
            in2 => \N__63647\,
            in3 => \N__51499\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n259\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18222\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18223\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60508\,
            in2 => \N__63382\,
            in3 => \N__51484\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n308\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18223\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18224\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63093\,
            in2 => \N__60496\,
            in3 => \N__51469\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n357\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18224\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18225\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66782\,
            in2 => \N__60481\,
            in3 => \N__51460\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n406\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18225\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18226\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_20_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60466\,
            in2 => \N__66600\,
            in3 => \N__51661\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n455\,
            ltout => OPEN,
            carryin => \bfn_20_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18227\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_20_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60673\,
            in2 => \N__66348\,
            in3 => \N__51649\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n504\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18227\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18228\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_20_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60661\,
            in2 => \N__66070\,
            in3 => \N__51637\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n553\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18228\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18229\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_20_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60649\,
            in2 => \N__65839\,
            in3 => \N__51622\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n602\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18229\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18230\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_20_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60637\,
            in2 => \N__65600\,
            in3 => \N__51604\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n651\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18230\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18231\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_20_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65352\,
            in2 => \N__60625\,
            in3 => \N__51589\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n700\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18231\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18232\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_20_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65170\,
            in2 => \N__60610\,
            in3 => \N__51574\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n754\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18232\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_LUT4_0_LC_20_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51571\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_20_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64888\,
            in2 => \N__64748\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n84\,
            ltout => OPEN,
            carryin => \bfn_20_28_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18309\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_20_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51742\,
            in2 => \N__64488\,
            in3 => \N__51736\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n130\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18309\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18310\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_20_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51733\,
            in2 => \N__64232\,
            in3 => \N__51727\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n179\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18310\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18311\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_20_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51724\,
            in2 => \N__63982\,
            in3 => \N__51718\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n228\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18311\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18312\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_20_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51715\,
            in2 => \N__63655\,
            in3 => \N__51709\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n277\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18312\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18313\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_20_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51706\,
            in2 => \N__63385\,
            in3 => \N__51700\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n326_adj_588\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18313\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18314\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_20_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51697\,
            in2 => \N__63095\,
            in3 => \N__51691\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n375_adj_587\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18314\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18315\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_20_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51688\,
            in2 => \N__66921\,
            in3 => \N__51682\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n424_adj_586\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18315\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18316\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_20_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51679\,
            in2 => \N__66625\,
            in3 => \N__51673\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n473_adj_585\,
            ltout => OPEN,
            carryin => \bfn_20_29_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18317\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_20_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51868\,
            in2 => \N__66346\,
            in3 => \N__51862\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n522_adj_584\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18317\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18318\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_20_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51859\,
            in2 => \N__66093\,
            in3 => \N__51853\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n571\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18318\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18319\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_20_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51850\,
            in2 => \N__65831\,
            in3 => \N__51844\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n620\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18319\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18320\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_20_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51841\,
            in2 => \N__65601\,
            in3 => \N__51835\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n669\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18320\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18321\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_20_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65361\,
            in2 => \N__51832\,
            in3 => \N__51823\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n718\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18321\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18322\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_20_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65192\,
            in2 => \N__51820\,
            in3 => \N__51796\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n778\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18322\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_LUT4_0_LC_20_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51793\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_21_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53888\,
            in2 => \N__54135\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n66\,
            ltout => OPEN,
            carryin => \bfn_21_7_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17596\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_21_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54084\,
            in2 => \N__51763\,
            in3 => \N__52009\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n115_adj_488\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17596\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17597\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_21_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54138\,
            in2 => \N__52006\,
            in3 => \N__51988\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n164_adj_466\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17597\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17598\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_21_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51985\,
            in2 => \N__54193\,
            in3 => \N__51967\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n213_adj_445\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17598\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17599\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_21_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51964\,
            in2 => \N__54136\,
            in3 => \N__51946\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n262\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17599\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17600\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_21_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51943\,
            in2 => \N__54194\,
            in3 => \N__51928\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n311\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17600\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17601\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_21_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51925\,
            in2 => \N__54137\,
            in3 => \N__51907\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n360_adj_484\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17601\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17602\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_21_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51904\,
            in2 => \N__54195\,
            in3 => \N__51889\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n409_adj_483\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17602\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17603\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_21_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51886\,
            in2 => \N__54252\,
            in3 => \N__51871\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n458_adj_468\,
            ltout => OPEN,
            carryin => \bfn_21_8_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17604\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54224\,
            in2 => \N__52183\,
            in3 => \N__52162\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n507_adj_447\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17604\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17605\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_21_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52159\,
            in2 => \N__54253\,
            in3 => \N__52144\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n556\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17605\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17606\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54228\,
            in2 => \N__52141\,
            in3 => \N__52120\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n605\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17606\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17607\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_21_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52117\,
            in2 => \N__54254\,
            in3 => \N__52099\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n654\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17607\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17608\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_21_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54232\,
            in2 => \N__52096\,
            in3 => \N__52072\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n703\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17608\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17609\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_21_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52069\,
            in2 => \N__52051\,
            in3 => \N__52030\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n758_adj_403\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17609\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_LUT4_0_LC_21_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52027\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54450\,
            in2 => \N__54796\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n60_adj_495\,
            ltout => OPEN,
            carryin => \bfn_21_9_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17566\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54750\,
            in2 => \N__52276\,
            in3 => \N__52267\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n109\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17566\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17567\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52264\,
            in2 => \N__54797\,
            in3 => \N__52258\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n158\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17567\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17568\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52255\,
            in2 => \N__54800\,
            in3 => \N__52249\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n207_adj_394\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17568\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17569\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52246\,
            in2 => \N__54798\,
            in3 => \N__52240\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n256_adj_392\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17569\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17570\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54757\,
            in2 => \N__52237\,
            in3 => \N__52228\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n305_adj_390\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17570\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17571\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52225\,
            in2 => \N__54799\,
            in3 => \N__52219\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n354\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17571\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17572\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54761\,
            in2 => \N__52216\,
            in3 => \N__52207\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n403\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17572\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17573\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52204\,
            in2 => \N__54768\,
            in3 => \N__52198\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n452\,
            ltout => OPEN,
            carryin => \bfn_21_10_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17574\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54705\,
            in2 => \N__52195\,
            in3 => \N__52186\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n501_adj_481\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17574\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17575\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52393\,
            in2 => \N__54769\,
            in3 => \N__52387\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n550_adj_441\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17575\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17576\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54709\,
            in2 => \N__52384\,
            in3 => \N__52375\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n599_adj_376\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17576\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17577\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52372\,
            in2 => \N__54770\,
            in3 => \N__52366\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n648\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17577\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17578\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54713\,
            in2 => \N__52363\,
            in3 => \N__52354\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n697_adj_444\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17578\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17579\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52351\,
            in2 => \N__52333\,
            in3 => \N__52312\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n750_adj_407\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17579\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_LUT4_0_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52309\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54801\,
            in2 => \N__58900\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n57_adj_491\,
            ltout => OPEN,
            carryin => \bfn_21_11_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17551\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58852\,
            in2 => \N__52291\,
            in3 => \N__52279\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n106_adj_509\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17551\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17552\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52510\,
            in2 => \N__58901\,
            in3 => \N__52501\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n155\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17552\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17553\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58856\,
            in2 => \N__52498\,
            in3 => \N__52486\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n204\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17553\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17554\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52483\,
            in2 => \N__58902\,
            in3 => \N__52474\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n253_adj_464\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17554\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17555\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58860\,
            in2 => \N__52471\,
            in3 => \N__52459\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n302\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17555\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17556\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52456\,
            in2 => \N__58903\,
            in3 => \N__52447\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n351_adj_396\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17556\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17557\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58864\,
            in2 => \N__52444\,
            in3 => \N__52432\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n400\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17557\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17558\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52429\,
            in2 => \N__58909\,
            in3 => \N__52420\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n449\,
            ltout => OPEN,
            carryin => \bfn_21_12_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17559\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58887\,
            in2 => \N__52417\,
            in3 => \N__52405\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n498\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17559\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17560\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52402\,
            in2 => \N__58910\,
            in3 => \N__52624\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n547\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17560\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17561\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58891\,
            in2 => \N__52621\,
            in3 => \N__52609\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n596\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17561\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17562\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52606\,
            in2 => \N__58911\,
            in3 => \N__52597\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n645\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17562\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17563\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58895\,
            in2 => \N__52594\,
            in3 => \N__52582\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n694\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17563\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17564\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52579\,
            in2 => \N__52558\,
            in3 => \N__52534\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n746_adj_409\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17564\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_LUT4_0_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52531\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13161_2_lut_3_lut_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__61389\,
            in1 => \N__67618\,
            in2 => \_gnd_net_\,
            in3 => \N__61454\,
            lcout => OPEN,
            ltout => \foc.dVoltage_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_119_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__67617\,
            in1 => \N__67978\,
            in2 => \N__52513\,
            in3 => \N__59071\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13174_2_lut_3_lut_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__68608\,
            in1 => \_gnd_net_\,
            in2 => \N__61479\,
            in3 => \N__61377\,
            lcout => \foc.dVoltage_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13168_2_lut_3_lut_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__61375\,
            in1 => \N__67899\,
            in2 => \_gnd_net_\,
            in3 => \N__61462\,
            lcout => \foc.dVoltage_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13169_2_lut_3_lut_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__68944\,
            in1 => \_gnd_net_\,
            in2 => \N__61478\,
            in3 => \N__61376\,
            lcout => \foc.dVoltage_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_118_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011100010"
        )
    port map (
            in0 => \N__61374\,
            in1 => \N__61461\,
            in2 => \N__68557\,
            in3 => \N__69208\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20548_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_121_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__68607\,
            in1 => \N__59104\,
            in2 => \N__52678\,
            in3 => \N__52675\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_124_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__59080\,
            in1 => \N__68943\,
            in2 => \N__52669\,
            in3 => \N__52666\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_127_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__59218\,
            in1 => \N__61501\,
            in2 => \N__52660\,
            in3 => \N__59203\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i62_4_lut_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001101"
        )
    port map (
            in0 => \N__61373\,
            in1 => \N__61306\,
            in2 => \N__52657\,
            in3 => \N__61460\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13207_2_lut_3_lut_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__52651\,
            in1 => \N__59298\,
            in2 => \_gnd_net_\,
            in3 => \N__59423\,
            lcout => OPEN,
            ltout => \foc.qVoltage_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111010"
        )
    port map (
            in0 => \N__52909\,
            in1 => \_gnd_net_\,
            in2 => \N__52654\,
            in3 => \N__52650\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_267_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__52684\,
            in1 => \N__52726\,
            in2 => \N__52960\,
            in3 => \N__59161\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_262_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001001100"
        )
    port map (
            in0 => \N__52874\,
            in1 => \N__59292\,
            in2 => \N__52942\,
            in3 => \N__59415\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1223_rep_3_4_lut_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__52903\,
            in1 => \N__52875\,
            in2 => \N__52857\,
            in3 => \N__52824\,
            lcout => \foc.Out_31__N_333\,
            ltout => \foc.Out_31__N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13211_2_lut_3_lut_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__52795\,
            in1 => \_gnd_net_\,
            in2 => \N__52891\,
            in3 => \N__59416\,
            lcout => \foc.qVoltage_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i12830_4_lut_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__52888\,
            in1 => \N__52876\,
            in2 => \N__52858\,
            in3 => \N__52825\,
            lcout => \foc.Out_31__N_332\,
            ltout => \foc.Out_31__N_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13216_2_lut_3_lut_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__52756\,
            in1 => \_gnd_net_\,
            in2 => \N__52804\,
            in3 => \N__59293\,
            lcout => OPEN,
            ltout => \foc.qVoltage_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_264_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__52801\,
            in1 => \N__52794\,
            in2 => \N__52759\,
            in3 => \N__52755\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13217_2_lut_3_lut_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__52722\,
            in1 => \N__59294\,
            in2 => \_gnd_net_\,
            in3 => \N__59417\,
            lcout => \foc.qVoltage_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60902\,
            in2 => \N__67467\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n57\,
            ltout => OPEN,
            carryin => \bfn_21_17_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55444\,
            in1 => \N__54826\,
            in2 => \N__58915\,
            in3 => \N__54820\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_4\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17736\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17737\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55448\,
            in1 => \N__54817\,
            in2 => \N__54568\,
            in3 => \N__54553\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_5\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17737\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17738\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55445\,
            in1 => \N__54550\,
            in2 => \N__54538\,
            in3 => \N__54286\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_6\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17738\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55449\,
            in1 => \N__54283\,
            in2 => \N__54271\,
            in3 => \N__54016\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_7\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17739\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55446\,
            in1 => \N__54013\,
            in2 => \N__53999\,
            in3 => \N__53743\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_8\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17740\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55450\,
            in1 => \N__53740\,
            in2 => \N__53723\,
            in3 => \N__53494\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_9\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17741\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55447\,
            in1 => \N__53491\,
            in2 => \N__53478\,
            in3 => \N__53227\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_10\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17742\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55451\,
            in1 => \N__53224\,
            in2 => \N__53136\,
            in3 => \N__52963\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_11\,
            ltout => OPEN,
            carryin => \bfn_21_18_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55454\,
            in1 => \N__56227\,
            in2 => \N__56215\,
            in3 => \N__55981\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_12\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17744\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55452\,
            in1 => \N__55978\,
            in2 => \N__55964\,
            in3 => \N__55753\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17745\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55455\,
            in1 => \N__55750\,
            in2 => \N__55737\,
            in3 => \N__55522\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_14\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17746\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__55453\,
            in1 => \N__55390\,
            in2 => \N__55377\,
            in3 => \N__55189\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17747\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55179\,
            in2 => \N__55048\,
            in3 => \N__55024\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n691\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17748\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55021\,
            in2 => \N__55009\,
            in3 => \N__54847\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n742\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17749\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_LUT4_0_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54844\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i5_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__56478\,
            in1 => \N__56363\,
            in2 => \_gnd_net_\,
            in3 => \N__62697\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i1_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__56361\,
            in1 => \N__56476\,
            in2 => \_gnd_net_\,
            in3 => \N__60151\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i3_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__56477\,
            in1 => \N__56362\,
            in2 => \_gnd_net_\,
            in3 => \N__60097\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i22_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__56330\,
            in1 => \_gnd_net_\,
            in2 => \N__56479\,
            in3 => \N__57419\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i0_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__60127\,
            in1 => \N__56329\,
            in2 => \_gnd_net_\,
            in3 => \N__56443\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i28_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__56448\,
            in1 => \_gnd_net_\,
            in2 => \N__56360\,
            in3 => \N__57938\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i25_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__58109\,
            in1 => \N__56447\,
            in2 => \_gnd_net_\,
            in3 => \N__56331\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_280_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__57635\,
            in1 => \N__57787\,
            in2 => \N__57718\,
            in3 => \N__60163\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_281_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__57420\,
            in1 => \N__57491\,
            in2 => \N__56233\,
            in3 => \N__57551\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_282_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__58169\,
            in1 => \N__58110\,
            in2 => \N__56230\,
            in3 => \N__58238\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i14382_4_lut_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__58040\,
            in1 => \N__57939\,
            in2 => \N__56611\,
            in3 => \N__57986\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64632\,
            in2 => \N__64844\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n57\,
            ltout => OPEN,
            carryin => \bfn_21_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18174\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56778\,
            in1 => \N__56602\,
            in2 => \N__64489\,
            in3 => \N__56596\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_4\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18174\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18175\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56782\,
            in1 => \N__64101\,
            in2 => \N__56593\,
            in3 => \N__56575\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_5\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18175\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18176\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56779\,
            in1 => \N__56572\,
            in2 => \N__63936\,
            in3 => \N__56560\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_6\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18176\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18177\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56783\,
            in1 => \N__56557\,
            in2 => \N__63609\,
            in3 => \N__56545\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_7\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18177\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18178\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56780\,
            in1 => \N__56542\,
            in2 => \N__63399\,
            in3 => \N__56530\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_8\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18178\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18179\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56784\,
            in1 => \N__56527\,
            in2 => \N__63065\,
            in3 => \N__56512\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_9\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18179\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18180\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56781\,
            in1 => \N__56509\,
            in2 => \N__66875\,
            in3 => \N__56497\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_10\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18180\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18181\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56801\,
            in1 => \N__56884\,
            in2 => \N__66521\,
            in3 => \N__56872\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_11\,
            ltout => OPEN,
            carryin => \bfn_21_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18182\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56804\,
            in1 => \N__56869\,
            in2 => \N__66261\,
            in3 => \N__56857\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_12\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18182\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18183\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56802\,
            in1 => \N__56854\,
            in2 => \N__66012\,
            in3 => \N__56842\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18183\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18184\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56805\,
            in1 => \N__56839\,
            in2 => \N__65791\,
            in3 => \N__56827\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_14\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18184\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18185\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__56803\,
            in1 => \N__56707\,
            in2 => \N__65570\,
            in3 => \N__56695\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18185\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18186\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65342\,
            in2 => \N__56692\,
            in3 => \N__56662\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n691\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18186\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18187\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56659\,
            in2 => \N__65178\,
            in3 => \N__56632\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n742\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18187\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_LUT4_0_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56629\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_2_lut_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57082\,
            in2 => \N__57073\,
            in3 => \_gnd_net_\,
            lcout => \Add_add_temp_4_adj_2416\,
            ltout => OPEN,
            carryin => \bfn_21_23_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15913\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_3_lut_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57061\,
            in2 => \N__57052\,
            in3 => \N__57040\,
            lcout => \Add_add_temp_5_adj_2415\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15913\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15914\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_4_lut_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57037\,
            in2 => \N__57028\,
            in3 => \N__57013\,
            lcout => \Add_add_temp_6_adj_2414\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15914\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15915\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_5_lut_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57010\,
            in2 => \N__57001\,
            in3 => \N__56989\,
            lcout => \Add_add_temp_7_adj_2413\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15915\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15916\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_6_lut_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56986\,
            in2 => \N__56980\,
            in3 => \N__56968\,
            lcout => \Add_add_temp_8_adj_2412\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15916\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15917\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_7_lut_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56965\,
            in2 => \N__56956\,
            in3 => \N__56944\,
            lcout => \Add_add_temp_9_adj_2411\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15917\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15918\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_8_lut_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56941\,
            in2 => \N__56932\,
            in3 => \N__56920\,
            lcout => \Add_add_temp_10_adj_2410\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15918\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15919\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_9_lut_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56917\,
            in2 => \N__56896\,
            in3 => \N__56887\,
            lcout => \Add_add_temp_11_adj_2409\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15919\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15920\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_10_lut_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57385\,
            in2 => \N__57367\,
            in3 => \N__57352\,
            lcout => \Add_add_temp_12_adj_2408\,
            ltout => OPEN,
            carryin => \bfn_21_24_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15921\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_11_lut_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57349\,
            in2 => \N__57340\,
            in3 => \N__57316\,
            lcout => \Add_add_temp_13_adj_2407\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15921\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15922\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_12_lut_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57313\,
            in2 => \N__57304\,
            in3 => \N__57280\,
            lcout => \Add_add_temp_14_adj_2406\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15922\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15923\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_13_lut_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57277\,
            in2 => \N__57253\,
            in3 => \N__57238\,
            lcout => \Add_add_temp_15_adj_2405\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15923\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15924\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_14_lut_LC_21_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57235\,
            in2 => \N__57223\,
            in3 => \N__57202\,
            lcout => \Add_add_temp_16_adj_2404\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15924\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15925\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_15_lut_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57199\,
            in2 => \N__57178\,
            in3 => \N__57163\,
            lcout => \Add_add_temp_17_adj_2403\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15925\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15926\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_16_lut_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57160\,
            in2 => \N__57136\,
            in3 => \N__57121\,
            lcout => \Add_add_temp_18_adj_2402\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15926\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15927\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_17_lut_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57118\,
            in2 => \N__57097\,
            in3 => \N__57862\,
            lcout => \Add_add_temp_19_adj_2401\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15927\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15928\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_18_lut_LC_21_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57859\,
            in2 => \N__57841\,
            in3 => \N__57823\,
            lcout => \Add_add_temp_20_adj_2400\,
            ltout => OPEN,
            carryin => \bfn_21_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15929\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_19_lut_LC_21_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57820\,
            in2 => \N__57802\,
            in3 => \N__57754\,
            lcout => \Add_add_temp_21_adj_2399\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15929\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15930\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_20_lut_LC_21_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57751\,
            in2 => \N__57733\,
            in3 => \N__57688\,
            lcout => \Add_add_temp_22_adj_2398\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15930\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15931\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_21_lut_LC_21_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57685\,
            in2 => \N__57658\,
            in3 => \N__57604\,
            lcout => \Add_add_temp_23_adj_2397\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15931\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15932\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_22_lut_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57601\,
            in2 => \N__57577\,
            in3 => \N__57532\,
            lcout => \Add_add_temp_24_adj_2396\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15932\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15933\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_23_lut_LC_21_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57529\,
            in2 => \N__57508\,
            in3 => \N__57466\,
            lcout => \Add_add_temp_25_adj_2395\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15933\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15934\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_24_lut_LC_21_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57456\,
            in2 => \N__57439\,
            in3 => \N__57388\,
            lcout => \Add_add_temp_26_adj_2394\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15934\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15935\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_25_lut_LC_21_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58279\,
            in2 => \N__58255\,
            in3 => \N__58216\,
            lcout => \Add_add_temp_27_adj_2393\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15935\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15936\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_26_lut_LC_21_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58212\,
            in2 => \N__58186\,
            in3 => \N__58150\,
            lcout => \Add_add_temp_28_adj_2392\,
            ltout => OPEN,
            carryin => \bfn_21_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15937\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_27_lut_LC_21_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58140\,
            in2 => \N__58126\,
            in3 => \N__58084\,
            lcout => \Add_add_temp_29_adj_2391\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15937\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15938\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_28_lut_LC_21_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58081\,
            in2 => \N__58057\,
            in3 => \N__58018\,
            lcout => \Add_add_temp_30_adj_2390\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15938\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15939\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_29_lut_LC_21_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58015\,
            in2 => \N__58403\,
            in3 => \N__57967\,
            lcout => \Add_add_temp_31_adj_2389\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15939\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15940\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_30_lut_LC_21_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58395\,
            in2 => \N__57963\,
            in3 => \N__57916\,
            lcout => \Add_add_temp_32_adj_2388\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15940\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15941\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_31_lut_LC_21_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57913\,
            in2 => \N__58404\,
            in3 => \N__57865\,
            lcout => \Add_add_temp_33_adj_2387\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15941\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15942\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_32_lut_LC_21_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58399\,
            in2 => \N__58519\,
            in3 => \N__58459\,
            lcout => \Add_add_temp_34_adj_2386\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15942\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15943\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_33_lut_LC_21_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__58456\,
            in1 => \_gnd_net_\,
            in2 => \N__58405\,
            in3 => \N__58372\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_21_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64899\,
            in2 => \N__64749\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n81\,
            ltout => OPEN,
            carryin => \bfn_21_28_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18294\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_21_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58339\,
            in2 => \N__64497\,
            in3 => \N__58333\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n127\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18294\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18295\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_21_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58330\,
            in2 => \N__64236\,
            in3 => \N__58324\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n176\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18295\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18296\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_21_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58321\,
            in2 => \N__63981\,
            in3 => \N__58315\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n225\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18296\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18297\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_21_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63630\,
            in2 => \N__58312\,
            in3 => \N__58303\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n274\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18297\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18298\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_21_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58300\,
            in2 => \N__63401\,
            in3 => \N__58294\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n323\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18298\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18299\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_21_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63094\,
            in2 => \N__58291\,
            in3 => \N__58282\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n372_adj_596\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18299\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18300\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_21_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66884\,
            in2 => \N__58615\,
            in3 => \N__58606\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n421_adj_595\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18300\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18301\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_21_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66638\,
            in2 => \N__58603\,
            in3 => \N__58594\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n470_adj_594\,
            ltout => OPEN,
            carryin => \bfn_21_29_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18302\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_21_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58591\,
            in2 => \N__66347\,
            in3 => \N__58585\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n519_adj_593\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18302\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18303\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_21_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58582\,
            in2 => \N__66094\,
            in3 => \N__58576\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n568_adj_592\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18303\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18304\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_21_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58573\,
            in2 => \N__65832\,
            in3 => \N__58567\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n617_adj_591\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18304\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18305\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_21_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58564\,
            in2 => \N__65602\,
            in3 => \N__58558\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n666\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18305\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18306\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_21_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65387\,
            in2 => \N__58555\,
            in3 => \N__58546\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n715\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18306\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18307\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_21_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65203\,
            in2 => \N__58543\,
            in3 => \N__58522\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n774_adj_589\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18307\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_LUT4_0_LC_21_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58936\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58865\,
            in2 => \N__60951\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n54\,
            ltout => OPEN,
            carryin => \bfn_22_11_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17536\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60914\,
            in2 => \N__58687\,
            in3 => \N__58678\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n103\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17536\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17537\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58675\,
            in2 => \N__60952\,
            in3 => \N__58669\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n152\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17537\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17538\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60918\,
            in2 => \N__58666\,
            in3 => \N__58657\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n201\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17538\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17539\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58654\,
            in2 => \N__60953\,
            in3 => \N__58648\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n250\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17539\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17540\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60922\,
            in2 => \N__58645\,
            in3 => \N__58636\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n299\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17540\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17541\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58633\,
            in2 => \N__60954\,
            in3 => \N__58627\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n348\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17541\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17542\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60926\,
            in2 => \N__58624\,
            in3 => \N__59065\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n397\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17542\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17543\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59062\,
            in2 => \N__60955\,
            in3 => \N__59056\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n446\,
            ltout => OPEN,
            carryin => \bfn_22_12_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17544\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60930\,
            in2 => \N__59053\,
            in3 => \N__59044\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n495\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17544\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17545\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59041\,
            in2 => \N__60956\,
            in3 => \N__59035\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n544\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17545\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17546\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60934\,
            in2 => \N__59032\,
            in3 => \N__59023\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n593\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17546\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17547\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59020\,
            in2 => \N__60957\,
            in3 => \N__59014\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n642\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17547\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17548\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60938\,
            in2 => \N__59011\,
            in3 => \N__59002\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n691_adj_440\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17548\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17549\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58999\,
            in2 => \N__58993\,
            in3 => \N__58954\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n742_adj_411\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17549\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_LUT4_0_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58951\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_117_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010101100"
        )
    port map (
            in0 => \N__69156\,
            in1 => \N__61378\,
            in2 => \N__61475\,
            in3 => \N__69108\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__59107\,
            in3 => \N__61156\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13171_2_lut_3_lut_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__61450\,
            in1 => \N__61381\,
            in2 => \_gnd_net_\,
            in3 => \N__68800\,
            lcout => \foc.dVoltage_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13164_2_lut_3_lut_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__61379\,
            in1 => \N__61449\,
            in2 => \_gnd_net_\,
            in3 => \N__68188\,
            lcout => OPEN,
            ltout => \foc.dVoltage_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i15_2_lut_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__59098\,
            in3 => \N__68187\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_120_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__68799\,
            in1 => \N__59095\,
            in2 => \N__59089\,
            in3 => \N__59086\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12820_4_lut_LC_22_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__69157\,
            in1 => \N__69109\,
            in2 => \N__69010\,
            in3 => \N__61162\,
            lcout => \foc.Out_31__N_332_adj_2312\,
            ltout => \foc.Out_31__N_332_adj_2312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13167_2_lut_3_lut_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__61380\,
            in1 => \_gnd_net_\,
            in2 => \N__59074\,
            in3 => \N__67977\,
            lcout => \foc.dVoltage_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1212_rep_6_4_lut_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__61294\,
            in1 => \N__61312\,
            in2 => \N__69006\,
            in3 => \N__69107\,
            lcout => \foc.Out_31__N_333_adj_2310\,
            ltout => \foc.Out_31__N_333_adj_2310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13173_2_lut_3_lut_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68659\,
            in2 => \N__59230\,
            in3 => \N__61459\,
            lcout => \foc.dVoltage_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13162_2_lut_3_lut_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__67555\,
            in1 => \N__61477\,
            in2 => \_gnd_net_\,
            in3 => \N__61371\,
            lcout => OPEN,
            ltout => \foc.dVoltage_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_126_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__59227\,
            in1 => \N__68658\,
            in2 => \N__59221\,
            in3 => \N__67554\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13170_2_lut_3_lut_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__61458\,
            in1 => \N__68872\,
            in2 => \_gnd_net_\,
            in3 => \N__61372\,
            lcout => OPEN,
            ltout => \foc.dVoltage_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_123_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__68871\,
            in1 => \N__67898\,
            in2 => \N__59212\,
            in3 => \N__59209\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13204_2_lut_3_lut_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__59197\,
            in1 => \N__59325\,
            in2 => \_gnd_net_\,
            in3 => \N__59443\,
            lcout => OPEN,
            ltout => \foc.qVoltage_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_263_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__59359\,
            in1 => \N__59196\,
            in2 => \N__59164\,
            in3 => \N__59239\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.equal_13244_i21_2_lut_3_lut_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000100010"
        )
    port map (
            in0 => \N__59429\,
            in1 => \N__59155\,
            in2 => \_gnd_net_\,
            in3 => \N__59306\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_268_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__59449\,
            in1 => \N__59481\,
            in2 => \N__59131\,
            in3 => \N__59128\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13208_2_lut_3_lut_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__59482\,
            in1 => \_gnd_net_\,
            in2 => \N__59441\,
            in3 => \N__59307\,
            lcout => \foc.qVoltage_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13214_2_lut_3_lut_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__59433\,
            in1 => \N__59358\,
            in2 => \_gnd_net_\,
            in3 => \N__59308\,
            lcout => \foc.qVoltage_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i30_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__61974\,
            in1 => \N__61629\,
            in2 => \_gnd_net_\,
            in3 => \N__61910\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i0_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__61907\,
            in1 => \N__61971\,
            in2 => \_gnd_net_\,
            in3 => \N__62551\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i27_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__61972\,
            in1 => \N__61908\,
            in2 => \_gnd_net_\,
            in3 => \N__61712\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i29_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__61973\,
            in1 => \N__61909\,
            in2 => \_gnd_net_\,
            in3 => \N__61597\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i6_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__61906\,
            in1 => \N__61970\,
            in2 => \_gnd_net_\,
            in3 => \N__62416\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i13327_4_lut_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__59614\,
            in1 => \N__61685\,
            in2 => \N__61716\,
            in3 => \N__61655\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_139_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__61592\,
            in1 => \N__62142\,
            in2 => \N__59233\,
            in3 => \N__61622\,
            lcout => \Saturate_out1_31__N_267\,
            ltout => \Saturate_out1_31__N_267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i18_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__62175\,
            in1 => \_gnd_net_\,
            in2 => \N__59491\,
            in3 => \N__61901\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i1_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__61902\,
            in1 => \N__62569\,
            in2 => \_gnd_net_\,
            in3 => \N__61966\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i3_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__61969\,
            in1 => \N__61905\,
            in2 => \_gnd_net_\,
            in3 => \N__62518\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i2_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__61904\,
            in1 => \N__61968\,
            in2 => \_gnd_net_\,
            in3 => \N__62490\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i20_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__61967\,
            in1 => \N__61903\,
            in2 => \_gnd_net_\,
            in3 => \N__59791\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i24_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__61911\,
            in1 => \N__61985\,
            in2 => \_gnd_net_\,
            in3 => \N__60005\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i25_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__61986\,
            in1 => \N__61912\,
            in2 => \_gnd_net_\,
            in3 => \N__59972\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_143_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__62307\,
            in1 => \N__62250\,
            in2 => \N__62284\,
            in3 => \N__61789\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19842_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_144_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__62226\,
            in1 => \N__62202\,
            in2 => \N__59488\,
            in3 => \N__62176\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_145_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__61551\,
            in1 => \N__62060\,
            in2 => \N__59485\,
            in3 => \N__59787\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_146_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__60007\,
            in1 => \N__59974\,
            in2 => \N__59620\,
            in3 => \N__61530\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_137_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__61550\,
            in1 => \N__62152\,
            in2 => \N__62064\,
            in3 => \N__59786\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20648_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_138_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__60006\,
            in1 => \N__59973\,
            in2 => \N__59617\,
            in3 => \N__61529\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_2_lut_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59608\,
            in2 => \N__59599\,
            in3 => \_gnd_net_\,
            lcout => \Add_add_temp_4\,
            ltout => OPEN,
            carryin => \bfn_22_19_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15973\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_3_lut_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59587\,
            in2 => \N__59578\,
            in3 => \N__59563\,
            lcout => \Add_add_temp_5\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15973\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15974\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_4_lut_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59560\,
            in2 => \N__59551\,
            in3 => \N__59539\,
            lcout => \Add_add_temp_6\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15974\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15975\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_5_lut_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59536\,
            in2 => \N__59527\,
            in3 => \N__59512\,
            lcout => \Add_add_temp_7\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15975\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15976\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_6_lut_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61561\,
            in2 => \N__59509\,
            in3 => \N__59494\,
            lcout => \Add_add_temp_8\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15976\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15977\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_7_lut_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62035\,
            in2 => \N__59749\,
            in3 => \N__59737\,
            lcout => \Add_add_temp_9\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15977\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15978\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_8_lut_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59734\,
            in2 => \N__59725\,
            in3 => \N__59710\,
            lcout => \Add_add_temp_10\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15978\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15979\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_9_lut_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59707\,
            in2 => \N__67510\,
            in3 => \N__59701\,
            lcout => \Add_add_temp_11\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15979\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15980\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_10_lut_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67492\,
            in2 => \N__59698\,
            in3 => \N__59686\,
            lcout => \Add_add_temp_12\,
            ltout => OPEN,
            carryin => \bfn_22_20_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15981\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_11_lut_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67210\,
            in2 => \N__59683\,
            in3 => \N__59671\,
            lcout => \Add_add_temp_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15981\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15982\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_12_lut_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67168\,
            in2 => \N__59668\,
            in3 => \N__59656\,
            lcout => \Add_add_temp_14\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15982\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15983\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_13_lut_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59653\,
            in2 => \N__67126\,
            in3 => \N__59644\,
            lcout => \Add_add_temp_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15983\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15984\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_14_lut_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67081\,
            in2 => \N__59641\,
            in3 => \N__59623\,
            lcout => \Add_add_temp_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15984\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15985\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_15_lut_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67042\,
            in2 => \N__59923\,
            in3 => \N__59908\,
            lcout => \Add_add_temp_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15985\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15986\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_16_lut_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67843\,
            in2 => \N__59905\,
            in3 => \N__59890\,
            lcout => \Add_add_temp_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15986\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15987\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_17_lut_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59887\,
            in2 => \N__67816\,
            in3 => \N__59875\,
            lcout => \Add_add_temp_19\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15987\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15988\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_18_lut_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67765\,
            in2 => \N__59872\,
            in3 => \N__59857\,
            lcout => \Add_add_temp_20\,
            ltout => OPEN,
            carryin => \bfn_22_21_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15989\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_19_lut_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67702\,
            in2 => \N__59854\,
            in3 => \N__59839\,
            lcout => \Add_add_temp_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15989\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15990\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_20_lut_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67651\,
            in2 => \N__59836\,
            in3 => \N__59821\,
            lcout => \Add_add_temp_22\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15990\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15991\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_21_lut_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59818\,
            in2 => \N__67588\,
            in3 => \N__59806\,
            lcout => \Add_add_temp_23\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15991\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15992\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_22_lut_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59803\,
            in2 => \N__68500\,
            in3 => \N__59770\,
            lcout => \Add_add_temp_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15992\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15993\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_23_lut_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68218\,
            in2 => \N__59767\,
            in3 => \N__59752\,
            lcout => \Add_add_temp_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15993\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15994\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_24_lut_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60055\,
            in2 => \N__68143\,
            in3 => \N__60043\,
            lcout => \Add_add_temp_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15994\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15995\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_25_lut_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68080\,
            in2 => \N__60040\,
            in3 => \N__60025\,
            lcout => \Add_add_temp_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15995\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15996\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_26_lut_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68017\,
            in2 => \N__60022\,
            in3 => \N__59992\,
            lcout => \Add_add_temp_28\,
            ltout => OPEN,
            carryin => \bfn_22_22_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15997\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_27_lut_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67933\,
            in2 => \N__59989\,
            in3 => \N__59956\,
            lcout => \Add_add_temp_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15997\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15998\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_28_lut_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68965\,
            in2 => \N__59953\,
            in3 => \N__59935\,
            lcout => \Add_add_temp_30\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15998\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15999\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_29_lut_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68910\,
            in2 => \N__60447\,
            in3 => \N__59932\,
            lcout => \Add_add_temp_31\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15999\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n16000\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_30_lut_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60441\,
            in2 => \N__68839\,
            in3 => \N__59929\,
            lcout => \Add_add_temp_32\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n16000\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n16001\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_31_lut_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60443\,
            in2 => \N__68770\,
            in3 => \N__59926\,
            lcout => \Add_add_temp_33\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n16001\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n16002\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_32_lut_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68698\,
            in2 => \N__60448\,
            in3 => \N__60451\,
            lcout => \Add_add_temp_34\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n16002\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n16003\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_33_lut_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60442\,
            in1 => \N__69045\,
            in2 => \_gnd_net_\,
            in3 => \N__60415\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i13263_4_lut_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__60556\,
            in1 => \N__60398\,
            in2 => \N__60375\,
            in3 => \N__60341\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n15200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_278_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__60321\,
            in1 => \N__60303\,
            in2 => \N__60292\,
            in3 => \N__60270\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20680_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_279_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__60251\,
            in1 => \N__60215\,
            in2 => \N__60199\,
            in3 => \N__60174\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_284_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__60111\,
            in1 => \N__60093\,
            in2 => \N__60147\,
            in3 => \N__60069\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_2_lut_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60140\,
            in2 => \_gnd_net_\,
            in3 => \N__60123\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_276_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__60110\,
            in1 => \N__60092\,
            in2 => \N__60079\,
            in3 => \N__60068\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n19761_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_277_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__62660\,
            in1 => \N__62687\,
            in2 => \N__60559\,
            in3 => \N__62714\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_22_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64914\,
            in2 => \N__64753\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n69\,
            ltout => OPEN,
            carryin => \bfn_22_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18234\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_22_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60550\,
            in2 => \N__64450\,
            in3 => \N__60535\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n115\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18234\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18235\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_22_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62629\,
            in2 => \N__64220\,
            in3 => \N__60523\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n164\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18235\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18236\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_22_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62620\,
            in2 => \N__63967\,
            in3 => \N__60511\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n213\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18236\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18237\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_22_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62611\,
            in2 => \N__63668\,
            in3 => \N__60499\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n262\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18237\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18238\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_22_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62602\,
            in2 => \N__63383\,
            in3 => \N__60484\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n311\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18238\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18239\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_22_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62593\,
            in2 => \N__63109\,
            in3 => \N__60469\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n360\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18239\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18240\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_22_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62584\,
            in2 => \N__66829\,
            in3 => \N__60454\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n409\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18240\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18241\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_22_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62575\,
            in2 => \N__66631\,
            in3 => \N__60664\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n458\,
            ltout => OPEN,
            carryin => \bfn_22_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18242\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_22_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62830\,
            in2 => \N__66349\,
            in3 => \N__60652\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n507\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18242\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18243\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_22_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62821\,
            in2 => \N__66086\,
            in3 => \N__60640\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n556\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18243\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18244\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_22_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62812\,
            in2 => \N__65828\,
            in3 => \N__60628\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n605\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18244\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18245\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_22_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62803\,
            in2 => \N__65596\,
            in3 => \N__60613\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n654\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18245\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18246\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_22_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65384\,
            in2 => \N__62794\,
            in3 => \N__60598\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n703\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18246\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18247\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_22_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65194\,
            in2 => \N__62782\,
            in3 => \N__60580\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n758\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18247\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_LUT4_0_LC_22_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60577\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_22_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64960\,
            in2 => \N__64758\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n78\,
            ltout => OPEN,
            carryin => \bfn_22_28_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18279\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_22_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60748\,
            in2 => \N__64496\,
            in3 => \N__60742\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n124\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18279\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18280\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_22_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60739\,
            in2 => \N__64243\,
            in3 => \N__60733\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n173\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18280\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18281\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_22_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60730\,
            in2 => \N__63979\,
            in3 => \N__60724\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n222\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18281\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18282\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_22_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60721\,
            in2 => \N__63669\,
            in3 => \N__60715\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n271\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18282\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18283\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_22_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60712\,
            in2 => \N__63405\,
            in3 => \N__60706\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n320\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18283\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18284\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_22_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60703\,
            in2 => \N__63131\,
            in3 => \N__60697\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n369\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18284\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18285\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_22_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66922\,
            in2 => \N__60694\,
            in3 => \N__60685\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n418\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18285\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18286\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_22_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60682\,
            in2 => \N__66640\,
            in3 => \N__60676\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n467\,
            ltout => OPEN,
            carryin => \bfn_22_29_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18287\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_22_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61063\,
            in2 => \N__66361\,
            in3 => \N__61057\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n516\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18287\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18288\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_22_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61054\,
            in2 => \N__66098\,
            in3 => \N__61048\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n565\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18288\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18289\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_22_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61045\,
            in2 => \N__65844\,
            in3 => \N__61039\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n614\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18289\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18290\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_22_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61036\,
            in2 => \N__65611\,
            in3 => \N__61030\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n663\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18290\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18291\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_22_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65388\,
            in2 => \N__61027\,
            in3 => \N__61018\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n712\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18291\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18292\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_22_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65201\,
            in2 => \N__61015\,
            in3 => \N__60991\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n770\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18292\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_LUT4_0_LC_22_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60988\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60939\,
            in2 => \N__67456\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_1\,
            ltout => OPEN,
            carryin => \bfn_23_11_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17521\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67413\,
            in2 => \N__61150\,
            in3 => \N__61141\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_2\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17521\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17522\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61138\,
            in2 => \N__67457\,
            in3 => \N__61132\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_3\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17522\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17523\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67417\,
            in2 => \N__61129\,
            in3 => \N__61120\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_4\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17523\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17524\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61117\,
            in2 => \N__67458\,
            in3 => \N__61111\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_5\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17524\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17525\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67421\,
            in2 => \N__61108\,
            in3 => \N__61099\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_6\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17525\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17526\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61096\,
            in2 => \N__67459\,
            in3 => \N__61090\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_7\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17526\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17527\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67425\,
            in2 => \N__61087\,
            in3 => \N__61078\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_8\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17527\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17528\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67426\,
            in2 => \N__61075\,
            in3 => \N__61066\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_9\,
            ltout => OPEN,
            carryin => \bfn_23_12_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17529\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61288\,
            in2 => \N__67460\,
            in3 => \N__61282\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_10\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17529\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17530\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61279\,
            in2 => \N__67463\,
            in3 => \N__61273\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_11\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17530\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17531\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_23_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61270\,
            in2 => \N__67461\,
            in3 => \N__61264\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_12\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17531\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17532\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61261\,
            in2 => \N__67464\,
            in3 => \N__61255\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17532\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17533\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61252\,
            in2 => \N__67462\,
            in3 => \N__61246\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_14\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17533\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n17534\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61243\,
            in2 => \N__61213\,
            in3 => \N__61183\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n738\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n17534\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_LUT4_0_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61180\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_20_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__69253\,
            in1 => \N__69204\,
            in2 => \N__69298\,
            in3 => \N__66976\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19932\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011001010"
        )
    port map (
            in0 => \N__61388\,
            in1 => \N__69294\,
            in2 => \N__61476\,
            in3 => \N__69252\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13172_2_lut_3_lut_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__68728\,
            in1 => \_gnd_net_\,
            in2 => \N__61480\,
            in3 => \N__61387\,
            lcout => OPEN,
            ltout => \foc.dVoltage_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_122_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__68106\,
            in1 => \N__68727\,
            in2 => \N__61507\,
            in3 => \N__61486\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_125_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__61492\,
            in1 => \N__68049\,
            in2 => \N__61504\,
            in3 => \N__61318\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.equal_13243_i14_2_lut_3_lut_3_lut_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__61382\,
            in1 => \N__68464\,
            in2 => \_gnd_net_\,
            in3 => \N__61469\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13165_2_lut_3_lut_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__68107\,
            in1 => \_gnd_net_\,
            in2 => \N__61390\,
            in3 => \N__61470\,
            lcout => \foc.dVoltage_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13166_2_lut_3_lut_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__61471\,
            in1 => \N__68050\,
            in2 => \_gnd_net_\,
            in3 => \N__61386\,
            lcout => \foc.dVoltage_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_53_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__66949\,
            in1 => \N__68550\,
            in2 => \N__69155\,
            in3 => \N__68601\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__67678\,
            in1 => \N__67732\,
            in2 => \_gnd_net_\,
            in3 => \N__67783\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_3_lut_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__69203\,
            in1 => \N__69251\,
            in2 => \_gnd_net_\,
            in3 => \N__69293\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1202_3_lut_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__67673\,
            in1 => \N__67728\,
            in2 => \_gnd_net_\,
            in3 => \N__67779\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_11_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__67610\,
            in1 => \N__68459\,
            in2 => \N__61510\,
            in3 => \N__67548\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i10_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__62395\,
            in1 => \N__62017\,
            in2 => \_gnd_net_\,
            in3 => \N__61888\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i11_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__62018\,
            in1 => \N__61891\,
            in2 => \_gnd_net_\,
            in3 => \N__61738\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i8_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__62347\,
            in1 => \N__61890\,
            in2 => \_gnd_net_\,
            in3 => \N__62021\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i13_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__61783\,
            in1 => \N__62019\,
            in2 => \_gnd_net_\,
            in3 => \N__61889\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i7_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__62020\,
            in1 => \N__61892\,
            in2 => \_gnd_net_\,
            in3 => \N__62443\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i26_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001110"
        )
    port map (
            in0 => \N__61656\,
            in1 => \N__61886\,
            in2 => \N__62015\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i28_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__61686\,
            in1 => \N__61885\,
            in2 => \_gnd_net_\,
            in3 => \N__61981\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i9_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001110"
        )
    port map (
            in0 => \N__62371\,
            in1 => \N__61887\,
            in2 => \N__62016\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i17_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__62230\,
            in1 => \N__61884\,
            in2 => \_gnd_net_\,
            in3 => \N__61977\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i747_4_lut_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__61717\,
            in1 => \N__61687\,
            in2 => \N__61660\,
            in3 => \N__61636\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_147_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__62143\,
            in1 => \N__61630\,
            in2 => \N__61600\,
            in3 => \N__61596\,
            lcout => \Saturate_out1_31__N_266\,
            ltout => \Saturate_out1_31__N_266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i12_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001110"
        )
    port map (
            in0 => \N__61975\,
            in1 => \N__61762\,
            in2 => \N__61564\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i15_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__62254\,
            in1 => \N__61883\,
            in2 => \_gnd_net_\,
            in3 => \N__61976\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i16_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__61894\,
            in1 => \N__62023\,
            in2 => \_gnd_net_\,
            in3 => \N__62311\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i4_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__62028\,
            in1 => \N__61899\,
            in2 => \_gnd_net_\,
            in3 => \N__62535\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i22_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__61897\,
            in1 => \N__62026\,
            in2 => \_gnd_net_\,
            in3 => \N__61555\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i23_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__62027\,
            in1 => \N__61898\,
            in2 => \_gnd_net_\,
            in3 => \N__61531\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i21_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__61896\,
            in1 => \N__62025\,
            in2 => \_gnd_net_\,
            in3 => \N__62065\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i14_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__62022\,
            in1 => \N__61893\,
            in2 => \_gnd_net_\,
            in3 => \N__62283\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i5_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__61900\,
            in1 => \N__62029\,
            in2 => \_gnd_net_\,
            in3 => \N__62460\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i19_LC_23_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__62024\,
            in1 => \N__61895\,
            in2 => \_gnd_net_\,
            in3 => \N__62203\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_140_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__62483\,
            in1 => \N__62565\,
            in2 => \N__62517\,
            in3 => \N__62534\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_141_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__62459\,
            in1 => \N__62435\,
            in2 => \N__61798\,
            in3 => \N__62411\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i729_4_lut_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__62367\,
            in1 => \N__62388\,
            in2 => \N__61795\,
            in3 => \N__62340\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n22_adj_519_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_142_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__61754\,
            in1 => \N__61776\,
            in2 => \N__61792\,
            in3 => \N__61731\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_133_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__62323\,
            in1 => \N__61775\,
            in2 => \N__61758\,
            in3 => \N__61730\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_130_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62564\,
            in2 => \_gnd_net_\,
            in3 => \N__62547\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_131_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__62536\,
            in1 => \N__62516\,
            in2 => \N__62494\,
            in3 => \N__62467\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19777_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_132_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__62461\,
            in1 => \N__62436\,
            in2 => \N__62419\,
            in3 => \N__62415\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i13268_4_lut_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__62387\,
            in1 => \N__62366\,
            in2 => \N__62350\,
            in3 => \N__62339\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_134_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__62317\,
            in1 => \N__62300\,
            in2 => \N__62279\,
            in3 => \N__62243\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.n19746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_136_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__62214\,
            in1 => \N__62190\,
            in2 => \N__62179\,
            in3 => \N__62165\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i31_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62130\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_285_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__62731\,
            in1 => \N__62721\,
            in2 => \N__62698\,
            in3 => \N__62667\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n20718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_23_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64910\,
            in2 => \N__64754\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n72\,
            ltout => OPEN,
            carryin => \bfn_23_25_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18249\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_23_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62635\,
            in2 => \N__64451\,
            in3 => \N__62623\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n118\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18249\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18250\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_23_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64261\,
            in2 => \N__64241\,
            in3 => \N__62614\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n167\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18250\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18251\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_23_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64000\,
            in2 => \N__63980\,
            in3 => \N__62605\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n216\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18251\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_23_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63706\,
            in2 => \N__63686\,
            in3 => \N__62596\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n265\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18252\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18253\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_23_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63424\,
            in2 => \N__63384\,
            in3 => \N__62587\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n314\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18253\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18254\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_23_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63148\,
            in2 => \N__63136\,
            in3 => \N__62578\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n363\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18254\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18255\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_23_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62845\,
            in2 => \N__66830\,
            in3 => \N__62833\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n412\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18255\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18256\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_23_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66649\,
            in2 => \N__66639\,
            in3 => \N__62824\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n461\,
            ltout => OPEN,
            carryin => \bfn_23_26_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18257\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_23_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66379\,
            in2 => \N__66359\,
            in3 => \N__62815\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n510\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18257\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18258\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_23_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66118\,
            in2 => \N__66099\,
            in3 => \N__62806\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n559\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18258\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18259\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_23_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65863\,
            in2 => \N__65829\,
            in3 => \N__62797\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n608\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18259\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18260\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_23_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65629\,
            in2 => \N__65609\,
            in3 => \N__62785\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n657\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18260\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18261\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_23_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65385\,
            in2 => \N__65404\,
            in3 => \N__62773\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n706\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18261\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18262\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_23_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65202\,
            in2 => \N__65218\,
            in3 => \N__62755\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n762\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18262\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_LUT4_0_LC_23_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62752\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_23_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64956\,
            in2 => \N__64759\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n75\,
            ltout => OPEN,
            carryin => \bfn_23_27_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18264\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_23_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64507\,
            in2 => \N__64501\,
            in3 => \N__64252\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n121\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18264\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18265\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_23_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64249\,
            in2 => \N__64242\,
            in3 => \N__63991\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n170\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18265\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18266\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_23_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63988\,
            in2 => \N__63974\,
            in3 => \N__63697\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n219\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18266\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18267\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_23_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63694\,
            in2 => \N__63687\,
            in3 => \N__63415\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n268\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18267\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18268\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_23_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63412\,
            in2 => \N__63406\,
            in3 => \N__63139\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n317\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18268\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18269\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_23_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63110\,
            in2 => \N__62854\,
            in3 => \N__62836\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n366\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18269\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18270\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_23_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66937\,
            in2 => \N__66920\,
            in3 => \N__66643\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n415\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18270\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18271\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_23_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66598\,
            in2 => \N__66388\,
            in3 => \N__66370\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n464\,
            ltout => OPEN,
            carryin => \bfn_23_28_0_\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18272\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_23_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66367\,
            in2 => \N__66360\,
            in3 => \N__66109\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n513\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18272\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18273\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_23_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66106\,
            in2 => \N__66100\,
            in3 => \N__65854\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n562\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18273\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18274\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_23_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65851\,
            in2 => \N__65843\,
            in3 => \N__65620\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n611\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18274\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18275\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_23_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65617\,
            in2 => \N__65610\,
            in3 => \N__65392\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n660\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18275\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18276\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_23_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65389\,
            in2 => \N__65227\,
            in3 => \N__65206\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n709\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18276\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18277\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_23_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65193\,
            in2 => \N__65038\,
            in3 => \N__67000\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n766\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_Q_Current_Control.n18277\,
            carryout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_LUT4_0_LC_23_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66997\,
            lcout => \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_19_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__66964\,
            in1 => \N__68594\,
            in2 => \N__68549\,
            in3 => \N__68649\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_15_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__67516\,
            in1 => \N__67964\,
            in2 => \N__67900\,
            in3 => \N__68942\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_17_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__68862\,
            in1 => \N__68721\,
            in2 => \N__66967\,
            in3 => \N__68793\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13232_4_lut_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__66943\,
            in1 => \N__68460\,
            in2 => \N__68179\,
            in3 => \N__67547\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13251_4_lut_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__68099\,
            in1 => \N__67970\,
            in2 => \N__66958\,
            in3 => \N__68047\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__68861\,
            in1 => \N__67885\,
            in2 => \N__66955\,
            in3 => \N__68936\,
            lcout => OPEN,
            ltout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_27_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__68720\,
            in1 => \N__68792\,
            in2 => \N__66952\,
            in3 => \N__68648\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12921_2_lut_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67611\,
            in2 => \_gnd_net_\,
            in3 => \N__67677\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n14851\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_14_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__68100\,
            in1 => \N__68048\,
            in2 => \N__68180\,
            in3 => \N__67522\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_2_lut_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67503\,
            in1 => \N__67485\,
            in2 => \N__67474\,
            in3 => \_gnd_net_\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20184\,
            ltout => OPEN,
            carryin => \bfn_24_16_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15568\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_3_lut_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67216\,
            in1 => \N__67203\,
            in2 => \N__67192\,
            in3 => \N__67177\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20186\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15568\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15569\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_4_lut_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67174\,
            in1 => \N__67161\,
            in2 => \N__67150\,
            in3 => \N__67135\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20188\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15569\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15570\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_5_lut_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67132\,
            in1 => \N__67116\,
            in2 => \N__67105\,
            in3 => \N__67090\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20190\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15570\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15571\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_6_lut_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67087\,
            in1 => \N__67077\,
            in2 => \N__67066\,
            in3 => \N__67051\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20192\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15571\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15572\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_lut_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67048\,
            in1 => \N__67032\,
            in2 => \N__67021\,
            in3 => \N__67003\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20194\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15572\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15573\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_0_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68418\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15573\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_1_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__68434\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_0_THRU_CO\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_8_lut_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67861\,
            in1 => \N__67855\,
            in2 => \N__67842\,
            in3 => \N__67825\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20196\,
            ltout => OPEN,
            carryin => \bfn_24_17_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15574\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_9_lut_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__67822\,
            in1 => \N__67809\,
            in2 => \N__67798\,
            in3 => \N__67768\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.n20198\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15574\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15575\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_10_lut_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67758\,
            in2 => \N__67747\,
            in3 => \N__67717\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15575\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15576\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_11_lut_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67714\,
            in2 => \N__67695\,
            in3 => \N__67654\,
            lcout => \foc.preSatVoltage_10_adj_2311\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15576\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15577\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_12_lut_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67650\,
            in2 => \N__67633\,
            in3 => \N__67591\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15577\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15578\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_13_lut_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67581\,
            in2 => \N__67570\,
            in3 => \N__67525\,
            lcout => \foc.preSatVoltage_12_adj_2330\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15578\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15579\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_lut_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68496\,
            in2 => \N__68479\,
            in3 => \N__68440\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15579\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15580\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_THRU_CRY_0_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68422\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15580\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15580_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_15_lut_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68214\,
            in2 => \N__68203\,
            in3 => \N__68146\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14\,
            ltout => OPEN,
            carryin => \bfn_24_18_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15581\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_16_lut_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68136\,
            in2 => \N__68125\,
            in3 => \N__68083\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_15\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15581\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15582\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_17_lut_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68076\,
            in2 => \N__68065\,
            in3 => \N__68020\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15582\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_18_lut_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68013\,
            in2 => \N__67996\,
            in3 => \N__67936\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15583\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_19_lut_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67929\,
            in2 => \N__67915\,
            in3 => \N__67864\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_18\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15584\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_20_lut_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68977\,
            in2 => \N__68961\,
            in3 => \N__68914\,
            lcout => \foc.preSatVoltage_19_adj_2329\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15585\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_21_lut_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68911\,
            in2 => \N__68890\,
            in3 => \N__68842\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_20\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15586\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15587\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_22_lut_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68829\,
            in2 => \N__68818\,
            in3 => \N__68773\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_21\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15587\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15588\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_23_lut_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68769\,
            in2 => \N__68746\,
            in3 => \N__68701\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_22\,
            ltout => OPEN,
            carryin => \bfn_24_19_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_24_lut_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68697\,
            in2 => \N__68674\,
            in3 => \N__68626\,
            lcout => \foc.preSatVoltage_23_adj_2328\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15589\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_25_lut_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69059\,
            in2 => \N__68623\,
            in3 => \N__68572\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15590\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_26_lut_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68569\,
            in2 => \N__69071\,
            in3 => \N__68518\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15591\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_27_lut_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69063\,
            in2 => \N__68515\,
            in3 => \N__69268\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15592\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_28_lut_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69265\,
            in2 => \N__69072\,
            in3 => \N__69226\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15593\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_29_lut_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69067\,
            in2 => \N__69223\,
            in3 => \N__69175\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15594\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15595\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_30_lut_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69172\,
            in2 => \N__69073\,
            in3 => \N__69130\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_29\,
            ltout => OPEN,
            carryin => \foc.u_DQ_Current_Control.u_D_Current_Control.n15595\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15596\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_31_lut_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69043\,
            in2 => \N__69127\,
            in3 => \N__69076\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30\,
            ltout => OPEN,
            carryin => \bfn_24_20_0_\,
            carryout => \foc.u_DQ_Current_Control.u_D_Current_Control.n15597\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_32_lut_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__69044\,
            in1 => \N__69025\,
            in2 => \_gnd_net_\,
            in3 => \N__69013\,
            lcout => \foc.u_DQ_Current_Control.u_D_Current_Control.Voltage_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
