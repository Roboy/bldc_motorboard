// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 16 2019 20:28:04

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    inout PIN_6;
    inout PIN_5;
    inout PIN_4;
    output PIN_3;
    output PIN_24;
    output PIN_23;
    output PIN_22;
    input PIN_21;
    input PIN_20;
    output PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    inout PIN_11;
    inout PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__81286;
    wire N__81285;
    wire N__81284;
    wire N__81277;
    wire N__81276;
    wire N__81275;
    wire N__81268;
    wire N__81267;
    wire N__81266;
    wire N__81259;
    wire N__81258;
    wire N__81257;
    wire N__81250;
    wire N__81249;
    wire N__81248;
    wire N__81241;
    wire N__81240;
    wire N__81239;
    wire N__81232;
    wire N__81231;
    wire N__81230;
    wire N__81223;
    wire N__81222;
    wire N__81221;
    wire N__81214;
    wire N__81213;
    wire N__81212;
    wire N__81205;
    wire N__81204;
    wire N__81203;
    wire N__81196;
    wire N__81195;
    wire N__81194;
    wire N__81187;
    wire N__81186;
    wire N__81185;
    wire N__81178;
    wire N__81177;
    wire N__81176;
    wire N__81169;
    wire N__81168;
    wire N__81167;
    wire N__81160;
    wire N__81159;
    wire N__81158;
    wire N__81151;
    wire N__81150;
    wire N__81149;
    wire N__81142;
    wire N__81141;
    wire N__81140;
    wire N__81133;
    wire N__81132;
    wire N__81131;
    wire N__81114;
    wire N__81111;
    wire N__81108;
    wire N__81105;
    wire N__81104;
    wire N__81103;
    wire N__81100;
    wire N__81097;
    wire N__81094;
    wire N__81091;
    wire N__81086;
    wire N__81081;
    wire N__81078;
    wire N__81075;
    wire N__81072;
    wire N__81071;
    wire N__81068;
    wire N__81065;
    wire N__81062;
    wire N__81059;
    wire N__81058;
    wire N__81057;
    wire N__81054;
    wire N__81051;
    wire N__81048;
    wire N__81045;
    wire N__81042;
    wire N__81039;
    wire N__81036;
    wire N__81033;
    wire N__81032;
    wire N__81031;
    wire N__81028;
    wire N__81025;
    wire N__81020;
    wire N__81015;
    wire N__81006;
    wire N__81003;
    wire N__81002;
    wire N__80999;
    wire N__80996;
    wire N__80991;
    wire N__80988;
    wire N__80987;
    wire N__80986;
    wire N__80983;
    wire N__80982;
    wire N__80979;
    wire N__80976;
    wire N__80975;
    wire N__80974;
    wire N__80973;
    wire N__80970;
    wire N__80967;
    wire N__80966;
    wire N__80963;
    wire N__80960;
    wire N__80957;
    wire N__80952;
    wire N__80951;
    wire N__80948;
    wire N__80945;
    wire N__80944;
    wire N__80943;
    wire N__80942;
    wire N__80941;
    wire N__80940;
    wire N__80937;
    wire N__80928;
    wire N__80925;
    wire N__80924;
    wire N__80923;
    wire N__80922;
    wire N__80921;
    wire N__80920;
    wire N__80919;
    wire N__80918;
    wire N__80913;
    wire N__80908;
    wire N__80905;
    wire N__80900;
    wire N__80899;
    wire N__80894;
    wire N__80889;
    wire N__80888;
    wire N__80885;
    wire N__80882;
    wire N__80875;
    wire N__80872;
    wire N__80871;
    wire N__80868;
    wire N__80867;
    wire N__80864;
    wire N__80859;
    wire N__80856;
    wire N__80853;
    wire N__80850;
    wire N__80847;
    wire N__80844;
    wire N__80843;
    wire N__80840;
    wire N__80837;
    wire N__80834;
    wire N__80831;
    wire N__80828;
    wire N__80825;
    wire N__80820;
    wire N__80813;
    wire N__80810;
    wire N__80807;
    wire N__80804;
    wire N__80799;
    wire N__80796;
    wire N__80793;
    wire N__80790;
    wire N__80787;
    wire N__80784;
    wire N__80781;
    wire N__80776;
    wire N__80769;
    wire N__80764;
    wire N__80757;
    wire N__80748;
    wire N__80747;
    wire N__80746;
    wire N__80743;
    wire N__80742;
    wire N__80741;
    wire N__80740;
    wire N__80739;
    wire N__80738;
    wire N__80737;
    wire N__80736;
    wire N__80735;
    wire N__80734;
    wire N__80733;
    wire N__80730;
    wire N__80729;
    wire N__80726;
    wire N__80723;
    wire N__80720;
    wire N__80719;
    wire N__80718;
    wire N__80715;
    wire N__80712;
    wire N__80711;
    wire N__80708;
    wire N__80707;
    wire N__80704;
    wire N__80703;
    wire N__80700;
    wire N__80697;
    wire N__80696;
    wire N__80693;
    wire N__80688;
    wire N__80685;
    wire N__80682;
    wire N__80679;
    wire N__80674;
    wire N__80673;
    wire N__80672;
    wire N__80671;
    wire N__80668;
    wire N__80665;
    wire N__80662;
    wire N__80659;
    wire N__80656;
    wire N__80655;
    wire N__80650;
    wire N__80647;
    wire N__80644;
    wire N__80641;
    wire N__80638;
    wire N__80635;
    wire N__80632;
    wire N__80627;
    wire N__80624;
    wire N__80619;
    wire N__80618;
    wire N__80617;
    wire N__80616;
    wire N__80615;
    wire N__80612;
    wire N__80609;
    wire N__80606;
    wire N__80605;
    wire N__80602;
    wire N__80595;
    wire N__80592;
    wire N__80589;
    wire N__80586;
    wire N__80581;
    wire N__80576;
    wire N__80575;
    wire N__80568;
    wire N__80565;
    wire N__80562;
    wire N__80557;
    wire N__80554;
    wire N__80549;
    wire N__80546;
    wire N__80543;
    wire N__80540;
    wire N__80535;
    wire N__80532;
    wire N__80527;
    wire N__80524;
    wire N__80521;
    wire N__80518;
    wire N__80515;
    wire N__80510;
    wire N__80509;
    wire N__80508;
    wire N__80505;
    wire N__80502;
    wire N__80497;
    wire N__80492;
    wire N__80487;
    wire N__80484;
    wire N__80481;
    wire N__80478;
    wire N__80471;
    wire N__80466;
    wire N__80463;
    wire N__80458;
    wire N__80453;
    wire N__80444;
    wire N__80433;
    wire N__80432;
    wire N__80431;
    wire N__80430;
    wire N__80429;
    wire N__80428;
    wire N__80427;
    wire N__80426;
    wire N__80425;
    wire N__80424;
    wire N__80423;
    wire N__80422;
    wire N__80421;
    wire N__80420;
    wire N__80419;
    wire N__80418;
    wire N__80417;
    wire N__80416;
    wire N__80415;
    wire N__80414;
    wire N__80413;
    wire N__80412;
    wire N__80407;
    wire N__80404;
    wire N__80403;
    wire N__80402;
    wire N__80401;
    wire N__80400;
    wire N__80399;
    wire N__80398;
    wire N__80397;
    wire N__80396;
    wire N__80395;
    wire N__80392;
    wire N__80389;
    wire N__80386;
    wire N__80385;
    wire N__80382;
    wire N__80379;
    wire N__80376;
    wire N__80373;
    wire N__80368;
    wire N__80365;
    wire N__80360;
    wire N__80355;
    wire N__80344;
    wire N__80341;
    wire N__80338;
    wire N__80329;
    wire N__80328;
    wire N__80325;
    wire N__80324;
    wire N__80323;
    wire N__80322;
    wire N__80321;
    wire N__80320;
    wire N__80319;
    wire N__80318;
    wire N__80315;
    wire N__80312;
    wire N__80307;
    wire N__80304;
    wire N__80299;
    wire N__80296;
    wire N__80293;
    wire N__80288;
    wire N__80283;
    wire N__80276;
    wire N__80267;
    wire N__80266;
    wire N__80265;
    wire N__80264;
    wire N__80263;
    wire N__80262;
    wire N__80261;
    wire N__80260;
    wire N__80259;
    wire N__80256;
    wire N__80253;
    wire N__80250;
    wire N__80241;
    wire N__80236;
    wire N__80233;
    wire N__80230;
    wire N__80227;
    wire N__80224;
    wire N__80221;
    wire N__80218;
    wire N__80213;
    wire N__80206;
    wire N__80203;
    wire N__80200;
    wire N__80197;
    wire N__80186;
    wire N__80183;
    wire N__80180;
    wire N__80171;
    wire N__80162;
    wire N__80155;
    wire N__80136;
    wire N__80135;
    wire N__80132;
    wire N__80131;
    wire N__80128;
    wire N__80125;
    wire N__80122;
    wire N__80119;
    wire N__80116;
    wire N__80113;
    wire N__80110;
    wire N__80107;
    wire N__80100;
    wire N__80099;
    wire N__80098;
    wire N__80097;
    wire N__80096;
    wire N__80095;
    wire N__80094;
    wire N__80093;
    wire N__80090;
    wire N__80087;
    wire N__80084;
    wire N__80081;
    wire N__80080;
    wire N__80079;
    wire N__80076;
    wire N__80073;
    wire N__80070;
    wire N__80067;
    wire N__80064;
    wire N__80061;
    wire N__80060;
    wire N__80055;
    wire N__80052;
    wire N__80051;
    wire N__80048;
    wire N__80045;
    wire N__80044;
    wire N__80041;
    wire N__80036;
    wire N__80033;
    wire N__80032;
    wire N__80031;
    wire N__80030;
    wire N__80029;
    wire N__80026;
    wire N__80023;
    wire N__80020;
    wire N__80017;
    wire N__80016;
    wire N__80013;
    wire N__80010;
    wire N__80009;
    wire N__80008;
    wire N__80007;
    wire N__80004;
    wire N__80001;
    wire N__79998;
    wire N__79995;
    wire N__79992;
    wire N__79989;
    wire N__79988;
    wire N__79987;
    wire N__79986;
    wire N__79985;
    wire N__79984;
    wire N__79983;
    wire N__79980;
    wire N__79975;
    wire N__79972;
    wire N__79967;
    wire N__79964;
    wire N__79961;
    wire N__79958;
    wire N__79955;
    wire N__79954;
    wire N__79953;
    wire N__79952;
    wire N__79949;
    wire N__79948;
    wire N__79947;
    wire N__79944;
    wire N__79941;
    wire N__79938;
    wire N__79929;
    wire N__79922;
    wire N__79919;
    wire N__79914;
    wire N__79911;
    wire N__79908;
    wire N__79901;
    wire N__79892;
    wire N__79889;
    wire N__79886;
    wire N__79883;
    wire N__79878;
    wire N__79875;
    wire N__79868;
    wire N__79865;
    wire N__79860;
    wire N__79857;
    wire N__79848;
    wire N__79845;
    wire N__79842;
    wire N__79833;
    wire N__79830;
    wire N__79827;
    wire N__79824;
    wire N__79821;
    wire N__79814;
    wire N__79811;
    wire N__79800;
    wire N__79797;
    wire N__79796;
    wire N__79793;
    wire N__79792;
    wire N__79791;
    wire N__79788;
    wire N__79787;
    wire N__79786;
    wire N__79785;
    wire N__79784;
    wire N__79781;
    wire N__79778;
    wire N__79777;
    wire N__79776;
    wire N__79769;
    wire N__79766;
    wire N__79763;
    wire N__79760;
    wire N__79759;
    wire N__79758;
    wire N__79757;
    wire N__79756;
    wire N__79751;
    wire N__79746;
    wire N__79743;
    wire N__79740;
    wire N__79737;
    wire N__79734;
    wire N__79729;
    wire N__79728;
    wire N__79727;
    wire N__79724;
    wire N__79721;
    wire N__79718;
    wire N__79709;
    wire N__79704;
    wire N__79703;
    wire N__79702;
    wire N__79699;
    wire N__79698;
    wire N__79695;
    wire N__79692;
    wire N__79689;
    wire N__79686;
    wire N__79681;
    wire N__79678;
    wire N__79677;
    wire N__79674;
    wire N__79671;
    wire N__79668;
    wire N__79665;
    wire N__79662;
    wire N__79653;
    wire N__79650;
    wire N__79649;
    wire N__79648;
    wire N__79647;
    wire N__79646;
    wire N__79641;
    wire N__79632;
    wire N__79629;
    wire N__79628;
    wire N__79627;
    wire N__79626;
    wire N__79623;
    wire N__79622;
    wire N__79619;
    wire N__79616;
    wire N__79613;
    wire N__79608;
    wire N__79605;
    wire N__79602;
    wire N__79599;
    wire N__79596;
    wire N__79593;
    wire N__79590;
    wire N__79589;
    wire N__79588;
    wire N__79587;
    wire N__79582;
    wire N__79579;
    wire N__79576;
    wire N__79571;
    wire N__79568;
    wire N__79565;
    wire N__79560;
    wire N__79557;
    wire N__79554;
    wire N__79551;
    wire N__79548;
    wire N__79543;
    wire N__79542;
    wire N__79537;
    wire N__79532;
    wire N__79527;
    wire N__79522;
    wire N__79519;
    wire N__79516;
    wire N__79513;
    wire N__79510;
    wire N__79505;
    wire N__79502;
    wire N__79491;
    wire N__79490;
    wire N__79489;
    wire N__79488;
    wire N__79485;
    wire N__79484;
    wire N__79483;
    wire N__79482;
    wire N__79481;
    wire N__79478;
    wire N__79477;
    wire N__79476;
    wire N__79473;
    wire N__79472;
    wire N__79471;
    wire N__79468;
    wire N__79465;
    wire N__79464;
    wire N__79463;
    wire N__79458;
    wire N__79457;
    wire N__79456;
    wire N__79453;
    wire N__79450;
    wire N__79447;
    wire N__79444;
    wire N__79443;
    wire N__79442;
    wire N__79441;
    wire N__79440;
    wire N__79439;
    wire N__79436;
    wire N__79433;
    wire N__79428;
    wire N__79425;
    wire N__79422;
    wire N__79421;
    wire N__79420;
    wire N__79415;
    wire N__79412;
    wire N__79407;
    wire N__79404;
    wire N__79399;
    wire N__79398;
    wire N__79397;
    wire N__79396;
    wire N__79393;
    wire N__79388;
    wire N__79385;
    wire N__79380;
    wire N__79373;
    wire N__79370;
    wire N__79367;
    wire N__79366;
    wire N__79365;
    wire N__79364;
    wire N__79363;
    wire N__79362;
    wire N__79361;
    wire N__79360;
    wire N__79359;
    wire N__79358;
    wire N__79357;
    wire N__79356;
    wire N__79355;
    wire N__79354;
    wire N__79351;
    wire N__79348;
    wire N__79345;
    wire N__79342;
    wire N__79337;
    wire N__79334;
    wire N__79327;
    wire N__79324;
    wire N__79321;
    wire N__79316;
    wire N__79311;
    wire N__79308;
    wire N__79305;
    wire N__79300;
    wire N__79295;
    wire N__79288;
    wire N__79277;
    wire N__79274;
    wire N__79269;
    wire N__79266;
    wire N__79261;
    wire N__79248;
    wire N__79227;
    wire N__79226;
    wire N__79223;
    wire N__79220;
    wire N__79217;
    wire N__79214;
    wire N__79209;
    wire N__79206;
    wire N__79205;
    wire N__79204;
    wire N__79203;
    wire N__79200;
    wire N__79197;
    wire N__79194;
    wire N__79193;
    wire N__79192;
    wire N__79191;
    wire N__79190;
    wire N__79189;
    wire N__79186;
    wire N__79185;
    wire N__79184;
    wire N__79183;
    wire N__79182;
    wire N__79177;
    wire N__79174;
    wire N__79173;
    wire N__79172;
    wire N__79169;
    wire N__79168;
    wire N__79167;
    wire N__79164;
    wire N__79161;
    wire N__79158;
    wire N__79155;
    wire N__79152;
    wire N__79149;
    wire N__79148;
    wire N__79145;
    wire N__79142;
    wire N__79141;
    wire N__79140;
    wire N__79137;
    wire N__79132;
    wire N__79129;
    wire N__79126;
    wire N__79125;
    wire N__79120;
    wire N__79117;
    wire N__79114;
    wire N__79111;
    wire N__79110;
    wire N__79109;
    wire N__79108;
    wire N__79107;
    wire N__79106;
    wire N__79101;
    wire N__79096;
    wire N__79093;
    wire N__79088;
    wire N__79085;
    wire N__79084;
    wire N__79083;
    wire N__79078;
    wire N__79075;
    wire N__79072;
    wire N__79069;
    wire N__79066;
    wire N__79063;
    wire N__79060;
    wire N__79055;
    wire N__79052;
    wire N__79051;
    wire N__79046;
    wire N__79043;
    wire N__79040;
    wire N__79037;
    wire N__79034;
    wire N__79029;
    wire N__79022;
    wire N__79019;
    wire N__79016;
    wire N__79009;
    wire N__79006;
    wire N__79001;
    wire N__78998;
    wire N__78995;
    wire N__78994;
    wire N__78985;
    wire N__78980;
    wire N__78979;
    wire N__78978;
    wire N__78975;
    wire N__78970;
    wire N__78963;
    wire N__78960;
    wire N__78955;
    wire N__78952;
    wire N__78949;
    wire N__78946;
    wire N__78943;
    wire N__78938;
    wire N__78933;
    wire N__78926;
    wire N__78915;
    wire N__78912;
    wire N__78911;
    wire N__78908;
    wire N__78905;
    wire N__78904;
    wire N__78901;
    wire N__78898;
    wire N__78897;
    wire N__78896;
    wire N__78895;
    wire N__78892;
    wire N__78891;
    wire N__78890;
    wire N__78887;
    wire N__78884;
    wire N__78881;
    wire N__78876;
    wire N__78873;
    wire N__78870;
    wire N__78867;
    wire N__78852;
    wire N__78849;
    wire N__78846;
    wire N__78843;
    wire N__78842;
    wire N__78841;
    wire N__78838;
    wire N__78833;
    wire N__78830;
    wire N__78825;
    wire N__78824;
    wire N__78823;
    wire N__78822;
    wire N__78821;
    wire N__78820;
    wire N__78819;
    wire N__78818;
    wire N__78817;
    wire N__78816;
    wire N__78815;
    wire N__78814;
    wire N__78813;
    wire N__78812;
    wire N__78811;
    wire N__78810;
    wire N__78809;
    wire N__78808;
    wire N__78807;
    wire N__78806;
    wire N__78805;
    wire N__78804;
    wire N__78803;
    wire N__78802;
    wire N__78801;
    wire N__78800;
    wire N__78799;
    wire N__78798;
    wire N__78797;
    wire N__78796;
    wire N__78795;
    wire N__78794;
    wire N__78793;
    wire N__78792;
    wire N__78791;
    wire N__78790;
    wire N__78789;
    wire N__78788;
    wire N__78787;
    wire N__78786;
    wire N__78785;
    wire N__78784;
    wire N__78783;
    wire N__78782;
    wire N__78781;
    wire N__78780;
    wire N__78779;
    wire N__78778;
    wire N__78777;
    wire N__78776;
    wire N__78775;
    wire N__78774;
    wire N__78773;
    wire N__78772;
    wire N__78771;
    wire N__78770;
    wire N__78769;
    wire N__78768;
    wire N__78767;
    wire N__78766;
    wire N__78765;
    wire N__78764;
    wire N__78763;
    wire N__78762;
    wire N__78761;
    wire N__78760;
    wire N__78759;
    wire N__78758;
    wire N__78757;
    wire N__78756;
    wire N__78755;
    wire N__78754;
    wire N__78753;
    wire N__78752;
    wire N__78751;
    wire N__78750;
    wire N__78749;
    wire N__78748;
    wire N__78747;
    wire N__78746;
    wire N__78745;
    wire N__78744;
    wire N__78743;
    wire N__78742;
    wire N__78741;
    wire N__78740;
    wire N__78739;
    wire N__78738;
    wire N__78737;
    wire N__78736;
    wire N__78735;
    wire N__78734;
    wire N__78733;
    wire N__78732;
    wire N__78731;
    wire N__78730;
    wire N__78729;
    wire N__78728;
    wire N__78727;
    wire N__78726;
    wire N__78725;
    wire N__78724;
    wire N__78723;
    wire N__78722;
    wire N__78721;
    wire N__78720;
    wire N__78719;
    wire N__78718;
    wire N__78717;
    wire N__78716;
    wire N__78715;
    wire N__78714;
    wire N__78713;
    wire N__78712;
    wire N__78711;
    wire N__78710;
    wire N__78709;
    wire N__78708;
    wire N__78707;
    wire N__78706;
    wire N__78705;
    wire N__78704;
    wire N__78703;
    wire N__78702;
    wire N__78701;
    wire N__78700;
    wire N__78699;
    wire N__78698;
    wire N__78697;
    wire N__78696;
    wire N__78695;
    wire N__78694;
    wire N__78693;
    wire N__78692;
    wire N__78691;
    wire N__78690;
    wire N__78689;
    wire N__78688;
    wire N__78687;
    wire N__78686;
    wire N__78685;
    wire N__78684;
    wire N__78683;
    wire N__78682;
    wire N__78681;
    wire N__78680;
    wire N__78679;
    wire N__78678;
    wire N__78677;
    wire N__78676;
    wire N__78675;
    wire N__78674;
    wire N__78673;
    wire N__78672;
    wire N__78671;
    wire N__78670;
    wire N__78669;
    wire N__78668;
    wire N__78667;
    wire N__78666;
    wire N__78665;
    wire N__78664;
    wire N__78663;
    wire N__78662;
    wire N__78661;
    wire N__78660;
    wire N__78659;
    wire N__78658;
    wire N__78657;
    wire N__78656;
    wire N__78655;
    wire N__78654;
    wire N__78653;
    wire N__78652;
    wire N__78651;
    wire N__78650;
    wire N__78649;
    wire N__78648;
    wire N__78647;
    wire N__78646;
    wire N__78645;
    wire N__78644;
    wire N__78643;
    wire N__78642;
    wire N__78641;
    wire N__78640;
    wire N__78639;
    wire N__78638;
    wire N__78637;
    wire N__78636;
    wire N__78635;
    wire N__78634;
    wire N__78633;
    wire N__78632;
    wire N__78631;
    wire N__78630;
    wire N__78629;
    wire N__78628;
    wire N__78627;
    wire N__78626;
    wire N__78625;
    wire N__78624;
    wire N__78623;
    wire N__78622;
    wire N__78621;
    wire N__78620;
    wire N__78619;
    wire N__78618;
    wire N__78617;
    wire N__78616;
    wire N__78615;
    wire N__78614;
    wire N__78613;
    wire N__78612;
    wire N__78611;
    wire N__78610;
    wire N__78609;
    wire N__78608;
    wire N__78607;
    wire N__78606;
    wire N__78605;
    wire N__78604;
    wire N__78603;
    wire N__78602;
    wire N__78601;
    wire N__78600;
    wire N__78599;
    wire N__78598;
    wire N__78597;
    wire N__78596;
    wire N__78595;
    wire N__78594;
    wire N__78593;
    wire N__78592;
    wire N__78591;
    wire N__78590;
    wire N__78589;
    wire N__78588;
    wire N__78587;
    wire N__78586;
    wire N__78585;
    wire N__78584;
    wire N__78583;
    wire N__78582;
    wire N__78581;
    wire N__78580;
    wire N__78579;
    wire N__78578;
    wire N__78577;
    wire N__78576;
    wire N__78575;
    wire N__78574;
    wire N__78573;
    wire N__78572;
    wire N__78571;
    wire N__78570;
    wire N__78569;
    wire N__78568;
    wire N__78567;
    wire N__78566;
    wire N__78565;
    wire N__78564;
    wire N__78563;
    wire N__78562;
    wire N__78033;
    wire N__78030;
    wire N__78027;
    wire N__78026;
    wire N__78025;
    wire N__78024;
    wire N__78021;
    wire N__78020;
    wire N__78019;
    wire N__78018;
    wire N__78017;
    wire N__78014;
    wire N__78009;
    wire N__78006;
    wire N__78003;
    wire N__77998;
    wire N__77995;
    wire N__77992;
    wire N__77987;
    wire N__77982;
    wire N__77979;
    wire N__77976;
    wire N__77971;
    wire N__77966;
    wire N__77963;
    wire N__77958;
    wire N__77957;
    wire N__77956;
    wire N__77955;
    wire N__77954;
    wire N__77951;
    wire N__77948;
    wire N__77945;
    wire N__77942;
    wire N__77939;
    wire N__77938;
    wire N__77933;
    wire N__77928;
    wire N__77925;
    wire N__77922;
    wire N__77919;
    wire N__77914;
    wire N__77911;
    wire N__77906;
    wire N__77903;
    wire N__77898;
    wire N__77895;
    wire N__77892;
    wire N__77889;
    wire N__77886;
    wire N__77883;
    wire N__77880;
    wire N__77879;
    wire N__77876;
    wire N__77873;
    wire N__77872;
    wire N__77869;
    wire N__77866;
    wire N__77863;
    wire N__77858;
    wire N__77857;
    wire N__77856;
    wire N__77853;
    wire N__77850;
    wire N__77847;
    wire N__77846;
    wire N__77845;
    wire N__77844;
    wire N__77841;
    wire N__77838;
    wire N__77833;
    wire N__77826;
    wire N__77817;
    wire N__77816;
    wire N__77813;
    wire N__77812;
    wire N__77811;
    wire N__77810;
    wire N__77807;
    wire N__77804;
    wire N__77799;
    wire N__77796;
    wire N__77793;
    wire N__77792;
    wire N__77789;
    wire N__77784;
    wire N__77781;
    wire N__77778;
    wire N__77777;
    wire N__77776;
    wire N__77771;
    wire N__77766;
    wire N__77761;
    wire N__77754;
    wire N__77751;
    wire N__77748;
    wire N__77745;
    wire N__77742;
    wire N__77739;
    wire N__77736;
    wire N__77733;
    wire N__77730;
    wire N__77727;
    wire N__77726;
    wire N__77723;
    wire N__77720;
    wire N__77715;
    wire N__77712;
    wire N__77709;
    wire N__77706;
    wire N__77705;
    wire N__77702;
    wire N__77699;
    wire N__77696;
    wire N__77693;
    wire N__77688;
    wire N__77687;
    wire N__77684;
    wire N__77681;
    wire N__77678;
    wire N__77675;
    wire N__77674;
    wire N__77673;
    wire N__77668;
    wire N__77663;
    wire N__77658;
    wire N__77655;
    wire N__77654;
    wire N__77651;
    wire N__77650;
    wire N__77649;
    wire N__77646;
    wire N__77643;
    wire N__77640;
    wire N__77639;
    wire N__77638;
    wire N__77635;
    wire N__77632;
    wire N__77629;
    wire N__77626;
    wire N__77623;
    wire N__77620;
    wire N__77617;
    wire N__77614;
    wire N__77611;
    wire N__77608;
    wire N__77605;
    wire N__77602;
    wire N__77593;
    wire N__77590;
    wire N__77583;
    wire N__77580;
    wire N__77579;
    wire N__77578;
    wire N__77575;
    wire N__77574;
    wire N__77573;
    wire N__77570;
    wire N__77569;
    wire N__77566;
    wire N__77563;
    wire N__77560;
    wire N__77557;
    wire N__77554;
    wire N__77551;
    wire N__77546;
    wire N__77543;
    wire N__77538;
    wire N__77535;
    wire N__77532;
    wire N__77529;
    wire N__77526;
    wire N__77517;
    wire N__77514;
    wire N__77511;
    wire N__77508;
    wire N__77505;
    wire N__77502;
    wire N__77501;
    wire N__77498;
    wire N__77495;
    wire N__77490;
    wire N__77489;
    wire N__77486;
    wire N__77483;
    wire N__77480;
    wire N__77477;
    wire N__77474;
    wire N__77471;
    wire N__77466;
    wire N__77463;
    wire N__77460;
    wire N__77457;
    wire N__77454;
    wire N__77453;
    wire N__77450;
    wire N__77447;
    wire N__77446;
    wire N__77441;
    wire N__77440;
    wire N__77437;
    wire N__77434;
    wire N__77431;
    wire N__77428;
    wire N__77421;
    wire N__77418;
    wire N__77417;
    wire N__77414;
    wire N__77411;
    wire N__77406;
    wire N__77405;
    wire N__77402;
    wire N__77399;
    wire N__77394;
    wire N__77393;
    wire N__77392;
    wire N__77391;
    wire N__77388;
    wire N__77383;
    wire N__77380;
    wire N__77377;
    wire N__77376;
    wire N__77373;
    wire N__77368;
    wire N__77365;
    wire N__77362;
    wire N__77355;
    wire N__77352;
    wire N__77351;
    wire N__77348;
    wire N__77345;
    wire N__77342;
    wire N__77341;
    wire N__77336;
    wire N__77333;
    wire N__77332;
    wire N__77329;
    wire N__77326;
    wire N__77323;
    wire N__77318;
    wire N__77315;
    wire N__77312;
    wire N__77307;
    wire N__77304;
    wire N__77301;
    wire N__77298;
    wire N__77295;
    wire N__77292;
    wire N__77291;
    wire N__77288;
    wire N__77287;
    wire N__77284;
    wire N__77281;
    wire N__77280;
    wire N__77277;
    wire N__77274;
    wire N__77273;
    wire N__77270;
    wire N__77267;
    wire N__77266;
    wire N__77261;
    wire N__77258;
    wire N__77255;
    wire N__77252;
    wire N__77249;
    wire N__77246;
    wire N__77243;
    wire N__77238;
    wire N__77229;
    wire N__77226;
    wire N__77223;
    wire N__77220;
    wire N__77217;
    wire N__77216;
    wire N__77213;
    wire N__77210;
    wire N__77209;
    wire N__77204;
    wire N__77201;
    wire N__77198;
    wire N__77195;
    wire N__77190;
    wire N__77189;
    wire N__77188;
    wire N__77187;
    wire N__77184;
    wire N__77181;
    wire N__77180;
    wire N__77177;
    wire N__77174;
    wire N__77171;
    wire N__77168;
    wire N__77165;
    wire N__77162;
    wire N__77151;
    wire N__77150;
    wire N__77147;
    wire N__77144;
    wire N__77141;
    wire N__77138;
    wire N__77133;
    wire N__77132;
    wire N__77131;
    wire N__77130;
    wire N__77129;
    wire N__77128;
    wire N__77125;
    wire N__77124;
    wire N__77123;
    wire N__77122;
    wire N__77121;
    wire N__77118;
    wire N__77115;
    wire N__77112;
    wire N__77111;
    wire N__77110;
    wire N__77107;
    wire N__77106;
    wire N__77103;
    wire N__77102;
    wire N__77101;
    wire N__77100;
    wire N__77099;
    wire N__77098;
    wire N__77093;
    wire N__77092;
    wire N__77091;
    wire N__77090;
    wire N__77087;
    wire N__77084;
    wire N__77081;
    wire N__77078;
    wire N__77075;
    wire N__77072;
    wire N__77069;
    wire N__77066;
    wire N__77065;
    wire N__77062;
    wire N__77059;
    wire N__77058;
    wire N__77055;
    wire N__77052;
    wire N__77049;
    wire N__77046;
    wire N__77045;
    wire N__77044;
    wire N__77041;
    wire N__77038;
    wire N__77035;
    wire N__77028;
    wire N__77023;
    wire N__77020;
    wire N__77017;
    wire N__77012;
    wire N__77009;
    wire N__77006;
    wire N__77003;
    wire N__76998;
    wire N__76997;
    wire N__76994;
    wire N__76985;
    wire N__76982;
    wire N__76979;
    wire N__76974;
    wire N__76963;
    wire N__76958;
    wire N__76955;
    wire N__76954;
    wire N__76949;
    wire N__76946;
    wire N__76945;
    wire N__76944;
    wire N__76941;
    wire N__76936;
    wire N__76933;
    wire N__76926;
    wire N__76923;
    wire N__76920;
    wire N__76917;
    wire N__76916;
    wire N__76913;
    wire N__76912;
    wire N__76909;
    wire N__76906;
    wire N__76903;
    wire N__76900;
    wire N__76895;
    wire N__76892;
    wire N__76887;
    wire N__76884;
    wire N__76883;
    wire N__76880;
    wire N__76877;
    wire N__76874;
    wire N__76865;
    wire N__76860;
    wire N__76855;
    wire N__76852;
    wire N__76845;
    wire N__76842;
    wire N__76833;
    wire N__76832;
    wire N__76829;
    wire N__76828;
    wire N__76825;
    wire N__76822;
    wire N__76819;
    wire N__76816;
    wire N__76815;
    wire N__76810;
    wire N__76807;
    wire N__76804;
    wire N__76801;
    wire N__76798;
    wire N__76797;
    wire N__76794;
    wire N__76791;
    wire N__76788;
    wire N__76785;
    wire N__76776;
    wire N__76773;
    wire N__76770;
    wire N__76767;
    wire N__76764;
    wire N__76761;
    wire N__76758;
    wire N__76755;
    wire N__76752;
    wire N__76749;
    wire N__76746;
    wire N__76743;
    wire N__76742;
    wire N__76741;
    wire N__76738;
    wire N__76735;
    wire N__76732;
    wire N__76727;
    wire N__76726;
    wire N__76723;
    wire N__76720;
    wire N__76717;
    wire N__76710;
    wire N__76707;
    wire N__76704;
    wire N__76701;
    wire N__76698;
    wire N__76695;
    wire N__76694;
    wire N__76693;
    wire N__76688;
    wire N__76687;
    wire N__76684;
    wire N__76683;
    wire N__76682;
    wire N__76679;
    wire N__76676;
    wire N__76675;
    wire N__76674;
    wire N__76671;
    wire N__76668;
    wire N__76665;
    wire N__76660;
    wire N__76657;
    wire N__76656;
    wire N__76655;
    wire N__76654;
    wire N__76653;
    wire N__76652;
    wire N__76649;
    wire N__76644;
    wire N__76641;
    wire N__76636;
    wire N__76631;
    wire N__76630;
    wire N__76629;
    wire N__76626;
    wire N__76625;
    wire N__76624;
    wire N__76623;
    wire N__76622;
    wire N__76617;
    wire N__76614;
    wire N__76613;
    wire N__76612;
    wire N__76611;
    wire N__76610;
    wire N__76607;
    wire N__76600;
    wire N__76599;
    wire N__76596;
    wire N__76595;
    wire N__76592;
    wire N__76589;
    wire N__76586;
    wire N__76583;
    wire N__76582;
    wire N__76579;
    wire N__76576;
    wire N__76573;
    wire N__76570;
    wire N__76567;
    wire N__76564;
    wire N__76559;
    wire N__76554;
    wire N__76551;
    wire N__76550;
    wire N__76549;
    wire N__76548;
    wire N__76545;
    wire N__76542;
    wire N__76539;
    wire N__76536;
    wire N__76531;
    wire N__76530;
    wire N__76529;
    wire N__76526;
    wire N__76525;
    wire N__76520;
    wire N__76513;
    wire N__76510;
    wire N__76505;
    wire N__76502;
    wire N__76499;
    wire N__76496;
    wire N__76493;
    wire N__76484;
    wire N__76481;
    wire N__76478;
    wire N__76475;
    wire N__76472;
    wire N__76469;
    wire N__76464;
    wire N__76459;
    wire N__76456;
    wire N__76449;
    wire N__76446;
    wire N__76443;
    wire N__76434;
    wire N__76429;
    wire N__76426;
    wire N__76423;
    wire N__76420;
    wire N__76417;
    wire N__76414;
    wire N__76411;
    wire N__76398;
    wire N__76395;
    wire N__76394;
    wire N__76393;
    wire N__76390;
    wire N__76389;
    wire N__76386;
    wire N__76385;
    wire N__76384;
    wire N__76383;
    wire N__76382;
    wire N__76379;
    wire N__76378;
    wire N__76375;
    wire N__76372;
    wire N__76369;
    wire N__76366;
    wire N__76365;
    wire N__76362;
    wire N__76359;
    wire N__76356;
    wire N__76355;
    wire N__76354;
    wire N__76351;
    wire N__76348;
    wire N__76343;
    wire N__76338;
    wire N__76335;
    wire N__76332;
    wire N__76329;
    wire N__76326;
    wire N__76325;
    wire N__76324;
    wire N__76321;
    wire N__76318;
    wire N__76317;
    wire N__76316;
    wire N__76315;
    wire N__76310;
    wire N__76305;
    wire N__76302;
    wire N__76295;
    wire N__76294;
    wire N__76293;
    wire N__76290;
    wire N__76289;
    wire N__76286;
    wire N__76285;
    wire N__76282;
    wire N__76279;
    wire N__76276;
    wire N__76275;
    wire N__76274;
    wire N__76271;
    wire N__76268;
    wire N__76265;
    wire N__76260;
    wire N__76257;
    wire N__76254;
    wire N__76251;
    wire N__76248;
    wire N__76245;
    wire N__76242;
    wire N__76239;
    wire N__76232;
    wire N__76229;
    wire N__76228;
    wire N__76227;
    wire N__76224;
    wire N__76221;
    wire N__76218;
    wire N__76215;
    wire N__76212;
    wire N__76209;
    wire N__76206;
    wire N__76199;
    wire N__76194;
    wire N__76191;
    wire N__76188;
    wire N__76183;
    wire N__76180;
    wire N__76175;
    wire N__76172;
    wire N__76167;
    wire N__76164;
    wire N__76161;
    wire N__76158;
    wire N__76155;
    wire N__76154;
    wire N__76153;
    wire N__76152;
    wire N__76151;
    wire N__76150;
    wire N__76149;
    wire N__76148;
    wire N__76135;
    wire N__76130;
    wire N__76125;
    wire N__76122;
    wire N__76117;
    wire N__76112;
    wire N__76107;
    wire N__76104;
    wire N__76099;
    wire N__76086;
    wire N__76083;
    wire N__76082;
    wire N__76079;
    wire N__76076;
    wire N__76071;
    wire N__76070;
    wire N__76067;
    wire N__76064;
    wire N__76061;
    wire N__76058;
    wire N__76053;
    wire N__76052;
    wire N__76049;
    wire N__76048;
    wire N__76047;
    wire N__76044;
    wire N__76041;
    wire N__76038;
    wire N__76037;
    wire N__76036;
    wire N__76033;
    wire N__76030;
    wire N__76027;
    wire N__76022;
    wire N__76019;
    wire N__76016;
    wire N__76013;
    wire N__76008;
    wire N__76005;
    wire N__75996;
    wire N__75993;
    wire N__75990;
    wire N__75989;
    wire N__75986;
    wire N__75983;
    wire N__75980;
    wire N__75977;
    wire N__75974;
    wire N__75969;
    wire N__75966;
    wire N__75963;
    wire N__75962;
    wire N__75959;
    wire N__75956;
    wire N__75951;
    wire N__75948;
    wire N__75947;
    wire N__75946;
    wire N__75943;
    wire N__75940;
    wire N__75939;
    wire N__75938;
    wire N__75935;
    wire N__75932;
    wire N__75929;
    wire N__75926;
    wire N__75923;
    wire N__75920;
    wire N__75913;
    wire N__75910;
    wire N__75909;
    wire N__75906;
    wire N__75903;
    wire N__75900;
    wire N__75897;
    wire N__75894;
    wire N__75891;
    wire N__75888;
    wire N__75883;
    wire N__75880;
    wire N__75873;
    wire N__75870;
    wire N__75867;
    wire N__75864;
    wire N__75861;
    wire N__75858;
    wire N__75857;
    wire N__75854;
    wire N__75851;
    wire N__75848;
    wire N__75847;
    wire N__75844;
    wire N__75841;
    wire N__75838;
    wire N__75831;
    wire N__75830;
    wire N__75827;
    wire N__75824;
    wire N__75823;
    wire N__75820;
    wire N__75815;
    wire N__75810;
    wire N__75807;
    wire N__75804;
    wire N__75801;
    wire N__75798;
    wire N__75795;
    wire N__75792;
    wire N__75789;
    wire N__75786;
    wire N__75785;
    wire N__75784;
    wire N__75779;
    wire N__75778;
    wire N__75775;
    wire N__75772;
    wire N__75769;
    wire N__75766;
    wire N__75765;
    wire N__75762;
    wire N__75757;
    wire N__75754;
    wire N__75751;
    wire N__75748;
    wire N__75745;
    wire N__75742;
    wire N__75739;
    wire N__75732;
    wire N__75731;
    wire N__75730;
    wire N__75729;
    wire N__75726;
    wire N__75719;
    wire N__75716;
    wire N__75713;
    wire N__75708;
    wire N__75705;
    wire N__75702;
    wire N__75701;
    wire N__75700;
    wire N__75697;
    wire N__75694;
    wire N__75691;
    wire N__75688;
    wire N__75685;
    wire N__75682;
    wire N__75679;
    wire N__75678;
    wire N__75675;
    wire N__75672;
    wire N__75669;
    wire N__75666;
    wire N__75663;
    wire N__75660;
    wire N__75657;
    wire N__75654;
    wire N__75649;
    wire N__75646;
    wire N__75641;
    wire N__75636;
    wire N__75633;
    wire N__75630;
    wire N__75627;
    wire N__75624;
    wire N__75621;
    wire N__75620;
    wire N__75615;
    wire N__75614;
    wire N__75613;
    wire N__75612;
    wire N__75611;
    wire N__75608;
    wire N__75605;
    wire N__75600;
    wire N__75597;
    wire N__75590;
    wire N__75587;
    wire N__75584;
    wire N__75579;
    wire N__75576;
    wire N__75573;
    wire N__75570;
    wire N__75567;
    wire N__75566;
    wire N__75563;
    wire N__75562;
    wire N__75559;
    wire N__75558;
    wire N__75555;
    wire N__75554;
    wire N__75553;
    wire N__75550;
    wire N__75549;
    wire N__75548;
    wire N__75545;
    wire N__75542;
    wire N__75539;
    wire N__75536;
    wire N__75533;
    wire N__75528;
    wire N__75525;
    wire N__75522;
    wire N__75507;
    wire N__75506;
    wire N__75501;
    wire N__75500;
    wire N__75499;
    wire N__75498;
    wire N__75495;
    wire N__75494;
    wire N__75493;
    wire N__75492;
    wire N__75489;
    wire N__75484;
    wire N__75481;
    wire N__75476;
    wire N__75473;
    wire N__75470;
    wire N__75467;
    wire N__75464;
    wire N__75461;
    wire N__75458;
    wire N__75455;
    wire N__75452;
    wire N__75449;
    wire N__75442;
    wire N__75439;
    wire N__75436;
    wire N__75433;
    wire N__75426;
    wire N__75423;
    wire N__75422;
    wire N__75421;
    wire N__75420;
    wire N__75417;
    wire N__75416;
    wire N__75415;
    wire N__75408;
    wire N__75407;
    wire N__75406;
    wire N__75403;
    wire N__75400;
    wire N__75399;
    wire N__75398;
    wire N__75397;
    wire N__75394;
    wire N__75393;
    wire N__75390;
    wire N__75385;
    wire N__75380;
    wire N__75375;
    wire N__75374;
    wire N__75373;
    wire N__75370;
    wire N__75367;
    wire N__75364;
    wire N__75359;
    wire N__75356;
    wire N__75353;
    wire N__75350;
    wire N__75347;
    wire N__75344;
    wire N__75341;
    wire N__75338;
    wire N__75337;
    wire N__75334;
    wire N__75331;
    wire N__75328;
    wire N__75327;
    wire N__75326;
    wire N__75321;
    wire N__75318;
    wire N__75313;
    wire N__75310;
    wire N__75307;
    wire N__75302;
    wire N__75301;
    wire N__75298;
    wire N__75295;
    wire N__75290;
    wire N__75287;
    wire N__75280;
    wire N__75277;
    wire N__75274;
    wire N__75261;
    wire N__75258;
    wire N__75257;
    wire N__75256;
    wire N__75255;
    wire N__75254;
    wire N__75253;
    wire N__75252;
    wire N__75251;
    wire N__75250;
    wire N__75249;
    wire N__75248;
    wire N__75245;
    wire N__75244;
    wire N__75243;
    wire N__75242;
    wire N__75239;
    wire N__75236;
    wire N__75233;
    wire N__75230;
    wire N__75229;
    wire N__75228;
    wire N__75225;
    wire N__75224;
    wire N__75219;
    wire N__75216;
    wire N__75211;
    wire N__75208;
    wire N__75205;
    wire N__75202;
    wire N__75199;
    wire N__75196;
    wire N__75195;
    wire N__75190;
    wire N__75187;
    wire N__75186;
    wire N__75185;
    wire N__75182;
    wire N__75179;
    wire N__75178;
    wire N__75177;
    wire N__75174;
    wire N__75171;
    wire N__75166;
    wire N__75163;
    wire N__75160;
    wire N__75153;
    wire N__75150;
    wire N__75147;
    wire N__75142;
    wire N__75139;
    wire N__75138;
    wire N__75137;
    wire N__75134;
    wire N__75131;
    wire N__75128;
    wire N__75125;
    wire N__75122;
    wire N__75117;
    wire N__75114;
    wire N__75113;
    wire N__75112;
    wire N__75111;
    wire N__75110;
    wire N__75103;
    wire N__75098;
    wire N__75093;
    wire N__75088;
    wire N__75085;
    wire N__75080;
    wire N__75077;
    wire N__75074;
    wire N__75071;
    wire N__75068;
    wire N__75065;
    wire N__75062;
    wire N__75057;
    wire N__75054;
    wire N__75051;
    wire N__75048;
    wire N__75047;
    wire N__75046;
    wire N__75041;
    wire N__75034;
    wire N__75029;
    wire N__75028;
    wire N__75027;
    wire N__75022;
    wire N__75019;
    wire N__75012;
    wire N__75007;
    wire N__75002;
    wire N__74999;
    wire N__74996;
    wire N__74993;
    wire N__74990;
    wire N__74987;
    wire N__74984;
    wire N__74977;
    wire N__74964;
    wire N__74963;
    wire N__74962;
    wire N__74961;
    wire N__74958;
    wire N__74955;
    wire N__74952;
    wire N__74949;
    wire N__74946;
    wire N__74943;
    wire N__74940;
    wire N__74937;
    wire N__74934;
    wire N__74933;
    wire N__74930;
    wire N__74927;
    wire N__74922;
    wire N__74919;
    wire N__74914;
    wire N__74911;
    wire N__74904;
    wire N__74903;
    wire N__74900;
    wire N__74897;
    wire N__74894;
    wire N__74893;
    wire N__74890;
    wire N__74887;
    wire N__74884;
    wire N__74881;
    wire N__74874;
    wire N__74871;
    wire N__74870;
    wire N__74867;
    wire N__74866;
    wire N__74863;
    wire N__74860;
    wire N__74857;
    wire N__74854;
    wire N__74851;
    wire N__74848;
    wire N__74841;
    wire N__74838;
    wire N__74837;
    wire N__74834;
    wire N__74831;
    wire N__74828;
    wire N__74825;
    wire N__74822;
    wire N__74817;
    wire N__74816;
    wire N__74815;
    wire N__74812;
    wire N__74811;
    wire N__74808;
    wire N__74805;
    wire N__74802;
    wire N__74799;
    wire N__74794;
    wire N__74789;
    wire N__74786;
    wire N__74783;
    wire N__74778;
    wire N__74775;
    wire N__74774;
    wire N__74773;
    wire N__74772;
    wire N__74769;
    wire N__74768;
    wire N__74765;
    wire N__74760;
    wire N__74757;
    wire N__74752;
    wire N__74745;
    wire N__74742;
    wire N__74739;
    wire N__74736;
    wire N__74733;
    wire N__74730;
    wire N__74727;
    wire N__74724;
    wire N__74721;
    wire N__74718;
    wire N__74715;
    wire N__74714;
    wire N__74713;
    wire N__74712;
    wire N__74709;
    wire N__74704;
    wire N__74701;
    wire N__74698;
    wire N__74695;
    wire N__74692;
    wire N__74689;
    wire N__74686;
    wire N__74679;
    wire N__74678;
    wire N__74675;
    wire N__74674;
    wire N__74673;
    wire N__74670;
    wire N__74667;
    wire N__74666;
    wire N__74663;
    wire N__74660;
    wire N__74659;
    wire N__74658;
    wire N__74655;
    wire N__74652;
    wire N__74647;
    wire N__74644;
    wire N__74643;
    wire N__74642;
    wire N__74637;
    wire N__74636;
    wire N__74633;
    wire N__74632;
    wire N__74631;
    wire N__74626;
    wire N__74625;
    wire N__74622;
    wire N__74619;
    wire N__74616;
    wire N__74613;
    wire N__74610;
    wire N__74607;
    wire N__74604;
    wire N__74601;
    wire N__74598;
    wire N__74595;
    wire N__74592;
    wire N__74589;
    wire N__74586;
    wire N__74581;
    wire N__74578;
    wire N__74573;
    wire N__74570;
    wire N__74563;
    wire N__74562;
    wire N__74559;
    wire N__74556;
    wire N__74553;
    wire N__74548;
    wire N__74545;
    wire N__74542;
    wire N__74529;
    wire N__74526;
    wire N__74525;
    wire N__74524;
    wire N__74521;
    wire N__74520;
    wire N__74517;
    wire N__74514;
    wire N__74511;
    wire N__74508;
    wire N__74507;
    wire N__74504;
    wire N__74501;
    wire N__74500;
    wire N__74499;
    wire N__74498;
    wire N__74493;
    wire N__74490;
    wire N__74487;
    wire N__74484;
    wire N__74481;
    wire N__74480;
    wire N__74477;
    wire N__74474;
    wire N__74471;
    wire N__74470;
    wire N__74469;
    wire N__74466;
    wire N__74459;
    wire N__74456;
    wire N__74453;
    wire N__74448;
    wire N__74447;
    wire N__74442;
    wire N__74441;
    wire N__74436;
    wire N__74429;
    wire N__74426;
    wire N__74423;
    wire N__74420;
    wire N__74417;
    wire N__74414;
    wire N__74407;
    wire N__74406;
    wire N__74403;
    wire N__74398;
    wire N__74395;
    wire N__74388;
    wire N__74387;
    wire N__74386;
    wire N__74383;
    wire N__74382;
    wire N__74381;
    wire N__74378;
    wire N__74375;
    wire N__74372;
    wire N__74369;
    wire N__74366;
    wire N__74365;
    wire N__74362;
    wire N__74359;
    wire N__74358;
    wire N__74355;
    wire N__74352;
    wire N__74349;
    wire N__74348;
    wire N__74345;
    wire N__74344;
    wire N__74341;
    wire N__74338;
    wire N__74335;
    wire N__74332;
    wire N__74329;
    wire N__74326;
    wire N__74323;
    wire N__74320;
    wire N__74317;
    wire N__74312;
    wire N__74309;
    wire N__74306;
    wire N__74303;
    wire N__74302;
    wire N__74297;
    wire N__74292;
    wire N__74289;
    wire N__74288;
    wire N__74285;
    wire N__74280;
    wire N__74279;
    wire N__74276;
    wire N__74273;
    wire N__74270;
    wire N__74267;
    wire N__74264;
    wire N__74259;
    wire N__74256;
    wire N__74247;
    wire N__74242;
    wire N__74239;
    wire N__74238;
    wire N__74235;
    wire N__74230;
    wire N__74227;
    wire N__74220;
    wire N__74217;
    wire N__74216;
    wire N__74213;
    wire N__74210;
    wire N__74209;
    wire N__74208;
    wire N__74207;
    wire N__74206;
    wire N__74205;
    wire N__74204;
    wire N__74203;
    wire N__74202;
    wire N__74197;
    wire N__74194;
    wire N__74189;
    wire N__74188;
    wire N__74187;
    wire N__74184;
    wire N__74181;
    wire N__74180;
    wire N__74179;
    wire N__74178;
    wire N__74171;
    wire N__74166;
    wire N__74163;
    wire N__74158;
    wire N__74157;
    wire N__74156;
    wire N__74151;
    wire N__74150;
    wire N__74147;
    wire N__74146;
    wire N__74145;
    wire N__74142;
    wire N__74139;
    wire N__74136;
    wire N__74135;
    wire N__74132;
    wire N__74127;
    wire N__74124;
    wire N__74121;
    wire N__74118;
    wire N__74117;
    wire N__74116;
    wire N__74115;
    wire N__74112;
    wire N__74111;
    wire N__74108;
    wire N__74105;
    wire N__74104;
    wire N__74101;
    wire N__74098;
    wire N__74095;
    wire N__74092;
    wire N__74089;
    wire N__74086;
    wire N__74081;
    wire N__74076;
    wire N__74073;
    wire N__74070;
    wire N__74069;
    wire N__74068;
    wire N__74067;
    wire N__74066;
    wire N__74063;
    wire N__74060;
    wire N__74057;
    wire N__74052;
    wire N__74051;
    wire N__74048;
    wire N__74045;
    wire N__74040;
    wire N__74035;
    wire N__74030;
    wire N__74025;
    wire N__74022;
    wire N__74021;
    wire N__74018;
    wire N__74015;
    wire N__74010;
    wire N__74003;
    wire N__74000;
    wire N__73997;
    wire N__73990;
    wire N__73981;
    wire N__73978;
    wire N__73975;
    wire N__73972;
    wire N__73967;
    wire N__73964;
    wire N__73957;
    wire N__73944;
    wire N__73943;
    wire N__73940;
    wire N__73939;
    wire N__73936;
    wire N__73933;
    wire N__73930;
    wire N__73927;
    wire N__73924;
    wire N__73921;
    wire N__73918;
    wire N__73915;
    wire N__73908;
    wire N__73905;
    wire N__73902;
    wire N__73901;
    wire N__73900;
    wire N__73899;
    wire N__73896;
    wire N__73893;
    wire N__73890;
    wire N__73887;
    wire N__73884;
    wire N__73881;
    wire N__73876;
    wire N__73873;
    wire N__73868;
    wire N__73863;
    wire N__73862;
    wire N__73861;
    wire N__73858;
    wire N__73855;
    wire N__73854;
    wire N__73851;
    wire N__73848;
    wire N__73843;
    wire N__73840;
    wire N__73837;
    wire N__73834;
    wire N__73831;
    wire N__73828;
    wire N__73825;
    wire N__73822;
    wire N__73817;
    wire N__73814;
    wire N__73809;
    wire N__73806;
    wire N__73803;
    wire N__73800;
    wire N__73797;
    wire N__73796;
    wire N__73793;
    wire N__73790;
    wire N__73787;
    wire N__73784;
    wire N__73779;
    wire N__73776;
    wire N__73773;
    wire N__73772;
    wire N__73769;
    wire N__73766;
    wire N__73763;
    wire N__73760;
    wire N__73755;
    wire N__73752;
    wire N__73751;
    wire N__73750;
    wire N__73747;
    wire N__73744;
    wire N__73741;
    wire N__73738;
    wire N__73735;
    wire N__73734;
    wire N__73727;
    wire N__73724;
    wire N__73719;
    wire N__73718;
    wire N__73717;
    wire N__73716;
    wire N__73715;
    wire N__73714;
    wire N__73711;
    wire N__73710;
    wire N__73709;
    wire N__73708;
    wire N__73707;
    wire N__73706;
    wire N__73705;
    wire N__73704;
    wire N__73703;
    wire N__73702;
    wire N__73697;
    wire N__73696;
    wire N__73695;
    wire N__73694;
    wire N__73693;
    wire N__73692;
    wire N__73691;
    wire N__73690;
    wire N__73689;
    wire N__73688;
    wire N__73687;
    wire N__73686;
    wire N__73685;
    wire N__73684;
    wire N__73681;
    wire N__73670;
    wire N__73669;
    wire N__73668;
    wire N__73667;
    wire N__73666;
    wire N__73665;
    wire N__73662;
    wire N__73659;
    wire N__73658;
    wire N__73655;
    wire N__73652;
    wire N__73651;
    wire N__73644;
    wire N__73641;
    wire N__73630;
    wire N__73623;
    wire N__73620;
    wire N__73615;
    wire N__73612;
    wire N__73611;
    wire N__73610;
    wire N__73609;
    wire N__73608;
    wire N__73605;
    wire N__73602;
    wire N__73599;
    wire N__73598;
    wire N__73597;
    wire N__73596;
    wire N__73595;
    wire N__73590;
    wire N__73587;
    wire N__73582;
    wire N__73579;
    wire N__73576;
    wire N__73573;
    wire N__73570;
    wire N__73567;
    wire N__73564;
    wire N__73561;
    wire N__73558;
    wire N__73551;
    wire N__73548;
    wire N__73543;
    wire N__73534;
    wire N__73529;
    wire N__73526;
    wire N__73523;
    wire N__73522;
    wire N__73521;
    wire N__73520;
    wire N__73519;
    wire N__73518;
    wire N__73513;
    wire N__73506;
    wire N__73503;
    wire N__73500;
    wire N__73497;
    wire N__73492;
    wire N__73489;
    wire N__73484;
    wire N__73479;
    wire N__73472;
    wire N__73467;
    wire N__73464;
    wire N__73461;
    wire N__73458;
    wire N__73453;
    wire N__73450;
    wire N__73447;
    wire N__73444;
    wire N__73441;
    wire N__73436;
    wire N__73431;
    wire N__73424;
    wire N__73401;
    wire N__73400;
    wire N__73397;
    wire N__73396;
    wire N__73393;
    wire N__73392;
    wire N__73389;
    wire N__73386;
    wire N__73383;
    wire N__73380;
    wire N__73377;
    wire N__73374;
    wire N__73369;
    wire N__73366;
    wire N__73361;
    wire N__73356;
    wire N__73353;
    wire N__73350;
    wire N__73349;
    wire N__73348;
    wire N__73347;
    wire N__73346;
    wire N__73343;
    wire N__73338;
    wire N__73337;
    wire N__73336;
    wire N__73335;
    wire N__73332;
    wire N__73331;
    wire N__73330;
    wire N__73327;
    wire N__73326;
    wire N__73321;
    wire N__73316;
    wire N__73313;
    wire N__73308;
    wire N__73307;
    wire N__73304;
    wire N__73301;
    wire N__73300;
    wire N__73299;
    wire N__73298;
    wire N__73295;
    wire N__73294;
    wire N__73293;
    wire N__73292;
    wire N__73291;
    wire N__73290;
    wire N__73289;
    wire N__73286;
    wire N__73283;
    wire N__73280;
    wire N__73277;
    wire N__73276;
    wire N__73273;
    wire N__73270;
    wire N__73267;
    wire N__73264;
    wire N__73261;
    wire N__73258;
    wire N__73255;
    wire N__73250;
    wire N__73245;
    wire N__73242;
    wire N__73239;
    wire N__73234;
    wire N__73229;
    wire N__73226;
    wire N__73223;
    wire N__73220;
    wire N__73215;
    wire N__73214;
    wire N__73211;
    wire N__73210;
    wire N__73209;
    wire N__73208;
    wire N__73207;
    wire N__73202;
    wire N__73201;
    wire N__73196;
    wire N__73187;
    wire N__73182;
    wire N__73179;
    wire N__73176;
    wire N__73173;
    wire N__73170;
    wire N__73167;
    wire N__73160;
    wire N__73157;
    wire N__73156;
    wire N__73155;
    wire N__73154;
    wire N__73153;
    wire N__73150;
    wire N__73147;
    wire N__73144;
    wire N__73137;
    wire N__73134;
    wire N__73131;
    wire N__73124;
    wire N__73121;
    wire N__73118;
    wire N__73113;
    wire N__73110;
    wire N__73103;
    wire N__73096;
    wire N__73083;
    wire N__73082;
    wire N__73081;
    wire N__73078;
    wire N__73075;
    wire N__73072;
    wire N__73067;
    wire N__73064;
    wire N__73059;
    wire N__73056;
    wire N__73055;
    wire N__73052;
    wire N__73049;
    wire N__73046;
    wire N__73043;
    wire N__73038;
    wire N__73035;
    wire N__73034;
    wire N__73033;
    wire N__73030;
    wire N__73027;
    wire N__73024;
    wire N__73021;
    wire N__73020;
    wire N__73015;
    wire N__73012;
    wire N__73009;
    wire N__73006;
    wire N__73003;
    wire N__72996;
    wire N__72993;
    wire N__72992;
    wire N__72991;
    wire N__72990;
    wire N__72989;
    wire N__72986;
    wire N__72983;
    wire N__72982;
    wire N__72981;
    wire N__72980;
    wire N__72979;
    wire N__72978;
    wire N__72977;
    wire N__72974;
    wire N__72971;
    wire N__72968;
    wire N__72967;
    wire N__72966;
    wire N__72965;
    wire N__72964;
    wire N__72961;
    wire N__72956;
    wire N__72949;
    wire N__72946;
    wire N__72943;
    wire N__72942;
    wire N__72941;
    wire N__72940;
    wire N__72939;
    wire N__72938;
    wire N__72937;
    wire N__72936;
    wire N__72935;
    wire N__72932;
    wire N__72929;
    wire N__72926;
    wire N__72925;
    wire N__72924;
    wire N__72923;
    wire N__72920;
    wire N__72917;
    wire N__72912;
    wire N__72909;
    wire N__72906;
    wire N__72903;
    wire N__72900;
    wire N__72899;
    wire N__72898;
    wire N__72893;
    wire N__72890;
    wire N__72887;
    wire N__72884;
    wire N__72881;
    wire N__72880;
    wire N__72875;
    wire N__72872;
    wire N__72869;
    wire N__72866;
    wire N__72863;
    wire N__72862;
    wire N__72861;
    wire N__72860;
    wire N__72857;
    wire N__72848;
    wire N__72845;
    wire N__72838;
    wire N__72835;
    wire N__72832;
    wire N__72829;
    wire N__72826;
    wire N__72821;
    wire N__72816;
    wire N__72813;
    wire N__72810;
    wire N__72805;
    wire N__72800;
    wire N__72797;
    wire N__72792;
    wire N__72789;
    wire N__72786;
    wire N__72781;
    wire N__72774;
    wire N__72771;
    wire N__72768;
    wire N__72765;
    wire N__72762;
    wire N__72759;
    wire N__72754;
    wire N__72751;
    wire N__72748;
    wire N__72745;
    wire N__72740;
    wire N__72737;
    wire N__72734;
    wire N__72729;
    wire N__72722;
    wire N__72717;
    wire N__72712;
    wire N__72705;
    wire N__72702;
    wire N__72693;
    wire N__72690;
    wire N__72689;
    wire N__72686;
    wire N__72683;
    wire N__72682;
    wire N__72681;
    wire N__72678;
    wire N__72675;
    wire N__72672;
    wire N__72669;
    wire N__72666;
    wire N__72663;
    wire N__72660;
    wire N__72657;
    wire N__72654;
    wire N__72651;
    wire N__72642;
    wire N__72639;
    wire N__72638;
    wire N__72635;
    wire N__72632;
    wire N__72631;
    wire N__72626;
    wire N__72623;
    wire N__72620;
    wire N__72617;
    wire N__72612;
    wire N__72609;
    wire N__72606;
    wire N__72603;
    wire N__72600;
    wire N__72597;
    wire N__72594;
    wire N__72591;
    wire N__72588;
    wire N__72587;
    wire N__72586;
    wire N__72585;
    wire N__72582;
    wire N__72581;
    wire N__72578;
    wire N__72577;
    wire N__72574;
    wire N__72571;
    wire N__72570;
    wire N__72567;
    wire N__72564;
    wire N__72563;
    wire N__72560;
    wire N__72559;
    wire N__72556;
    wire N__72553;
    wire N__72550;
    wire N__72547;
    wire N__72542;
    wire N__72539;
    wire N__72536;
    wire N__72533;
    wire N__72530;
    wire N__72529;
    wire N__72528;
    wire N__72521;
    wire N__72518;
    wire N__72515;
    wire N__72508;
    wire N__72503;
    wire N__72500;
    wire N__72489;
    wire N__72486;
    wire N__72483;
    wire N__72482;
    wire N__72479;
    wire N__72476;
    wire N__72473;
    wire N__72472;
    wire N__72469;
    wire N__72468;
    wire N__72465;
    wire N__72464;
    wire N__72463;
    wire N__72460;
    wire N__72457;
    wire N__72454;
    wire N__72451;
    wire N__72448;
    wire N__72445;
    wire N__72442;
    wire N__72439;
    wire N__72436;
    wire N__72433;
    wire N__72430;
    wire N__72417;
    wire N__72414;
    wire N__72413;
    wire N__72410;
    wire N__72407;
    wire N__72404;
    wire N__72401;
    wire N__72398;
    wire N__72397;
    wire N__72396;
    wire N__72393;
    wire N__72390;
    wire N__72387;
    wire N__72384;
    wire N__72377;
    wire N__72372;
    wire N__72371;
    wire N__72370;
    wire N__72367;
    wire N__72366;
    wire N__72361;
    wire N__72360;
    wire N__72357;
    wire N__72354;
    wire N__72351;
    wire N__72348;
    wire N__72347;
    wire N__72342;
    wire N__72337;
    wire N__72334;
    wire N__72329;
    wire N__72326;
    wire N__72321;
    wire N__72320;
    wire N__72319;
    wire N__72318;
    wire N__72315;
    wire N__72310;
    wire N__72309;
    wire N__72306;
    wire N__72303;
    wire N__72300;
    wire N__72299;
    wire N__72296;
    wire N__72293;
    wire N__72288;
    wire N__72285;
    wire N__72284;
    wire N__72283;
    wire N__72280;
    wire N__72277;
    wire N__72274;
    wire N__72271;
    wire N__72268;
    wire N__72265;
    wire N__72252;
    wire N__72251;
    wire N__72246;
    wire N__72243;
    wire N__72242;
    wire N__72239;
    wire N__72238;
    wire N__72237;
    wire N__72234;
    wire N__72231;
    wire N__72226;
    wire N__72219;
    wire N__72216;
    wire N__72215;
    wire N__72214;
    wire N__72211;
    wire N__72210;
    wire N__72207;
    wire N__72206;
    wire N__72203;
    wire N__72200;
    wire N__72197;
    wire N__72196;
    wire N__72195;
    wire N__72192;
    wire N__72187;
    wire N__72182;
    wire N__72179;
    wire N__72176;
    wire N__72165;
    wire N__72162;
    wire N__72161;
    wire N__72158;
    wire N__72155;
    wire N__72154;
    wire N__72153;
    wire N__72152;
    wire N__72149;
    wire N__72146;
    wire N__72143;
    wire N__72138;
    wire N__72135;
    wire N__72130;
    wire N__72123;
    wire N__72120;
    wire N__72117;
    wire N__72114;
    wire N__72111;
    wire N__72110;
    wire N__72107;
    wire N__72104;
    wire N__72103;
    wire N__72100;
    wire N__72095;
    wire N__72090;
    wire N__72089;
    wire N__72088;
    wire N__72085;
    wire N__72082;
    wire N__72079;
    wire N__72078;
    wire N__72075;
    wire N__72072;
    wire N__72067;
    wire N__72060;
    wire N__72057;
    wire N__72054;
    wire N__72051;
    wire N__72050;
    wire N__72049;
    wire N__72046;
    wire N__72041;
    wire N__72036;
    wire N__72033;
    wire N__72032;
    wire N__72029;
    wire N__72026;
    wire N__72021;
    wire N__72018;
    wire N__72017;
    wire N__72014;
    wire N__72011;
    wire N__72006;
    wire N__72003;
    wire N__72002;
    wire N__72001;
    wire N__71998;
    wire N__71995;
    wire N__71992;
    wire N__71989;
    wire N__71988;
    wire N__71981;
    wire N__71978;
    wire N__71975;
    wire N__71970;
    wire N__71969;
    wire N__71968;
    wire N__71967;
    wire N__71966;
    wire N__71963;
    wire N__71960;
    wire N__71959;
    wire N__71958;
    wire N__71957;
    wire N__71954;
    wire N__71953;
    wire N__71950;
    wire N__71947;
    wire N__71946;
    wire N__71945;
    wire N__71944;
    wire N__71943;
    wire N__71940;
    wire N__71939;
    wire N__71938;
    wire N__71937;
    wire N__71936;
    wire N__71931;
    wire N__71928;
    wire N__71925;
    wire N__71922;
    wire N__71921;
    wire N__71918;
    wire N__71917;
    wire N__71916;
    wire N__71915;
    wire N__71914;
    wire N__71913;
    wire N__71910;
    wire N__71907;
    wire N__71906;
    wire N__71903;
    wire N__71902;
    wire N__71897;
    wire N__71894;
    wire N__71891;
    wire N__71888;
    wire N__71887;
    wire N__71884;
    wire N__71879;
    wire N__71876;
    wire N__71875;
    wire N__71872;
    wire N__71867;
    wire N__71866;
    wire N__71863;
    wire N__71860;
    wire N__71855;
    wire N__71850;
    wire N__71847;
    wire N__71842;
    wire N__71837;
    wire N__71834;
    wire N__71831;
    wire N__71828;
    wire N__71825;
    wire N__71822;
    wire N__71817;
    wire N__71816;
    wire N__71811;
    wire N__71808;
    wire N__71805;
    wire N__71802;
    wire N__71799;
    wire N__71796;
    wire N__71793;
    wire N__71790;
    wire N__71787;
    wire N__71782;
    wire N__71781;
    wire N__71778;
    wire N__71773;
    wire N__71768;
    wire N__71763;
    wire N__71762;
    wire N__71761;
    wire N__71758;
    wire N__71753;
    wire N__71744;
    wire N__71741;
    wire N__71734;
    wire N__71731;
    wire N__71726;
    wire N__71723;
    wire N__71720;
    wire N__71715;
    wire N__71712;
    wire N__71709;
    wire N__71706;
    wire N__71701;
    wire N__71692;
    wire N__71679;
    wire N__71676;
    wire N__71675;
    wire N__71674;
    wire N__71673;
    wire N__71670;
    wire N__71667;
    wire N__71662;
    wire N__71659;
    wire N__71656;
    wire N__71653;
    wire N__71646;
    wire N__71645;
    wire N__71642;
    wire N__71639;
    wire N__71636;
    wire N__71635;
    wire N__71632;
    wire N__71631;
    wire N__71628;
    wire N__71627;
    wire N__71624;
    wire N__71621;
    wire N__71618;
    wire N__71615;
    wire N__71612;
    wire N__71609;
    wire N__71606;
    wire N__71603;
    wire N__71598;
    wire N__71589;
    wire N__71588;
    wire N__71585;
    wire N__71582;
    wire N__71579;
    wire N__71576;
    wire N__71573;
    wire N__71572;
    wire N__71569;
    wire N__71566;
    wire N__71563;
    wire N__71560;
    wire N__71553;
    wire N__71552;
    wire N__71549;
    wire N__71546;
    wire N__71545;
    wire N__71544;
    wire N__71543;
    wire N__71542;
    wire N__71539;
    wire N__71538;
    wire N__71537;
    wire N__71536;
    wire N__71533;
    wire N__71530;
    wire N__71529;
    wire N__71526;
    wire N__71523;
    wire N__71520;
    wire N__71519;
    wire N__71516;
    wire N__71513;
    wire N__71510;
    wire N__71507;
    wire N__71506;
    wire N__71505;
    wire N__71504;
    wire N__71499;
    wire N__71496;
    wire N__71493;
    wire N__71490;
    wire N__71487;
    wire N__71484;
    wire N__71483;
    wire N__71482;
    wire N__71477;
    wire N__71474;
    wire N__71473;
    wire N__71472;
    wire N__71471;
    wire N__71468;
    wire N__71465;
    wire N__71462;
    wire N__71459;
    wire N__71458;
    wire N__71457;
    wire N__71456;
    wire N__71455;
    wire N__71454;
    wire N__71451;
    wire N__71448;
    wire N__71445;
    wire N__71442;
    wire N__71437;
    wire N__71432;
    wire N__71429;
    wire N__71428;
    wire N__71425;
    wire N__71418;
    wire N__71409;
    wire N__71406;
    wire N__71403;
    wire N__71398;
    wire N__71395;
    wire N__71394;
    wire N__71391;
    wire N__71388;
    wire N__71379;
    wire N__71376;
    wire N__71373;
    wire N__71372;
    wire N__71369;
    wire N__71366;
    wire N__71355;
    wire N__71352;
    wire N__71351;
    wire N__71350;
    wire N__71349;
    wire N__71348;
    wire N__71347;
    wire N__71344;
    wire N__71341;
    wire N__71338;
    wire N__71333;
    wire N__71330;
    wire N__71321;
    wire N__71310;
    wire N__71295;
    wire N__71292;
    wire N__71289;
    wire N__71286;
    wire N__71283;
    wire N__71280;
    wire N__71277;
    wire N__71274;
    wire N__71271;
    wire N__71270;
    wire N__71269;
    wire N__71268;
    wire N__71265;
    wire N__71260;
    wire N__71257;
    wire N__71254;
    wire N__71247;
    wire N__71246;
    wire N__71243;
    wire N__71242;
    wire N__71239;
    wire N__71236;
    wire N__71233;
    wire N__71230;
    wire N__71225;
    wire N__71220;
    wire N__71219;
    wire N__71216;
    wire N__71213;
    wire N__71210;
    wire N__71209;
    wire N__71206;
    wire N__71203;
    wire N__71200;
    wire N__71197;
    wire N__71192;
    wire N__71187;
    wire N__71184;
    wire N__71181;
    wire N__71178;
    wire N__71177;
    wire N__71176;
    wire N__71175;
    wire N__71172;
    wire N__71169;
    wire N__71166;
    wire N__71163;
    wire N__71158;
    wire N__71155;
    wire N__71148;
    wire N__71145;
    wire N__71142;
    wire N__71139;
    wire N__71136;
    wire N__71133;
    wire N__71130;
    wire N__71127;
    wire N__71126;
    wire N__71123;
    wire N__71120;
    wire N__71119;
    wire N__71118;
    wire N__71117;
    wire N__71116;
    wire N__71115;
    wire N__71114;
    wire N__71113;
    wire N__71110;
    wire N__71107;
    wire N__71104;
    wire N__71101;
    wire N__71100;
    wire N__71099;
    wire N__71096;
    wire N__71095;
    wire N__71094;
    wire N__71093;
    wire N__71092;
    wire N__71091;
    wire N__71088;
    wire N__71081;
    wire N__71080;
    wire N__71079;
    wire N__71078;
    wire N__71077;
    wire N__71068;
    wire N__71065;
    wire N__71062;
    wire N__71059;
    wire N__71054;
    wire N__71051;
    wire N__71046;
    wire N__71041;
    wire N__71036;
    wire N__71033;
    wire N__71032;
    wire N__71031;
    wire N__71030;
    wire N__71027;
    wire N__71024;
    wire N__71019;
    wire N__71016;
    wire N__71005;
    wire N__71002;
    wire N__70999;
    wire N__70994;
    wire N__70989;
    wire N__70982;
    wire N__70971;
    wire N__70968;
    wire N__70965;
    wire N__70962;
    wire N__70959;
    wire N__70958;
    wire N__70955;
    wire N__70952;
    wire N__70949;
    wire N__70946;
    wire N__70943;
    wire N__70940;
    wire N__70937;
    wire N__70932;
    wire N__70929;
    wire N__70926;
    wire N__70923;
    wire N__70922;
    wire N__70919;
    wire N__70916;
    wire N__70915;
    wire N__70910;
    wire N__70907;
    wire N__70902;
    wire N__70899;
    wire N__70896;
    wire N__70893;
    wire N__70890;
    wire N__70887;
    wire N__70886;
    wire N__70885;
    wire N__70880;
    wire N__70877;
    wire N__70876;
    wire N__70873;
    wire N__70870;
    wire N__70867;
    wire N__70864;
    wire N__70861;
    wire N__70854;
    wire N__70851;
    wire N__70850;
    wire N__70849;
    wire N__70848;
    wire N__70847;
    wire N__70844;
    wire N__70841;
    wire N__70838;
    wire N__70835;
    wire N__70832;
    wire N__70827;
    wire N__70818;
    wire N__70815;
    wire N__70812;
    wire N__70809;
    wire N__70808;
    wire N__70805;
    wire N__70802;
    wire N__70799;
    wire N__70796;
    wire N__70793;
    wire N__70788;
    wire N__70787;
    wire N__70784;
    wire N__70781;
    wire N__70778;
    wire N__70775;
    wire N__70774;
    wire N__70771;
    wire N__70768;
    wire N__70765;
    wire N__70760;
    wire N__70757;
    wire N__70754;
    wire N__70749;
    wire N__70746;
    wire N__70743;
    wire N__70742;
    wire N__70741;
    wire N__70738;
    wire N__70735;
    wire N__70732;
    wire N__70727;
    wire N__70724;
    wire N__70721;
    wire N__70716;
    wire N__70715;
    wire N__70712;
    wire N__70709;
    wire N__70706;
    wire N__70701;
    wire N__70698;
    wire N__70695;
    wire N__70694;
    wire N__70691;
    wire N__70688;
    wire N__70683;
    wire N__70680;
    wire N__70677;
    wire N__70674;
    wire N__70673;
    wire N__70672;
    wire N__70669;
    wire N__70666;
    wire N__70663;
    wire N__70660;
    wire N__70659;
    wire N__70658;
    wire N__70655;
    wire N__70652;
    wire N__70649;
    wire N__70646;
    wire N__70645;
    wire N__70642;
    wire N__70637;
    wire N__70632;
    wire N__70627;
    wire N__70620;
    wire N__70619;
    wire N__70618;
    wire N__70615;
    wire N__70612;
    wire N__70609;
    wire N__70602;
    wire N__70599;
    wire N__70598;
    wire N__70595;
    wire N__70592;
    wire N__70591;
    wire N__70588;
    wire N__70585;
    wire N__70582;
    wire N__70575;
    wire N__70572;
    wire N__70571;
    wire N__70568;
    wire N__70565;
    wire N__70562;
    wire N__70559;
    wire N__70556;
    wire N__70551;
    wire N__70550;
    wire N__70549;
    wire N__70548;
    wire N__70545;
    wire N__70542;
    wire N__70537;
    wire N__70534;
    wire N__70531;
    wire N__70528;
    wire N__70527;
    wire N__70524;
    wire N__70519;
    wire N__70516;
    wire N__70513;
    wire N__70506;
    wire N__70505;
    wire N__70502;
    wire N__70499;
    wire N__70498;
    wire N__70495;
    wire N__70492;
    wire N__70489;
    wire N__70482;
    wire N__70479;
    wire N__70476;
    wire N__70473;
    wire N__70470;
    wire N__70469;
    wire N__70466;
    wire N__70463;
    wire N__70458;
    wire N__70455;
    wire N__70452;
    wire N__70449;
    wire N__70446;
    wire N__70445;
    wire N__70444;
    wire N__70443;
    wire N__70440;
    wire N__70439;
    wire N__70432;
    wire N__70429;
    wire N__70426;
    wire N__70425;
    wire N__70422;
    wire N__70417;
    wire N__70414;
    wire N__70411;
    wire N__70408;
    wire N__70401;
    wire N__70400;
    wire N__70397;
    wire N__70394;
    wire N__70391;
    wire N__70388;
    wire N__70387;
    wire N__70384;
    wire N__70381;
    wire N__70378;
    wire N__70373;
    wire N__70368;
    wire N__70365;
    wire N__70362;
    wire N__70359;
    wire N__70356;
    wire N__70353;
    wire N__70352;
    wire N__70349;
    wire N__70348;
    wire N__70347;
    wire N__70344;
    wire N__70341;
    wire N__70338;
    wire N__70335;
    wire N__70332;
    wire N__70329;
    wire N__70328;
    wire N__70325;
    wire N__70322;
    wire N__70319;
    wire N__70316;
    wire N__70313;
    wire N__70310;
    wire N__70299;
    wire N__70298;
    wire N__70297;
    wire N__70294;
    wire N__70291;
    wire N__70288;
    wire N__70285;
    wire N__70284;
    wire N__70281;
    wire N__70278;
    wire N__70277;
    wire N__70274;
    wire N__70271;
    wire N__70268;
    wire N__70265;
    wire N__70264;
    wire N__70261;
    wire N__70258;
    wire N__70253;
    wire N__70250;
    wire N__70247;
    wire N__70244;
    wire N__70233;
    wire N__70230;
    wire N__70229;
    wire N__70226;
    wire N__70225;
    wire N__70222;
    wire N__70219;
    wire N__70216;
    wire N__70215;
    wire N__70212;
    wire N__70209;
    wire N__70206;
    wire N__70203;
    wire N__70194;
    wire N__70193;
    wire N__70188;
    wire N__70187;
    wire N__70186;
    wire N__70183;
    wire N__70180;
    wire N__70179;
    wire N__70178;
    wire N__70175;
    wire N__70174;
    wire N__70173;
    wire N__70172;
    wire N__70171;
    wire N__70170;
    wire N__70169;
    wire N__70168;
    wire N__70167;
    wire N__70166;
    wire N__70165;
    wire N__70164;
    wire N__70159;
    wire N__70156;
    wire N__70155;
    wire N__70154;
    wire N__70153;
    wire N__70152;
    wire N__70151;
    wire N__70150;
    wire N__70149;
    wire N__70148;
    wire N__70147;
    wire N__70146;
    wire N__70145;
    wire N__70144;
    wire N__70143;
    wire N__70142;
    wire N__70141;
    wire N__70140;
    wire N__70139;
    wire N__70138;
    wire N__70131;
    wire N__70128;
    wire N__70121;
    wire N__70116;
    wire N__70107;
    wire N__70102;
    wire N__70097;
    wire N__70094;
    wire N__70091;
    wire N__70088;
    wire N__70087;
    wire N__70084;
    wire N__70083;
    wire N__70082;
    wire N__70081;
    wire N__70080;
    wire N__70079;
    wire N__70078;
    wire N__70075;
    wire N__70070;
    wire N__70063;
    wire N__70058;
    wire N__70055;
    wire N__70048;
    wire N__70045;
    wire N__70038;
    wire N__70031;
    wire N__70024;
    wire N__70023;
    wire N__70022;
    wire N__70019;
    wire N__70018;
    wire N__70017;
    wire N__70016;
    wire N__70015;
    wire N__70014;
    wire N__70005;
    wire N__69998;
    wire N__69993;
    wire N__69988;
    wire N__69979;
    wire N__69974;
    wire N__69969;
    wire N__69966;
    wire N__69963;
    wire N__69954;
    wire N__69951;
    wire N__69946;
    wire N__69941;
    wire N__69938;
    wire N__69935;
    wire N__69928;
    wire N__69925;
    wire N__69920;
    wire N__69917;
    wire N__69912;
    wire N__69903;
    wire N__69902;
    wire N__69899;
    wire N__69898;
    wire N__69895;
    wire N__69894;
    wire N__69891;
    wire N__69888;
    wire N__69885;
    wire N__69884;
    wire N__69881;
    wire N__69878;
    wire N__69873;
    wire N__69870;
    wire N__69867;
    wire N__69862;
    wire N__69861;
    wire N__69860;
    wire N__69857;
    wire N__69852;
    wire N__69847;
    wire N__69844;
    wire N__69837;
    wire N__69834;
    wire N__69833;
    wire N__69832;
    wire N__69829;
    wire N__69826;
    wire N__69825;
    wire N__69822;
    wire N__69819;
    wire N__69814;
    wire N__69811;
    wire N__69804;
    wire N__69801;
    wire N__69800;
    wire N__69797;
    wire N__69794;
    wire N__69793;
    wire N__69792;
    wire N__69789;
    wire N__69788;
    wire N__69785;
    wire N__69780;
    wire N__69777;
    wire N__69774;
    wire N__69765;
    wire N__69762;
    wire N__69761;
    wire N__69760;
    wire N__69759;
    wire N__69758;
    wire N__69755;
    wire N__69752;
    wire N__69747;
    wire N__69744;
    wire N__69741;
    wire N__69738;
    wire N__69735;
    wire N__69732;
    wire N__69729;
    wire N__69728;
    wire N__69725;
    wire N__69720;
    wire N__69717;
    wire N__69714;
    wire N__69709;
    wire N__69702;
    wire N__69701;
    wire N__69700;
    wire N__69697;
    wire N__69694;
    wire N__69693;
    wire N__69690;
    wire N__69687;
    wire N__69684;
    wire N__69681;
    wire N__69672;
    wire N__69669;
    wire N__69666;
    wire N__69663;
    wire N__69660;
    wire N__69657;
    wire N__69654;
    wire N__69651;
    wire N__69648;
    wire N__69645;
    wire N__69644;
    wire N__69641;
    wire N__69640;
    wire N__69637;
    wire N__69634;
    wire N__69631;
    wire N__69630;
    wire N__69627;
    wire N__69624;
    wire N__69619;
    wire N__69616;
    wire N__69609;
    wire N__69608;
    wire N__69605;
    wire N__69602;
    wire N__69599;
    wire N__69596;
    wire N__69593;
    wire N__69590;
    wire N__69585;
    wire N__69584;
    wire N__69583;
    wire N__69582;
    wire N__69581;
    wire N__69580;
    wire N__69577;
    wire N__69574;
    wire N__69567;
    wire N__69564;
    wire N__69561;
    wire N__69558;
    wire N__69557;
    wire N__69554;
    wire N__69551;
    wire N__69550;
    wire N__69549;
    wire N__69548;
    wire N__69547;
    wire N__69546;
    wire N__69543;
    wire N__69540;
    wire N__69537;
    wire N__69532;
    wire N__69525;
    wire N__69522;
    wire N__69519;
    wire N__69504;
    wire N__69501;
    wire N__69500;
    wire N__69495;
    wire N__69492;
    wire N__69491;
    wire N__69488;
    wire N__69485;
    wire N__69482;
    wire N__69481;
    wire N__69480;
    wire N__69475;
    wire N__69472;
    wire N__69469;
    wire N__69462;
    wire N__69461;
    wire N__69460;
    wire N__69459;
    wire N__69454;
    wire N__69451;
    wire N__69450;
    wire N__69447;
    wire N__69444;
    wire N__69441;
    wire N__69438;
    wire N__69437;
    wire N__69434;
    wire N__69431;
    wire N__69426;
    wire N__69423;
    wire N__69420;
    wire N__69415;
    wire N__69412;
    wire N__69411;
    wire N__69410;
    wire N__69407;
    wire N__69402;
    wire N__69399;
    wire N__69396;
    wire N__69387;
    wire N__69384;
    wire N__69381;
    wire N__69380;
    wire N__69377;
    wire N__69376;
    wire N__69373;
    wire N__69370;
    wire N__69367;
    wire N__69364;
    wire N__69363;
    wire N__69362;
    wire N__69355;
    wire N__69354;
    wire N__69351;
    wire N__69348;
    wire N__69345;
    wire N__69342;
    wire N__69337;
    wire N__69330;
    wire N__69329;
    wire N__69326;
    wire N__69325;
    wire N__69322;
    wire N__69321;
    wire N__69320;
    wire N__69317;
    wire N__69314;
    wire N__69313;
    wire N__69310;
    wire N__69305;
    wire N__69302;
    wire N__69301;
    wire N__69298;
    wire N__69295;
    wire N__69288;
    wire N__69285;
    wire N__69276;
    wire N__69275;
    wire N__69272;
    wire N__69267;
    wire N__69264;
    wire N__69263;
    wire N__69262;
    wire N__69255;
    wire N__69252;
    wire N__69249;
    wire N__69246;
    wire N__69243;
    wire N__69240;
    wire N__69237;
    wire N__69236;
    wire N__69235;
    wire N__69228;
    wire N__69227;
    wire N__69226;
    wire N__69225;
    wire N__69224;
    wire N__69223;
    wire N__69220;
    wire N__69215;
    wire N__69212;
    wire N__69211;
    wire N__69210;
    wire N__69205;
    wire N__69204;
    wire N__69201;
    wire N__69200;
    wire N__69199;
    wire N__69196;
    wire N__69195;
    wire N__69194;
    wire N__69191;
    wire N__69186;
    wire N__69185;
    wire N__69184;
    wire N__69183;
    wire N__69182;
    wire N__69181;
    wire N__69180;
    wire N__69177;
    wire N__69174;
    wire N__69171;
    wire N__69170;
    wire N__69167;
    wire N__69166;
    wire N__69163;
    wire N__69162;
    wire N__69161;
    wire N__69158;
    wire N__69157;
    wire N__69156;
    wire N__69151;
    wire N__69150;
    wire N__69147;
    wire N__69144;
    wire N__69141;
    wire N__69136;
    wire N__69129;
    wire N__69124;
    wire N__69121;
    wire N__69118;
    wire N__69117;
    wire N__69112;
    wire N__69109;
    wire N__69104;
    wire N__69101;
    wire N__69098;
    wire N__69095;
    wire N__69092;
    wire N__69091;
    wire N__69088;
    wire N__69085;
    wire N__69078;
    wire N__69075;
    wire N__69072;
    wire N__69069;
    wire N__69068;
    wire N__69065;
    wire N__69062;
    wire N__69059;
    wire N__69050;
    wire N__69047;
    wire N__69044;
    wire N__69041;
    wire N__69038;
    wire N__69035;
    wire N__69032;
    wire N__69025;
    wire N__69022;
    wire N__69019;
    wire N__69012;
    wire N__69007;
    wire N__69000;
    wire N__68995;
    wire N__68982;
    wire N__68979;
    wire N__68976;
    wire N__68973;
    wire N__68970;
    wire N__68969;
    wire N__68966;
    wire N__68963;
    wire N__68960;
    wire N__68959;
    wire N__68958;
    wire N__68957;
    wire N__68954;
    wire N__68951;
    wire N__68948;
    wire N__68945;
    wire N__68942;
    wire N__68931;
    wire N__68928;
    wire N__68927;
    wire N__68924;
    wire N__68923;
    wire N__68920;
    wire N__68917;
    wire N__68914;
    wire N__68911;
    wire N__68908;
    wire N__68901;
    wire N__68900;
    wire N__68895;
    wire N__68892;
    wire N__68889;
    wire N__68886;
    wire N__68883;
    wire N__68880;
    wire N__68879;
    wire N__68876;
    wire N__68873;
    wire N__68870;
    wire N__68867;
    wire N__68864;
    wire N__68861;
    wire N__68858;
    wire N__68855;
    wire N__68850;
    wire N__68849;
    wire N__68848;
    wire N__68847;
    wire N__68846;
    wire N__68845;
    wire N__68844;
    wire N__68843;
    wire N__68842;
    wire N__68841;
    wire N__68840;
    wire N__68837;
    wire N__68832;
    wire N__68829;
    wire N__68826;
    wire N__68821;
    wire N__68814;
    wire N__68811;
    wire N__68796;
    wire N__68795;
    wire N__68794;
    wire N__68793;
    wire N__68790;
    wire N__68787;
    wire N__68782;
    wire N__68781;
    wire N__68780;
    wire N__68777;
    wire N__68774;
    wire N__68771;
    wire N__68766;
    wire N__68757;
    wire N__68756;
    wire N__68753;
    wire N__68752;
    wire N__68751;
    wire N__68750;
    wire N__68749;
    wire N__68746;
    wire N__68743;
    wire N__68740;
    wire N__68737;
    wire N__68734;
    wire N__68733;
    wire N__68732;
    wire N__68729;
    wire N__68728;
    wire N__68727;
    wire N__68726;
    wire N__68723;
    wire N__68716;
    wire N__68713;
    wire N__68710;
    wire N__68707;
    wire N__68702;
    wire N__68699;
    wire N__68696;
    wire N__68679;
    wire N__68678;
    wire N__68677;
    wire N__68672;
    wire N__68671;
    wire N__68670;
    wire N__68669;
    wire N__68666;
    wire N__68663;
    wire N__68660;
    wire N__68655;
    wire N__68646;
    wire N__68645;
    wire N__68642;
    wire N__68639;
    wire N__68634;
    wire N__68633;
    wire N__68628;
    wire N__68625;
    wire N__68624;
    wire N__68623;
    wire N__68622;
    wire N__68619;
    wire N__68612;
    wire N__68607;
    wire N__68604;
    wire N__68601;
    wire N__68600;
    wire N__68597;
    wire N__68594;
    wire N__68593;
    wire N__68588;
    wire N__68585;
    wire N__68582;
    wire N__68579;
    wire N__68576;
    wire N__68571;
    wire N__68570;
    wire N__68567;
    wire N__68564;
    wire N__68559;
    wire N__68556;
    wire N__68555;
    wire N__68552;
    wire N__68549;
    wire N__68546;
    wire N__68545;
    wire N__68544;
    wire N__68543;
    wire N__68542;
    wire N__68539;
    wire N__68536;
    wire N__68533;
    wire N__68532;
    wire N__68531;
    wire N__68528;
    wire N__68527;
    wire N__68524;
    wire N__68521;
    wire N__68518;
    wire N__68513;
    wire N__68512;
    wire N__68511;
    wire N__68510;
    wire N__68507;
    wire N__68504;
    wire N__68501;
    wire N__68498;
    wire N__68497;
    wire N__68496;
    wire N__68495;
    wire N__68490;
    wire N__68485;
    wire N__68482;
    wire N__68477;
    wire N__68472;
    wire N__68467;
    wire N__68464;
    wire N__68459;
    wire N__68442;
    wire N__68441;
    wire N__68438;
    wire N__68437;
    wire N__68434;
    wire N__68433;
    wire N__68432;
    wire N__68429;
    wire N__68426;
    wire N__68423;
    wire N__68422;
    wire N__68419;
    wire N__68416;
    wire N__68411;
    wire N__68408;
    wire N__68405;
    wire N__68402;
    wire N__68399;
    wire N__68396;
    wire N__68395;
    wire N__68390;
    wire N__68387;
    wire N__68382;
    wire N__68379;
    wire N__68370;
    wire N__68367;
    wire N__68366;
    wire N__68365;
    wire N__68362;
    wire N__68359;
    wire N__68356;
    wire N__68353;
    wire N__68350;
    wire N__68349;
    wire N__68346;
    wire N__68343;
    wire N__68340;
    wire N__68337;
    wire N__68334;
    wire N__68331;
    wire N__68328;
    wire N__68319;
    wire N__68316;
    wire N__68313;
    wire N__68312;
    wire N__68311;
    wire N__68308;
    wire N__68305;
    wire N__68302;
    wire N__68295;
    wire N__68292;
    wire N__68289;
    wire N__68286;
    wire N__68283;
    wire N__68280;
    wire N__68279;
    wire N__68278;
    wire N__68275;
    wire N__68270;
    wire N__68267;
    wire N__68262;
    wire N__68261;
    wire N__68258;
    wire N__68255;
    wire N__68252;
    wire N__68247;
    wire N__68244;
    wire N__68241;
    wire N__68240;
    wire N__68237;
    wire N__68232;
    wire N__68229;
    wire N__68228;
    wire N__68223;
    wire N__68220;
    wire N__68217;
    wire N__68216;
    wire N__68215;
    wire N__68212;
    wire N__68209;
    wire N__68206;
    wire N__68203;
    wire N__68200;
    wire N__68197;
    wire N__68190;
    wire N__68189;
    wire N__68186;
    wire N__68183;
    wire N__68180;
    wire N__68177;
    wire N__68174;
    wire N__68171;
    wire N__68168;
    wire N__68163;
    wire N__68162;
    wire N__68161;
    wire N__68160;
    wire N__68157;
    wire N__68150;
    wire N__68145;
    wire N__68142;
    wire N__68141;
    wire N__68140;
    wire N__68137;
    wire N__68132;
    wire N__68127;
    wire N__68126;
    wire N__68123;
    wire N__68122;
    wire N__68121;
    wire N__68120;
    wire N__68117;
    wire N__68114;
    wire N__68111;
    wire N__68110;
    wire N__68109;
    wire N__68108;
    wire N__68105;
    wire N__68102;
    wire N__68097;
    wire N__68096;
    wire N__68095;
    wire N__68094;
    wire N__68093;
    wire N__68090;
    wire N__68083;
    wire N__68082;
    wire N__68081;
    wire N__68078;
    wire N__68073;
    wire N__68068;
    wire N__68063;
    wire N__68058;
    wire N__68053;
    wire N__68040;
    wire N__68039;
    wire N__68038;
    wire N__68035;
    wire N__68034;
    wire N__68031;
    wire N__68030;
    wire N__68029;
    wire N__68028;
    wire N__68025;
    wire N__68022;
    wire N__68019;
    wire N__68014;
    wire N__68009;
    wire N__67998;
    wire N__67995;
    wire N__67992;
    wire N__67989;
    wire N__67986;
    wire N__67985;
    wire N__67984;
    wire N__67981;
    wire N__67978;
    wire N__67975;
    wire N__67972;
    wire N__67969;
    wire N__67968;
    wire N__67967;
    wire N__67964;
    wire N__67959;
    wire N__67956;
    wire N__67953;
    wire N__67944;
    wire N__67943;
    wire N__67942;
    wire N__67941;
    wire N__67938;
    wire N__67935;
    wire N__67934;
    wire N__67931;
    wire N__67928;
    wire N__67925;
    wire N__67922;
    wire N__67919;
    wire N__67916;
    wire N__67915;
    wire N__67914;
    wire N__67911;
    wire N__67908;
    wire N__67903;
    wire N__67900;
    wire N__67895;
    wire N__67884;
    wire N__67883;
    wire N__67880;
    wire N__67877;
    wire N__67874;
    wire N__67873;
    wire N__67870;
    wire N__67867;
    wire N__67864;
    wire N__67863;
    wire N__67862;
    wire N__67859;
    wire N__67856;
    wire N__67853;
    wire N__67850;
    wire N__67847;
    wire N__67844;
    wire N__67841;
    wire N__67838;
    wire N__67835;
    wire N__67824;
    wire N__67821;
    wire N__67820;
    wire N__67819;
    wire N__67816;
    wire N__67813;
    wire N__67810;
    wire N__67805;
    wire N__67802;
    wire N__67797;
    wire N__67794;
    wire N__67793;
    wire N__67792;
    wire N__67789;
    wire N__67786;
    wire N__67783;
    wire N__67780;
    wire N__67773;
    wire N__67770;
    wire N__67767;
    wire N__67764;
    wire N__67761;
    wire N__67758;
    wire N__67755;
    wire N__67752;
    wire N__67749;
    wire N__67748;
    wire N__67745;
    wire N__67742;
    wire N__67739;
    wire N__67736;
    wire N__67733;
    wire N__67730;
    wire N__67725;
    wire N__67722;
    wire N__67719;
    wire N__67716;
    wire N__67713;
    wire N__67710;
    wire N__67707;
    wire N__67706;
    wire N__67703;
    wire N__67700;
    wire N__67695;
    wire N__67692;
    wire N__67689;
    wire N__67686;
    wire N__67683;
    wire N__67680;
    wire N__67677;
    wire N__67674;
    wire N__67671;
    wire N__67668;
    wire N__67665;
    wire N__67664;
    wire N__67661;
    wire N__67658;
    wire N__67657;
    wire N__67652;
    wire N__67649;
    wire N__67648;
    wire N__67645;
    wire N__67644;
    wire N__67641;
    wire N__67640;
    wire N__67637;
    wire N__67634;
    wire N__67631;
    wire N__67628;
    wire N__67625;
    wire N__67622;
    wire N__67621;
    wire N__67620;
    wire N__67617;
    wire N__67614;
    wire N__67607;
    wire N__67602;
    wire N__67593;
    wire N__67592;
    wire N__67591;
    wire N__67588;
    wire N__67585;
    wire N__67582;
    wire N__67577;
    wire N__67574;
    wire N__67571;
    wire N__67566;
    wire N__67563;
    wire N__67560;
    wire N__67559;
    wire N__67556;
    wire N__67553;
    wire N__67552;
    wire N__67551;
    wire N__67550;
    wire N__67549;
    wire N__67544;
    wire N__67539;
    wire N__67536;
    wire N__67533;
    wire N__67532;
    wire N__67529;
    wire N__67522;
    wire N__67519;
    wire N__67516;
    wire N__67513;
    wire N__67506;
    wire N__67505;
    wire N__67502;
    wire N__67501;
    wire N__67500;
    wire N__67499;
    wire N__67496;
    wire N__67493;
    wire N__67492;
    wire N__67491;
    wire N__67488;
    wire N__67483;
    wire N__67480;
    wire N__67477;
    wire N__67472;
    wire N__67461;
    wire N__67458;
    wire N__67455;
    wire N__67452;
    wire N__67449;
    wire N__67446;
    wire N__67443;
    wire N__67440;
    wire N__67437;
    wire N__67434;
    wire N__67431;
    wire N__67428;
    wire N__67425;
    wire N__67422;
    wire N__67419;
    wire N__67416;
    wire N__67415;
    wire N__67412;
    wire N__67409;
    wire N__67406;
    wire N__67403;
    wire N__67398;
    wire N__67395;
    wire N__67392;
    wire N__67389;
    wire N__67386;
    wire N__67383;
    wire N__67380;
    wire N__67377;
    wire N__67376;
    wire N__67373;
    wire N__67370;
    wire N__67365;
    wire N__67362;
    wire N__67361;
    wire N__67358;
    wire N__67355;
    wire N__67352;
    wire N__67351;
    wire N__67348;
    wire N__67345;
    wire N__67342;
    wire N__67335;
    wire N__67332;
    wire N__67329;
    wire N__67328;
    wire N__67327;
    wire N__67324;
    wire N__67321;
    wire N__67318;
    wire N__67315;
    wire N__67314;
    wire N__67313;
    wire N__67310;
    wire N__67307;
    wire N__67304;
    wire N__67301;
    wire N__67298;
    wire N__67297;
    wire N__67296;
    wire N__67287;
    wire N__67284;
    wire N__67281;
    wire N__67278;
    wire N__67275;
    wire N__67272;
    wire N__67269;
    wire N__67260;
    wire N__67257;
    wire N__67256;
    wire N__67255;
    wire N__67252;
    wire N__67251;
    wire N__67250;
    wire N__67249;
    wire N__67248;
    wire N__67243;
    wire N__67240;
    wire N__67235;
    wire N__67230;
    wire N__67223;
    wire N__67218;
    wire N__67215;
    wire N__67214;
    wire N__67213;
    wire N__67212;
    wire N__67209;
    wire N__67204;
    wire N__67201;
    wire N__67194;
    wire N__67193;
    wire N__67190;
    wire N__67187;
    wire N__67184;
    wire N__67181;
    wire N__67180;
    wire N__67177;
    wire N__67174;
    wire N__67171;
    wire N__67164;
    wire N__67163;
    wire N__67160;
    wire N__67157;
    wire N__67152;
    wire N__67151;
    wire N__67150;
    wire N__67149;
    wire N__67148;
    wire N__67147;
    wire N__67144;
    wire N__67141;
    wire N__67140;
    wire N__67137;
    wire N__67128;
    wire N__67125;
    wire N__67122;
    wire N__67121;
    wire N__67118;
    wire N__67115;
    wire N__67112;
    wire N__67109;
    wire N__67106;
    wire N__67099;
    wire N__67096;
    wire N__67089;
    wire N__67086;
    wire N__67083;
    wire N__67082;
    wire N__67079;
    wire N__67076;
    wire N__67071;
    wire N__67070;
    wire N__67067;
    wire N__67064;
    wire N__67061;
    wire N__67056;
    wire N__67055;
    wire N__67052;
    wire N__67049;
    wire N__67046;
    wire N__67043;
    wire N__67038;
    wire N__67037;
    wire N__67034;
    wire N__67033;
    wire N__67030;
    wire N__67027;
    wire N__67024;
    wire N__67021;
    wire N__67018;
    wire N__67015;
    wire N__67012;
    wire N__67005;
    wire N__67002;
    wire N__66999;
    wire N__66998;
    wire N__66995;
    wire N__66992;
    wire N__66987;
    wire N__66986;
    wire N__66985;
    wire N__66984;
    wire N__66979;
    wire N__66976;
    wire N__66973;
    wire N__66970;
    wire N__66965;
    wire N__66962;
    wire N__66957;
    wire N__66954;
    wire N__66951;
    wire N__66950;
    wire N__66947;
    wire N__66944;
    wire N__66939;
    wire N__66936;
    wire N__66933;
    wire N__66930;
    wire N__66929;
    wire N__66926;
    wire N__66923;
    wire N__66920;
    wire N__66919;
    wire N__66916;
    wire N__66913;
    wire N__66910;
    wire N__66903;
    wire N__66900;
    wire N__66899;
    wire N__66898;
    wire N__66897;
    wire N__66894;
    wire N__66893;
    wire N__66890;
    wire N__66887;
    wire N__66884;
    wire N__66881;
    wire N__66878;
    wire N__66875;
    wire N__66872;
    wire N__66871;
    wire N__66864;
    wire N__66863;
    wire N__66858;
    wire N__66855;
    wire N__66852;
    wire N__66849;
    wire N__66846;
    wire N__66841;
    wire N__66838;
    wire N__66831;
    wire N__66828;
    wire N__66827;
    wire N__66824;
    wire N__66821;
    wire N__66818;
    wire N__66813;
    wire N__66812;
    wire N__66811;
    wire N__66808;
    wire N__66807;
    wire N__66802;
    wire N__66799;
    wire N__66796;
    wire N__66793;
    wire N__66790;
    wire N__66787;
    wire N__66784;
    wire N__66781;
    wire N__66776;
    wire N__66771;
    wire N__66768;
    wire N__66765;
    wire N__66762;
    wire N__66759;
    wire N__66756;
    wire N__66753;
    wire N__66752;
    wire N__66751;
    wire N__66750;
    wire N__66747;
    wire N__66746;
    wire N__66743;
    wire N__66740;
    wire N__66737;
    wire N__66734;
    wire N__66731;
    wire N__66724;
    wire N__66721;
    wire N__66714;
    wire N__66711;
    wire N__66710;
    wire N__66709;
    wire N__66706;
    wire N__66703;
    wire N__66700;
    wire N__66697;
    wire N__66694;
    wire N__66687;
    wire N__66684;
    wire N__66681;
    wire N__66678;
    wire N__66675;
    wire N__66672;
    wire N__66669;
    wire N__66666;
    wire N__66663;
    wire N__66662;
    wire N__66661;
    wire N__66658;
    wire N__66655;
    wire N__66654;
    wire N__66651;
    wire N__66650;
    wire N__66647;
    wire N__66644;
    wire N__66641;
    wire N__66638;
    wire N__66637;
    wire N__66634;
    wire N__66629;
    wire N__66624;
    wire N__66621;
    wire N__66612;
    wire N__66609;
    wire N__66608;
    wire N__66605;
    wire N__66602;
    wire N__66597;
    wire N__66594;
    wire N__66593;
    wire N__66590;
    wire N__66587;
    wire N__66584;
    wire N__66579;
    wire N__66576;
    wire N__66573;
    wire N__66570;
    wire N__66569;
    wire N__66566;
    wire N__66565;
    wire N__66562;
    wire N__66559;
    wire N__66556;
    wire N__66553;
    wire N__66552;
    wire N__66549;
    wire N__66546;
    wire N__66543;
    wire N__66540;
    wire N__66537;
    wire N__66532;
    wire N__66525;
    wire N__66522;
    wire N__66521;
    wire N__66518;
    wire N__66517;
    wire N__66514;
    wire N__66511;
    wire N__66506;
    wire N__66501;
    wire N__66500;
    wire N__66497;
    wire N__66496;
    wire N__66495;
    wire N__66492;
    wire N__66487;
    wire N__66484;
    wire N__66481;
    wire N__66478;
    wire N__66475;
    wire N__66470;
    wire N__66465;
    wire N__66464;
    wire N__66461;
    wire N__66458;
    wire N__66455;
    wire N__66452;
    wire N__66447;
    wire N__66444;
    wire N__66441;
    wire N__66438;
    wire N__66435;
    wire N__66432;
    wire N__66431;
    wire N__66430;
    wire N__66427;
    wire N__66426;
    wire N__66425;
    wire N__66422;
    wire N__66419;
    wire N__66416;
    wire N__66411;
    wire N__66408;
    wire N__66403;
    wire N__66396;
    wire N__66393;
    wire N__66392;
    wire N__66389;
    wire N__66386;
    wire N__66381;
    wire N__66378;
    wire N__66375;
    wire N__66372;
    wire N__66369;
    wire N__66366;
    wire N__66365;
    wire N__66364;
    wire N__66361;
    wire N__66356;
    wire N__66355;
    wire N__66352;
    wire N__66349;
    wire N__66346;
    wire N__66339;
    wire N__66336;
    wire N__66335;
    wire N__66334;
    wire N__66333;
    wire N__66330;
    wire N__66327;
    wire N__66322;
    wire N__66315;
    wire N__66312;
    wire N__66309;
    wire N__66306;
    wire N__66303;
    wire N__66302;
    wire N__66299;
    wire N__66296;
    wire N__66293;
    wire N__66288;
    wire N__66285;
    wire N__66282;
    wire N__66279;
    wire N__66276;
    wire N__66273;
    wire N__66272;
    wire N__66271;
    wire N__66268;
    wire N__66265;
    wire N__66262;
    wire N__66259;
    wire N__66256;
    wire N__66253;
    wire N__66246;
    wire N__66243;
    wire N__66242;
    wire N__66239;
    wire N__66236;
    wire N__66233;
    wire N__66228;
    wire N__66227;
    wire N__66224;
    wire N__66221;
    wire N__66220;
    wire N__66217;
    wire N__66214;
    wire N__66211;
    wire N__66208;
    wire N__66205;
    wire N__66202;
    wire N__66199;
    wire N__66196;
    wire N__66189;
    wire N__66186;
    wire N__66183;
    wire N__66180;
    wire N__66177;
    wire N__66174;
    wire N__66173;
    wire N__66170;
    wire N__66167;
    wire N__66162;
    wire N__66161;
    wire N__66160;
    wire N__66157;
    wire N__66154;
    wire N__66151;
    wire N__66146;
    wire N__66143;
    wire N__66138;
    wire N__66135;
    wire N__66134;
    wire N__66133;
    wire N__66130;
    wire N__66125;
    wire N__66122;
    wire N__66117;
    wire N__66116;
    wire N__66113;
    wire N__66110;
    wire N__66107;
    wire N__66102;
    wire N__66099;
    wire N__66098;
    wire N__66097;
    wire N__66096;
    wire N__66093;
    wire N__66090;
    wire N__66087;
    wire N__66084;
    wire N__66081;
    wire N__66078;
    wire N__66073;
    wire N__66070;
    wire N__66063;
    wire N__66060;
    wire N__66057;
    wire N__66054;
    wire N__66053;
    wire N__66052;
    wire N__66049;
    wire N__66044;
    wire N__66041;
    wire N__66038;
    wire N__66033;
    wire N__66032;
    wire N__66027;
    wire N__66024;
    wire N__66021;
    wire N__66018;
    wire N__66017;
    wire N__66016;
    wire N__66011;
    wire N__66010;
    wire N__66007;
    wire N__66006;
    wire N__66003;
    wire N__66000;
    wire N__65995;
    wire N__65988;
    wire N__65987;
    wire N__65984;
    wire N__65981;
    wire N__65980;
    wire N__65977;
    wire N__65972;
    wire N__65969;
    wire N__65964;
    wire N__65961;
    wire N__65960;
    wire N__65959;
    wire N__65956;
    wire N__65953;
    wire N__65950;
    wire N__65947;
    wire N__65944;
    wire N__65941;
    wire N__65938;
    wire N__65931;
    wire N__65928;
    wire N__65927;
    wire N__65924;
    wire N__65921;
    wire N__65918;
    wire N__65915;
    wire N__65910;
    wire N__65907;
    wire N__65904;
    wire N__65903;
    wire N__65902;
    wire N__65899;
    wire N__65896;
    wire N__65893;
    wire N__65888;
    wire N__65885;
    wire N__65884;
    wire N__65881;
    wire N__65878;
    wire N__65875;
    wire N__65872;
    wire N__65869;
    wire N__65862;
    wire N__65861;
    wire N__65858;
    wire N__65855;
    wire N__65854;
    wire N__65853;
    wire N__65850;
    wire N__65847;
    wire N__65846;
    wire N__65841;
    wire N__65836;
    wire N__65835;
    wire N__65832;
    wire N__65829;
    wire N__65826;
    wire N__65823;
    wire N__65814;
    wire N__65811;
    wire N__65808;
    wire N__65805;
    wire N__65802;
    wire N__65799;
    wire N__65798;
    wire N__65795;
    wire N__65792;
    wire N__65787;
    wire N__65786;
    wire N__65783;
    wire N__65780;
    wire N__65779;
    wire N__65776;
    wire N__65773;
    wire N__65772;
    wire N__65769;
    wire N__65766;
    wire N__65763;
    wire N__65760;
    wire N__65757;
    wire N__65748;
    wire N__65747;
    wire N__65744;
    wire N__65741;
    wire N__65738;
    wire N__65735;
    wire N__65732;
    wire N__65729;
    wire N__65726;
    wire N__65721;
    wire N__65718;
    wire N__65717;
    wire N__65714;
    wire N__65711;
    wire N__65706;
    wire N__65705;
    wire N__65704;
    wire N__65703;
    wire N__65698;
    wire N__65697;
    wire N__65696;
    wire N__65691;
    wire N__65688;
    wire N__65685;
    wire N__65682;
    wire N__65679;
    wire N__65678;
    wire N__65675;
    wire N__65670;
    wire N__65667;
    wire N__65664;
    wire N__65655;
    wire N__65654;
    wire N__65651;
    wire N__65646;
    wire N__65643;
    wire N__65640;
    wire N__65639;
    wire N__65638;
    wire N__65637;
    wire N__65634;
    wire N__65633;
    wire N__65632;
    wire N__65631;
    wire N__65630;
    wire N__65627;
    wire N__65624;
    wire N__65621;
    wire N__65618;
    wire N__65613;
    wire N__65608;
    wire N__65595;
    wire N__65592;
    wire N__65591;
    wire N__65588;
    wire N__65585;
    wire N__65580;
    wire N__65577;
    wire N__65576;
    wire N__65573;
    wire N__65570;
    wire N__65567;
    wire N__65564;
    wire N__65561;
    wire N__65558;
    wire N__65553;
    wire N__65550;
    wire N__65549;
    wire N__65546;
    wire N__65543;
    wire N__65538;
    wire N__65535;
    wire N__65532;
    wire N__65529;
    wire N__65526;
    wire N__65525;
    wire N__65522;
    wire N__65519;
    wire N__65516;
    wire N__65511;
    wire N__65510;
    wire N__65507;
    wire N__65504;
    wire N__65501;
    wire N__65498;
    wire N__65493;
    wire N__65492;
    wire N__65489;
    wire N__65486;
    wire N__65481;
    wire N__65478;
    wire N__65475;
    wire N__65472;
    wire N__65469;
    wire N__65466;
    wire N__65463;
    wire N__65460;
    wire N__65457;
    wire N__65454;
    wire N__65453;
    wire N__65450;
    wire N__65447;
    wire N__65444;
    wire N__65441;
    wire N__65436;
    wire N__65435;
    wire N__65430;
    wire N__65427;
    wire N__65426;
    wire N__65423;
    wire N__65420;
    wire N__65419;
    wire N__65416;
    wire N__65413;
    wire N__65410;
    wire N__65407;
    wire N__65406;
    wire N__65405;
    wire N__65398;
    wire N__65395;
    wire N__65392;
    wire N__65385;
    wire N__65382;
    wire N__65379;
    wire N__65376;
    wire N__65373;
    wire N__65370;
    wire N__65369;
    wire N__65368;
    wire N__65365;
    wire N__65362;
    wire N__65359;
    wire N__65356;
    wire N__65353;
    wire N__65350;
    wire N__65347;
    wire N__65344;
    wire N__65337;
    wire N__65336;
    wire N__65335;
    wire N__65332;
    wire N__65331;
    wire N__65328;
    wire N__65327;
    wire N__65324;
    wire N__65319;
    wire N__65316;
    wire N__65313;
    wire N__65304;
    wire N__65301;
    wire N__65298;
    wire N__65297;
    wire N__65296;
    wire N__65295;
    wire N__65292;
    wire N__65287;
    wire N__65286;
    wire N__65283;
    wire N__65278;
    wire N__65275;
    wire N__65272;
    wire N__65269;
    wire N__65266;
    wire N__65263;
    wire N__65260;
    wire N__65253;
    wire N__65250;
    wire N__65247;
    wire N__65244;
    wire N__65241;
    wire N__65238;
    wire N__65235;
    wire N__65232;
    wire N__65229;
    wire N__65226;
    wire N__65223;
    wire N__65222;
    wire N__65221;
    wire N__65220;
    wire N__65217;
    wire N__65214;
    wire N__65209;
    wire N__65202;
    wire N__65201;
    wire N__65200;
    wire N__65197;
    wire N__65194;
    wire N__65193;
    wire N__65190;
    wire N__65185;
    wire N__65184;
    wire N__65181;
    wire N__65178;
    wire N__65175;
    wire N__65172;
    wire N__65163;
    wire N__65160;
    wire N__65157;
    wire N__65154;
    wire N__65151;
    wire N__65150;
    wire N__65147;
    wire N__65144;
    wire N__65143;
    wire N__65140;
    wire N__65137;
    wire N__65134;
    wire N__65127;
    wire N__65126;
    wire N__65121;
    wire N__65118;
    wire N__65115;
    wire N__65112;
    wire N__65111;
    wire N__65110;
    wire N__65109;
    wire N__65108;
    wire N__65105;
    wire N__65102;
    wire N__65097;
    wire N__65096;
    wire N__65093;
    wire N__65088;
    wire N__65085;
    wire N__65082;
    wire N__65079;
    wire N__65074;
    wire N__65073;
    wire N__65070;
    wire N__65069;
    wire N__65068;
    wire N__65065;
    wire N__65062;
    wire N__65059;
    wire N__65056;
    wire N__65051;
    wire N__65040;
    wire N__65039;
    wire N__65036;
    wire N__65035;
    wire N__65032;
    wire N__65029;
    wire N__65026;
    wire N__65023;
    wire N__65020;
    wire N__65017;
    wire N__65010;
    wire N__65009;
    wire N__65006;
    wire N__65003;
    wire N__65000;
    wire N__64997;
    wire N__64994;
    wire N__64989;
    wire N__64988;
    wire N__64987;
    wire N__64986;
    wire N__64983;
    wire N__64980;
    wire N__64977;
    wire N__64974;
    wire N__64971;
    wire N__64968;
    wire N__64967;
    wire N__64966;
    wire N__64965;
    wire N__64962;
    wire N__64959;
    wire N__64956;
    wire N__64953;
    wire N__64950;
    wire N__64947;
    wire N__64944;
    wire N__64939;
    wire N__64936;
    wire N__64931;
    wire N__64928;
    wire N__64923;
    wire N__64914;
    wire N__64911;
    wire N__64908;
    wire N__64905;
    wire N__64902;
    wire N__64901;
    wire N__64898;
    wire N__64897;
    wire N__64894;
    wire N__64891;
    wire N__64888;
    wire N__64885;
    wire N__64884;
    wire N__64883;
    wire N__64880;
    wire N__64877;
    wire N__64874;
    wire N__64873;
    wire N__64868;
    wire N__64863;
    wire N__64860;
    wire N__64857;
    wire N__64854;
    wire N__64851;
    wire N__64848;
    wire N__64839;
    wire N__64838;
    wire N__64835;
    wire N__64834;
    wire N__64831;
    wire N__64828;
    wire N__64827;
    wire N__64824;
    wire N__64821;
    wire N__64820;
    wire N__64819;
    wire N__64818;
    wire N__64817;
    wire N__64814;
    wire N__64811;
    wire N__64808;
    wire N__64805;
    wire N__64796;
    wire N__64793;
    wire N__64788;
    wire N__64779;
    wire N__64778;
    wire N__64777;
    wire N__64774;
    wire N__64773;
    wire N__64772;
    wire N__64769;
    wire N__64768;
    wire N__64765;
    wire N__64764;
    wire N__64761;
    wire N__64756;
    wire N__64755;
    wire N__64752;
    wire N__64749;
    wire N__64746;
    wire N__64743;
    wire N__64738;
    wire N__64737;
    wire N__64734;
    wire N__64733;
    wire N__64728;
    wire N__64725;
    wire N__64724;
    wire N__64719;
    wire N__64716;
    wire N__64713;
    wire N__64710;
    wire N__64705;
    wire N__64702;
    wire N__64697;
    wire N__64686;
    wire N__64683;
    wire N__64680;
    wire N__64677;
    wire N__64674;
    wire N__64673;
    wire N__64670;
    wire N__64667;
    wire N__64662;
    wire N__64659;
    wire N__64656;
    wire N__64655;
    wire N__64652;
    wire N__64649;
    wire N__64644;
    wire N__64641;
    wire N__64638;
    wire N__64635;
    wire N__64634;
    wire N__64633;
    wire N__64630;
    wire N__64625;
    wire N__64622;
    wire N__64619;
    wire N__64614;
    wire N__64613;
    wire N__64610;
    wire N__64607;
    wire N__64606;
    wire N__64605;
    wire N__64602;
    wire N__64599;
    wire N__64596;
    wire N__64593;
    wire N__64590;
    wire N__64585;
    wire N__64582;
    wire N__64581;
    wire N__64578;
    wire N__64573;
    wire N__64570;
    wire N__64563;
    wire N__64562;
    wire N__64557;
    wire N__64554;
    wire N__64551;
    wire N__64548;
    wire N__64545;
    wire N__64544;
    wire N__64541;
    wire N__64538;
    wire N__64535;
    wire N__64532;
    wire N__64531;
    wire N__64530;
    wire N__64529;
    wire N__64524;
    wire N__64521;
    wire N__64516;
    wire N__64513;
    wire N__64506;
    wire N__64503;
    wire N__64502;
    wire N__64501;
    wire N__64498;
    wire N__64495;
    wire N__64492;
    wire N__64491;
    wire N__64490;
    wire N__64487;
    wire N__64484;
    wire N__64481;
    wire N__64478;
    wire N__64475;
    wire N__64472;
    wire N__64465;
    wire N__64458;
    wire N__64457;
    wire N__64454;
    wire N__64451;
    wire N__64450;
    wire N__64447;
    wire N__64444;
    wire N__64441;
    wire N__64440;
    wire N__64437;
    wire N__64434;
    wire N__64431;
    wire N__64428;
    wire N__64423;
    wire N__64416;
    wire N__64413;
    wire N__64410;
    wire N__64409;
    wire N__64406;
    wire N__64403;
    wire N__64400;
    wire N__64397;
    wire N__64394;
    wire N__64389;
    wire N__64386;
    wire N__64383;
    wire N__64380;
    wire N__64377;
    wire N__64374;
    wire N__64373;
    wire N__64370;
    wire N__64367;
    wire N__64364;
    wire N__64361;
    wire N__64360;
    wire N__64355;
    wire N__64352;
    wire N__64347;
    wire N__64346;
    wire N__64345;
    wire N__64342;
    wire N__64341;
    wire N__64340;
    wire N__64337;
    wire N__64334;
    wire N__64331;
    wire N__64328;
    wire N__64325;
    wire N__64322;
    wire N__64317;
    wire N__64314;
    wire N__64311;
    wire N__64306;
    wire N__64303;
    wire N__64300;
    wire N__64293;
    wire N__64290;
    wire N__64287;
    wire N__64284;
    wire N__64283;
    wire N__64280;
    wire N__64275;
    wire N__64272;
    wire N__64269;
    wire N__64266;
    wire N__64263;
    wire N__64262;
    wire N__64261;
    wire N__64260;
    wire N__64259;
    wire N__64256;
    wire N__64251;
    wire N__64246;
    wire N__64239;
    wire N__64236;
    wire N__64233;
    wire N__64230;
    wire N__64229;
    wire N__64226;
    wire N__64223;
    wire N__64220;
    wire N__64217;
    wire N__64212;
    wire N__64211;
    wire N__64206;
    wire N__64203;
    wire N__64200;
    wire N__64197;
    wire N__64194;
    wire N__64191;
    wire N__64188;
    wire N__64185;
    wire N__64182;
    wire N__64179;
    wire N__64178;
    wire N__64177;
    wire N__64174;
    wire N__64169;
    wire N__64168;
    wire N__64165;
    wire N__64162;
    wire N__64159;
    wire N__64158;
    wire N__64153;
    wire N__64148;
    wire N__64143;
    wire N__64140;
    wire N__64139;
    wire N__64138;
    wire N__64135;
    wire N__64134;
    wire N__64133;
    wire N__64130;
    wire N__64127;
    wire N__64124;
    wire N__64121;
    wire N__64118;
    wire N__64115;
    wire N__64112;
    wire N__64107;
    wire N__64104;
    wire N__64099;
    wire N__64096;
    wire N__64089;
    wire N__64086;
    wire N__64085;
    wire N__64082;
    wire N__64079;
    wire N__64076;
    wire N__64073;
    wire N__64068;
    wire N__64065;
    wire N__64062;
    wire N__64059;
    wire N__64056;
    wire N__64053;
    wire N__64050;
    wire N__64049;
    wire N__64048;
    wire N__64045;
    wire N__64042;
    wire N__64039;
    wire N__64034;
    wire N__64033;
    wire N__64030;
    wire N__64027;
    wire N__64024;
    wire N__64017;
    wire N__64014;
    wire N__64013;
    wire N__64012;
    wire N__64009;
    wire N__64008;
    wire N__64007;
    wire N__64006;
    wire N__64003;
    wire N__64000;
    wire N__63997;
    wire N__63994;
    wire N__63989;
    wire N__63986;
    wire N__63983;
    wire N__63972;
    wire N__63969;
    wire N__63966;
    wire N__63965;
    wire N__63962;
    wire N__63961;
    wire N__63958;
    wire N__63955;
    wire N__63952;
    wire N__63945;
    wire N__63942;
    wire N__63939;
    wire N__63936;
    wire N__63933;
    wire N__63932;
    wire N__63929;
    wire N__63926;
    wire N__63921;
    wire N__63918;
    wire N__63917;
    wire N__63914;
    wire N__63911;
    wire N__63908;
    wire N__63907;
    wire N__63906;
    wire N__63903;
    wire N__63900;
    wire N__63895;
    wire N__63888;
    wire N__63885;
    wire N__63882;
    wire N__63879;
    wire N__63878;
    wire N__63877;
    wire N__63874;
    wire N__63871;
    wire N__63868;
    wire N__63865;
    wire N__63860;
    wire N__63855;
    wire N__63852;
    wire N__63849;
    wire N__63848;
    wire N__63847;
    wire N__63846;
    wire N__63843;
    wire N__63838;
    wire N__63835;
    wire N__63828;
    wire N__63825;
    wire N__63824;
    wire N__63821;
    wire N__63818;
    wire N__63813;
    wire N__63810;
    wire N__63807;
    wire N__63804;
    wire N__63803;
    wire N__63798;
    wire N__63795;
    wire N__63792;
    wire N__63791;
    wire N__63790;
    wire N__63789;
    wire N__63788;
    wire N__63787;
    wire N__63786;
    wire N__63783;
    wire N__63782;
    wire N__63779;
    wire N__63776;
    wire N__63771;
    wire N__63768;
    wire N__63765;
    wire N__63762;
    wire N__63759;
    wire N__63750;
    wire N__63741;
    wire N__63740;
    wire N__63739;
    wire N__63736;
    wire N__63735;
    wire N__63732;
    wire N__63731;
    wire N__63728;
    wire N__63727;
    wire N__63724;
    wire N__63719;
    wire N__63716;
    wire N__63713;
    wire N__63710;
    wire N__63705;
    wire N__63702;
    wire N__63697;
    wire N__63694;
    wire N__63687;
    wire N__63686;
    wire N__63685;
    wire N__63684;
    wire N__63681;
    wire N__63680;
    wire N__63677;
    wire N__63672;
    wire N__63669;
    wire N__63666;
    wire N__63657;
    wire N__63654;
    wire N__63653;
    wire N__63650;
    wire N__63647;
    wire N__63642;
    wire N__63639;
    wire N__63636;
    wire N__63635;
    wire N__63634;
    wire N__63631;
    wire N__63626;
    wire N__63621;
    wire N__63618;
    wire N__63615;
    wire N__63612;
    wire N__63609;
    wire N__63606;
    wire N__63603;
    wire N__63600;
    wire N__63599;
    wire N__63598;
    wire N__63595;
    wire N__63592;
    wire N__63589;
    wire N__63582;
    wire N__63579;
    wire N__63576;
    wire N__63573;
    wire N__63570;
    wire N__63567;
    wire N__63564;
    wire N__63561;
    wire N__63560;
    wire N__63557;
    wire N__63554;
    wire N__63551;
    wire N__63548;
    wire N__63543;
    wire N__63542;
    wire N__63539;
    wire N__63536;
    wire N__63533;
    wire N__63530;
    wire N__63527;
    wire N__63524;
    wire N__63523;
    wire N__63522;
    wire N__63517;
    wire N__63512;
    wire N__63507;
    wire N__63506;
    wire N__63503;
    wire N__63500;
    wire N__63499;
    wire N__63496;
    wire N__63493;
    wire N__63490;
    wire N__63487;
    wire N__63484;
    wire N__63479;
    wire N__63474;
    wire N__63471;
    wire N__63468;
    wire N__63465;
    wire N__63464;
    wire N__63461;
    wire N__63458;
    wire N__63453;
    wire N__63450;
    wire N__63447;
    wire N__63444;
    wire N__63441;
    wire N__63440;
    wire N__63437;
    wire N__63434;
    wire N__63431;
    wire N__63430;
    wire N__63427;
    wire N__63424;
    wire N__63421;
    wire N__63418;
    wire N__63413;
    wire N__63412;
    wire N__63409;
    wire N__63406;
    wire N__63403;
    wire N__63400;
    wire N__63397;
    wire N__63394;
    wire N__63391;
    wire N__63388;
    wire N__63381;
    wire N__63380;
    wire N__63379;
    wire N__63378;
    wire N__63375;
    wire N__63372;
    wire N__63367;
    wire N__63364;
    wire N__63359;
    wire N__63356;
    wire N__63353;
    wire N__63348;
    wire N__63347;
    wire N__63346;
    wire N__63345;
    wire N__63342;
    wire N__63339;
    wire N__63332;
    wire N__63329;
    wire N__63328;
    wire N__63325;
    wire N__63322;
    wire N__63319;
    wire N__63316;
    wire N__63313;
    wire N__63306;
    wire N__63303;
    wire N__63300;
    wire N__63299;
    wire N__63296;
    wire N__63295;
    wire N__63292;
    wire N__63289;
    wire N__63286;
    wire N__63279;
    wire N__63276;
    wire N__63273;
    wire N__63270;
    wire N__63267;
    wire N__63264;
    wire N__63263;
    wire N__63260;
    wire N__63257;
    wire N__63254;
    wire N__63251;
    wire N__63246;
    wire N__63243;
    wire N__63242;
    wire N__63241;
    wire N__63240;
    wire N__63237;
    wire N__63234;
    wire N__63231;
    wire N__63230;
    wire N__63227;
    wire N__63226;
    wire N__63223;
    wire N__63218;
    wire N__63215;
    wire N__63212;
    wire N__63211;
    wire N__63208;
    wire N__63203;
    wire N__63198;
    wire N__63195;
    wire N__63192;
    wire N__63185;
    wire N__63182;
    wire N__63179;
    wire N__63174;
    wire N__63171;
    wire N__63170;
    wire N__63167;
    wire N__63164;
    wire N__63159;
    wire N__63156;
    wire N__63153;
    wire N__63152;
    wire N__63149;
    wire N__63148;
    wire N__63145;
    wire N__63142;
    wire N__63141;
    wire N__63138;
    wire N__63135;
    wire N__63132;
    wire N__63129;
    wire N__63120;
    wire N__63117;
    wire N__63114;
    wire N__63111;
    wire N__63108;
    wire N__63107;
    wire N__63102;
    wire N__63099;
    wire N__63096;
    wire N__63093;
    wire N__63090;
    wire N__63089;
    wire N__63086;
    wire N__63083;
    wire N__63080;
    wire N__63077;
    wire N__63074;
    wire N__63069;
    wire N__63066;
    wire N__63063;
    wire N__63060;
    wire N__63057;
    wire N__63054;
    wire N__63051;
    wire N__63048;
    wire N__63045;
    wire N__63042;
    wire N__63039;
    wire N__63036;
    wire N__63033;
    wire N__63032;
    wire N__63029;
    wire N__63026;
    wire N__63021;
    wire N__63018;
    wire N__63015;
    wire N__63012;
    wire N__63011;
    wire N__63008;
    wire N__63005;
    wire N__63002;
    wire N__62999;
    wire N__62994;
    wire N__62991;
    wire N__62988;
    wire N__62985;
    wire N__62982;
    wire N__62981;
    wire N__62980;
    wire N__62977;
    wire N__62974;
    wire N__62971;
    wire N__62968;
    wire N__62965;
    wire N__62962;
    wire N__62959;
    wire N__62956;
    wire N__62953;
    wire N__62948;
    wire N__62943;
    wire N__62940;
    wire N__62939;
    wire N__62934;
    wire N__62931;
    wire N__62928;
    wire N__62927;
    wire N__62924;
    wire N__62921;
    wire N__62920;
    wire N__62919;
    wire N__62916;
    wire N__62911;
    wire N__62908;
    wire N__62905;
    wire N__62900;
    wire N__62895;
    wire N__62894;
    wire N__62891;
    wire N__62888;
    wire N__62887;
    wire N__62886;
    wire N__62881;
    wire N__62876;
    wire N__62875;
    wire N__62872;
    wire N__62869;
    wire N__62866;
    wire N__62859;
    wire N__62858;
    wire N__62855;
    wire N__62854;
    wire N__62849;
    wire N__62848;
    wire N__62847;
    wire N__62844;
    wire N__62841;
    wire N__62838;
    wire N__62835;
    wire N__62832;
    wire N__62829;
    wire N__62826;
    wire N__62823;
    wire N__62820;
    wire N__62815;
    wire N__62808;
    wire N__62807;
    wire N__62806;
    wire N__62803;
    wire N__62800;
    wire N__62799;
    wire N__62796;
    wire N__62795;
    wire N__62792;
    wire N__62787;
    wire N__62784;
    wire N__62781;
    wire N__62774;
    wire N__62769;
    wire N__62768;
    wire N__62767;
    wire N__62766;
    wire N__62759;
    wire N__62758;
    wire N__62757;
    wire N__62756;
    wire N__62753;
    wire N__62750;
    wire N__62743;
    wire N__62742;
    wire N__62735;
    wire N__62732;
    wire N__62727;
    wire N__62724;
    wire N__62721;
    wire N__62720;
    wire N__62715;
    wire N__62712;
    wire N__62711;
    wire N__62710;
    wire N__62705;
    wire N__62702;
    wire N__62699;
    wire N__62696;
    wire N__62693;
    wire N__62688;
    wire N__62687;
    wire N__62686;
    wire N__62683;
    wire N__62682;
    wire N__62677;
    wire N__62674;
    wire N__62671;
    wire N__62668;
    wire N__62667;
    wire N__62666;
    wire N__62663;
    wire N__62658;
    wire N__62655;
    wire N__62652;
    wire N__62643;
    wire N__62640;
    wire N__62639;
    wire N__62638;
    wire N__62635;
    wire N__62632;
    wire N__62629;
    wire N__62624;
    wire N__62621;
    wire N__62616;
    wire N__62615;
    wire N__62614;
    wire N__62613;
    wire N__62610;
    wire N__62607;
    wire N__62604;
    wire N__62603;
    wire N__62598;
    wire N__62595;
    wire N__62592;
    wire N__62591;
    wire N__62588;
    wire N__62585;
    wire N__62582;
    wire N__62579;
    wire N__62574;
    wire N__62571;
    wire N__62566;
    wire N__62559;
    wire N__62556;
    wire N__62553;
    wire N__62550;
    wire N__62549;
    wire N__62546;
    wire N__62543;
    wire N__62538;
    wire N__62535;
    wire N__62532;
    wire N__62529;
    wire N__62528;
    wire N__62527;
    wire N__62526;
    wire N__62523;
    wire N__62518;
    wire N__62515;
    wire N__62512;
    wire N__62509;
    wire N__62506;
    wire N__62503;
    wire N__62500;
    wire N__62493;
    wire N__62490;
    wire N__62487;
    wire N__62484;
    wire N__62483;
    wire N__62480;
    wire N__62477;
    wire N__62476;
    wire N__62471;
    wire N__62468;
    wire N__62463;
    wire N__62460;
    wire N__62459;
    wire N__62458;
    wire N__62455;
    wire N__62452;
    wire N__62449;
    wire N__62446;
    wire N__62445;
    wire N__62442;
    wire N__62439;
    wire N__62436;
    wire N__62433;
    wire N__62424;
    wire N__62423;
    wire N__62420;
    wire N__62417;
    wire N__62412;
    wire N__62411;
    wire N__62408;
    wire N__62407;
    wire N__62404;
    wire N__62401;
    wire N__62398;
    wire N__62397;
    wire N__62396;
    wire N__62389;
    wire N__62386;
    wire N__62383;
    wire N__62380;
    wire N__62379;
    wire N__62376;
    wire N__62371;
    wire N__62368;
    wire N__62361;
    wire N__62360;
    wire N__62357;
    wire N__62356;
    wire N__62355;
    wire N__62354;
    wire N__62353;
    wire N__62350;
    wire N__62345;
    wire N__62338;
    wire N__62331;
    wire N__62328;
    wire N__62325;
    wire N__62322;
    wire N__62319;
    wire N__62318;
    wire N__62317;
    wire N__62316;
    wire N__62313;
    wire N__62310;
    wire N__62309;
    wire N__62306;
    wire N__62303;
    wire N__62300;
    wire N__62297;
    wire N__62296;
    wire N__62295;
    wire N__62294;
    wire N__62291;
    wire N__62286;
    wire N__62281;
    wire N__62278;
    wire N__62275;
    wire N__62272;
    wire N__62271;
    wire N__62268;
    wire N__62265;
    wire N__62262;
    wire N__62259;
    wire N__62254;
    wire N__62253;
    wire N__62250;
    wire N__62245;
    wire N__62244;
    wire N__62241;
    wire N__62236;
    wire N__62233;
    wire N__62228;
    wire N__62225;
    wire N__62222;
    wire N__62219;
    wire N__62216;
    wire N__62213;
    wire N__62210;
    wire N__62207;
    wire N__62204;
    wire N__62201;
    wire N__62198;
    wire N__62197;
    wire N__62194;
    wire N__62191;
    wire N__62188;
    wire N__62185;
    wire N__62182;
    wire N__62179;
    wire N__62166;
    wire N__62163;
    wire N__62160;
    wire N__62157;
    wire N__62154;
    wire N__62151;
    wire N__62148;
    wire N__62145;
    wire N__62142;
    wire N__62141;
    wire N__62136;
    wire N__62133;
    wire N__62132;
    wire N__62127;
    wire N__62124;
    wire N__62123;
    wire N__62120;
    wire N__62119;
    wire N__62116;
    wire N__62113;
    wire N__62110;
    wire N__62107;
    wire N__62102;
    wire N__62099;
    wire N__62096;
    wire N__62091;
    wire N__62088;
    wire N__62085;
    wire N__62084;
    wire N__62081;
    wire N__62078;
    wire N__62075;
    wire N__62072;
    wire N__62071;
    wire N__62070;
    wire N__62069;
    wire N__62064;
    wire N__62057;
    wire N__62052;
    wire N__62049;
    wire N__62046;
    wire N__62043;
    wire N__62040;
    wire N__62037;
    wire N__62034;
    wire N__62033;
    wire N__62030;
    wire N__62027;
    wire N__62022;
    wire N__62019;
    wire N__62016;
    wire N__62013;
    wire N__62010;
    wire N__62009;
    wire N__62006;
    wire N__62003;
    wire N__62000;
    wire N__61995;
    wire N__61992;
    wire N__61991;
    wire N__61988;
    wire N__61987;
    wire N__61984;
    wire N__61981;
    wire N__61978;
    wire N__61975;
    wire N__61972;
    wire N__61969;
    wire N__61962;
    wire N__61959;
    wire N__61956;
    wire N__61953;
    wire N__61950;
    wire N__61949;
    wire N__61946;
    wire N__61943;
    wire N__61938;
    wire N__61935;
    wire N__61934;
    wire N__61931;
    wire N__61928;
    wire N__61927;
    wire N__61926;
    wire N__61921;
    wire N__61916;
    wire N__61913;
    wire N__61910;
    wire N__61905;
    wire N__61902;
    wire N__61901;
    wire N__61898;
    wire N__61897;
    wire N__61894;
    wire N__61891;
    wire N__61890;
    wire N__61887;
    wire N__61884;
    wire N__61881;
    wire N__61878;
    wire N__61875;
    wire N__61872;
    wire N__61867;
    wire N__61860;
    wire N__61859;
    wire N__61856;
    wire N__61853;
    wire N__61852;
    wire N__61851;
    wire N__61846;
    wire N__61841;
    wire N__61838;
    wire N__61833;
    wire N__61830;
    wire N__61827;
    wire N__61824;
    wire N__61821;
    wire N__61818;
    wire N__61815;
    wire N__61812;
    wire N__61811;
    wire N__61808;
    wire N__61805;
    wire N__61800;
    wire N__61797;
    wire N__61796;
    wire N__61793;
    wire N__61792;
    wire N__61789;
    wire N__61786;
    wire N__61783;
    wire N__61782;
    wire N__61781;
    wire N__61774;
    wire N__61771;
    wire N__61768;
    wire N__61767;
    wire N__61762;
    wire N__61759;
    wire N__61756;
    wire N__61753;
    wire N__61746;
    wire N__61745;
    wire N__61742;
    wire N__61741;
    wire N__61740;
    wire N__61739;
    wire N__61738;
    wire N__61735;
    wire N__61732;
    wire N__61725;
    wire N__61720;
    wire N__61719;
    wire N__61716;
    wire N__61711;
    wire N__61708;
    wire N__61703;
    wire N__61698;
    wire N__61695;
    wire N__61692;
    wire N__61691;
    wire N__61688;
    wire N__61685;
    wire N__61680;
    wire N__61677;
    wire N__61674;
    wire N__61671;
    wire N__61668;
    wire N__61665;
    wire N__61662;
    wire N__61659;
    wire N__61658;
    wire N__61655;
    wire N__61652;
    wire N__61649;
    wire N__61648;
    wire N__61645;
    wire N__61642;
    wire N__61639;
    wire N__61634;
    wire N__61629;
    wire N__61626;
    wire N__61623;
    wire N__61620;
    wire N__61617;
    wire N__61616;
    wire N__61613;
    wire N__61610;
    wire N__61607;
    wire N__61604;
    wire N__61601;
    wire N__61596;
    wire N__61593;
    wire N__61590;
    wire N__61589;
    wire N__61586;
    wire N__61583;
    wire N__61582;
    wire N__61579;
    wire N__61576;
    wire N__61573;
    wire N__61570;
    wire N__61567;
    wire N__61560;
    wire N__61557;
    wire N__61554;
    wire N__61553;
    wire N__61552;
    wire N__61549;
    wire N__61548;
    wire N__61545;
    wire N__61542;
    wire N__61541;
    wire N__61538;
    wire N__61535;
    wire N__61530;
    wire N__61527;
    wire N__61524;
    wire N__61521;
    wire N__61518;
    wire N__61515;
    wire N__61512;
    wire N__61503;
    wire N__61500;
    wire N__61497;
    wire N__61494;
    wire N__61491;
    wire N__61488;
    wire N__61487;
    wire N__61482;
    wire N__61479;
    wire N__61476;
    wire N__61475;
    wire N__61470;
    wire N__61467;
    wire N__61466;
    wire N__61463;
    wire N__61460;
    wire N__61457;
    wire N__61454;
    wire N__61451;
    wire N__61448;
    wire N__61443;
    wire N__61440;
    wire N__61437;
    wire N__61434;
    wire N__61433;
    wire N__61430;
    wire N__61429;
    wire N__61426;
    wire N__61425;
    wire N__61424;
    wire N__61421;
    wire N__61418;
    wire N__61415;
    wire N__61412;
    wire N__61409;
    wire N__61404;
    wire N__61399;
    wire N__61392;
    wire N__61391;
    wire N__61388;
    wire N__61385;
    wire N__61384;
    wire N__61381;
    wire N__61380;
    wire N__61377;
    wire N__61374;
    wire N__61371;
    wire N__61368;
    wire N__61363;
    wire N__61360;
    wire N__61357;
    wire N__61352;
    wire N__61347;
    wire N__61344;
    wire N__61341;
    wire N__61338;
    wire N__61335;
    wire N__61334;
    wire N__61333;
    wire N__61330;
    wire N__61327;
    wire N__61324;
    wire N__61321;
    wire N__61316;
    wire N__61313;
    wire N__61310;
    wire N__61305;
    wire N__61302;
    wire N__61299;
    wire N__61298;
    wire N__61295;
    wire N__61294;
    wire N__61293;
    wire N__61292;
    wire N__61289;
    wire N__61288;
    wire N__61285;
    wire N__61282;
    wire N__61277;
    wire N__61272;
    wire N__61263;
    wire N__61262;
    wire N__61259;
    wire N__61256;
    wire N__61255;
    wire N__61252;
    wire N__61249;
    wire N__61246;
    wire N__61245;
    wire N__61242;
    wire N__61239;
    wire N__61236;
    wire N__61235;
    wire N__61232;
    wire N__61227;
    wire N__61224;
    wire N__61221;
    wire N__61212;
    wire N__61209;
    wire N__61206;
    wire N__61203;
    wire N__61200;
    wire N__61197;
    wire N__61194;
    wire N__61191;
    wire N__61188;
    wire N__61185;
    wire N__61182;
    wire N__61179;
    wire N__61176;
    wire N__61175;
    wire N__61172;
    wire N__61169;
    wire N__61166;
    wire N__61163;
    wire N__61160;
    wire N__61157;
    wire N__61152;
    wire N__61149;
    wire N__61146;
    wire N__61143;
    wire N__61142;
    wire N__61139;
    wire N__61136;
    wire N__61133;
    wire N__61128;
    wire N__61125;
    wire N__61122;
    wire N__61119;
    wire N__61116;
    wire N__61113;
    wire N__61112;
    wire N__61111;
    wire N__61104;
    wire N__61101;
    wire N__61098;
    wire N__61095;
    wire N__61094;
    wire N__61091;
    wire N__61088;
    wire N__61083;
    wire N__61080;
    wire N__61077;
    wire N__61074;
    wire N__61071;
    wire N__61068;
    wire N__61065;
    wire N__61064;
    wire N__61061;
    wire N__61058;
    wire N__61057;
    wire N__61054;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61044;
    wire N__61043;
    wire N__61040;
    wire N__61037;
    wire N__61036;
    wire N__61035;
    wire N__61032;
    wire N__61031;
    wire N__61030;
    wire N__61025;
    wire N__61020;
    wire N__61017;
    wire N__61014;
    wire N__61011;
    wire N__61008;
    wire N__61005;
    wire N__60998;
    wire N__60987;
    wire N__60984;
    wire N__60981;
    wire N__60978;
    wire N__60975;
    wire N__60972;
    wire N__60969;
    wire N__60966;
    wire N__60963;
    wire N__60960;
    wire N__60957;
    wire N__60954;
    wire N__60953;
    wire N__60952;
    wire N__60949;
    wire N__60946;
    wire N__60943;
    wire N__60942;
    wire N__60939;
    wire N__60934;
    wire N__60931;
    wire N__60924;
    wire N__60921;
    wire N__60918;
    wire N__60915;
    wire N__60912;
    wire N__60909;
    wire N__60906;
    wire N__60905;
    wire N__60900;
    wire N__60899;
    wire N__60896;
    wire N__60895;
    wire N__60892;
    wire N__60891;
    wire N__60888;
    wire N__60885;
    wire N__60884;
    wire N__60883;
    wire N__60882;
    wire N__60877;
    wire N__60874;
    wire N__60867;
    wire N__60864;
    wire N__60855;
    wire N__60854;
    wire N__60851;
    wire N__60850;
    wire N__60847;
    wire N__60844;
    wire N__60841;
    wire N__60836;
    wire N__60835;
    wire N__60834;
    wire N__60829;
    wire N__60824;
    wire N__60819;
    wire N__60818;
    wire N__60817;
    wire N__60814;
    wire N__60809;
    wire N__60806;
    wire N__60803;
    wire N__60798;
    wire N__60797;
    wire N__60796;
    wire N__60793;
    wire N__60792;
    wire N__60789;
    wire N__60786;
    wire N__60783;
    wire N__60780;
    wire N__60775;
    wire N__60774;
    wire N__60773;
    wire N__60770;
    wire N__60765;
    wire N__60760;
    wire N__60753;
    wire N__60750;
    wire N__60747;
    wire N__60746;
    wire N__60743;
    wire N__60742;
    wire N__60741;
    wire N__60738;
    wire N__60737;
    wire N__60734;
    wire N__60731;
    wire N__60728;
    wire N__60723;
    wire N__60714;
    wire N__60711;
    wire N__60708;
    wire N__60705;
    wire N__60702;
    wire N__60699;
    wire N__60696;
    wire N__60693;
    wire N__60690;
    wire N__60687;
    wire N__60686;
    wire N__60683;
    wire N__60680;
    wire N__60677;
    wire N__60674;
    wire N__60671;
    wire N__60666;
    wire N__60663;
    wire N__60660;
    wire N__60657;
    wire N__60654;
    wire N__60651;
    wire N__60648;
    wire N__60645;
    wire N__60644;
    wire N__60641;
    wire N__60638;
    wire N__60637;
    wire N__60636;
    wire N__60635;
    wire N__60634;
    wire N__60633;
    wire N__60632;
    wire N__60631;
    wire N__60628;
    wire N__60625;
    wire N__60620;
    wire N__60617;
    wire N__60610;
    wire N__60607;
    wire N__60594;
    wire N__60591;
    wire N__60588;
    wire N__60585;
    wire N__60582;
    wire N__60579;
    wire N__60576;
    wire N__60573;
    wire N__60570;
    wire N__60567;
    wire N__60566;
    wire N__60563;
    wire N__60562;
    wire N__60559;
    wire N__60558;
    wire N__60557;
    wire N__60554;
    wire N__60553;
    wire N__60552;
    wire N__60549;
    wire N__60548;
    wire N__60547;
    wire N__60546;
    wire N__60545;
    wire N__60542;
    wire N__60537;
    wire N__60536;
    wire N__60535;
    wire N__60534;
    wire N__60533;
    wire N__60530;
    wire N__60527;
    wire N__60524;
    wire N__60521;
    wire N__60518;
    wire N__60515;
    wire N__60512;
    wire N__60511;
    wire N__60508;
    wire N__60507;
    wire N__60504;
    wire N__60501;
    wire N__60494;
    wire N__60491;
    wire N__60490;
    wire N__60481;
    wire N__60478;
    wire N__60475;
    wire N__60470;
    wire N__60465;
    wire N__60458;
    wire N__60453;
    wire N__60438;
    wire N__60435;
    wire N__60432;
    wire N__60431;
    wire N__60428;
    wire N__60427;
    wire N__60424;
    wire N__60421;
    wire N__60418;
    wire N__60417;
    wire N__60416;
    wire N__60415;
    wire N__60414;
    wire N__60413;
    wire N__60410;
    wire N__60409;
    wire N__60408;
    wire N__60405;
    wire N__60394;
    wire N__60391;
    wire N__60388;
    wire N__60387;
    wire N__60386;
    wire N__60385;
    wire N__60382;
    wire N__60379;
    wire N__60378;
    wire N__60377;
    wire N__60372;
    wire N__60369;
    wire N__60366;
    wire N__60363;
    wire N__60360;
    wire N__60357;
    wire N__60354;
    wire N__60347;
    wire N__60342;
    wire N__60327;
    wire N__60324;
    wire N__60321;
    wire N__60318;
    wire N__60315;
    wire N__60312;
    wire N__60309;
    wire N__60306;
    wire N__60305;
    wire N__60304;
    wire N__60303;
    wire N__60302;
    wire N__60301;
    wire N__60298;
    wire N__60297;
    wire N__60296;
    wire N__60295;
    wire N__60292;
    wire N__60289;
    wire N__60284;
    wire N__60283;
    wire N__60280;
    wire N__60277;
    wire N__60274;
    wire N__60269;
    wire N__60266;
    wire N__60261;
    wire N__60258;
    wire N__60243;
    wire N__60240;
    wire N__60239;
    wire N__60236;
    wire N__60235;
    wire N__60234;
    wire N__60231;
    wire N__60230;
    wire N__60229;
    wire N__60228;
    wire N__60227;
    wire N__60224;
    wire N__60219;
    wire N__60212;
    wire N__60209;
    wire N__60208;
    wire N__60205;
    wire N__60204;
    wire N__60203;
    wire N__60198;
    wire N__60195;
    wire N__60188;
    wire N__60187;
    wire N__60186;
    wire N__60183;
    wire N__60180;
    wire N__60173;
    wire N__60168;
    wire N__60159;
    wire N__60156;
    wire N__60155;
    wire N__60152;
    wire N__60149;
    wire N__60148;
    wire N__60143;
    wire N__60140;
    wire N__60135;
    wire N__60132;
    wire N__60131;
    wire N__60128;
    wire N__60125;
    wire N__60120;
    wire N__60117;
    wire N__60116;
    wire N__60113;
    wire N__60110;
    wire N__60107;
    wire N__60102;
    wire N__60099;
    wire N__60096;
    wire N__60093;
    wire N__60090;
    wire N__60087;
    wire N__60084;
    wire N__60081;
    wire N__60080;
    wire N__60077;
    wire N__60074;
    wire N__60071;
    wire N__60068;
    wire N__60063;
    wire N__60062;
    wire N__60061;
    wire N__60060;
    wire N__60057;
    wire N__60054;
    wire N__60049;
    wire N__60048;
    wire N__60045;
    wire N__60040;
    wire N__60037;
    wire N__60030;
    wire N__60029;
    wire N__60026;
    wire N__60023;
    wire N__60020;
    wire N__60017;
    wire N__60012;
    wire N__60009;
    wire N__60006;
    wire N__60003;
    wire N__60000;
    wire N__59997;
    wire N__59994;
    wire N__59991;
    wire N__59988;
    wire N__59985;
    wire N__59982;
    wire N__59979;
    wire N__59976;
    wire N__59973;
    wire N__59970;
    wire N__59967;
    wire N__59964;
    wire N__59961;
    wire N__59958;
    wire N__59955;
    wire N__59952;
    wire N__59949;
    wire N__59946;
    wire N__59943;
    wire N__59940;
    wire N__59937;
    wire N__59934;
    wire N__59931;
    wire N__59928;
    wire N__59925;
    wire N__59922;
    wire N__59919;
    wire N__59916;
    wire N__59913;
    wire N__59912;
    wire N__59909;
    wire N__59906;
    wire N__59901;
    wire N__59898;
    wire N__59897;
    wire N__59896;
    wire N__59893;
    wire N__59890;
    wire N__59887;
    wire N__59880;
    wire N__59877;
    wire N__59876;
    wire N__59875;
    wire N__59872;
    wire N__59869;
    wire N__59868;
    wire N__59867;
    wire N__59864;
    wire N__59861;
    wire N__59858;
    wire N__59853;
    wire N__59850;
    wire N__59845;
    wire N__59838;
    wire N__59835;
    wire N__59832;
    wire N__59829;
    wire N__59826;
    wire N__59823;
    wire N__59820;
    wire N__59817;
    wire N__59814;
    wire N__59811;
    wire N__59808;
    wire N__59805;
    wire N__59802;
    wire N__59799;
    wire N__59796;
    wire N__59793;
    wire N__59790;
    wire N__59787;
    wire N__59786;
    wire N__59783;
    wire N__59782;
    wire N__59777;
    wire N__59774;
    wire N__59771;
    wire N__59768;
    wire N__59763;
    wire N__59760;
    wire N__59757;
    wire N__59754;
    wire N__59751;
    wire N__59748;
    wire N__59745;
    wire N__59742;
    wire N__59739;
    wire N__59738;
    wire N__59735;
    wire N__59732;
    wire N__59731;
    wire N__59730;
    wire N__59725;
    wire N__59724;
    wire N__59721;
    wire N__59720;
    wire N__59717;
    wire N__59714;
    wire N__59711;
    wire N__59706;
    wire N__59703;
    wire N__59702;
    wire N__59699;
    wire N__59692;
    wire N__59689;
    wire N__59686;
    wire N__59683;
    wire N__59676;
    wire N__59673;
    wire N__59670;
    wire N__59667;
    wire N__59664;
    wire N__59663;
    wire N__59660;
    wire N__59657;
    wire N__59654;
    wire N__59651;
    wire N__59648;
    wire N__59645;
    wire N__59640;
    wire N__59637;
    wire N__59636;
    wire N__59633;
    wire N__59630;
    wire N__59629;
    wire N__59628;
    wire N__59625;
    wire N__59622;
    wire N__59619;
    wire N__59616;
    wire N__59613;
    wire N__59610;
    wire N__59607;
    wire N__59604;
    wire N__59601;
    wire N__59598;
    wire N__59589;
    wire N__59588;
    wire N__59587;
    wire N__59582;
    wire N__59579;
    wire N__59578;
    wire N__59575;
    wire N__59570;
    wire N__59567;
    wire N__59562;
    wire N__59561;
    wire N__59558;
    wire N__59557;
    wire N__59556;
    wire N__59553;
    wire N__59550;
    wire N__59545;
    wire N__59542;
    wire N__59539;
    wire N__59532;
    wire N__59529;
    wire N__59526;
    wire N__59525;
    wire N__59524;
    wire N__59521;
    wire N__59516;
    wire N__59513;
    wire N__59508;
    wire N__59505;
    wire N__59502;
    wire N__59499;
    wire N__59496;
    wire N__59493;
    wire N__59490;
    wire N__59487;
    wire N__59484;
    wire N__59481;
    wire N__59480;
    wire N__59479;
    wire N__59476;
    wire N__59471;
    wire N__59468;
    wire N__59463;
    wire N__59460;
    wire N__59457;
    wire N__59456;
    wire N__59453;
    wire N__59450;
    wire N__59445;
    wire N__59442;
    wire N__59441;
    wire N__59440;
    wire N__59435;
    wire N__59434;
    wire N__59433;
    wire N__59430;
    wire N__59427;
    wire N__59424;
    wire N__59421;
    wire N__59418;
    wire N__59415;
    wire N__59412;
    wire N__59403;
    wire N__59400;
    wire N__59397;
    wire N__59394;
    wire N__59391;
    wire N__59388;
    wire N__59385;
    wire N__59382;
    wire N__59379;
    wire N__59376;
    wire N__59373;
    wire N__59370;
    wire N__59367;
    wire N__59366;
    wire N__59363;
    wire N__59360;
    wire N__59355;
    wire N__59352;
    wire N__59349;
    wire N__59348;
    wire N__59345;
    wire N__59342;
    wire N__59339;
    wire N__59334;
    wire N__59333;
    wire N__59330;
    wire N__59329;
    wire N__59326;
    wire N__59321;
    wire N__59316;
    wire N__59313;
    wire N__59310;
    wire N__59307;
    wire N__59304;
    wire N__59301;
    wire N__59300;
    wire N__59297;
    wire N__59294;
    wire N__59289;
    wire N__59286;
    wire N__59283;
    wire N__59282;
    wire N__59281;
    wire N__59280;
    wire N__59277;
    wire N__59270;
    wire N__59265;
    wire N__59262;
    wire N__59261;
    wire N__59260;
    wire N__59259;
    wire N__59256;
    wire N__59253;
    wire N__59250;
    wire N__59247;
    wire N__59244;
    wire N__59243;
    wire N__59240;
    wire N__59237;
    wire N__59232;
    wire N__59231;
    wire N__59228;
    wire N__59225;
    wire N__59220;
    wire N__59215;
    wire N__59208;
    wire N__59207;
    wire N__59206;
    wire N__59205;
    wire N__59202;
    wire N__59199;
    wire N__59198;
    wire N__59197;
    wire N__59194;
    wire N__59191;
    wire N__59190;
    wire N__59187;
    wire N__59184;
    wire N__59179;
    wire N__59176;
    wire N__59173;
    wire N__59170;
    wire N__59165;
    wire N__59162;
    wire N__59157;
    wire N__59154;
    wire N__59149;
    wire N__59148;
    wire N__59143;
    wire N__59140;
    wire N__59137;
    wire N__59130;
    wire N__59129;
    wire N__59126;
    wire N__59125;
    wire N__59122;
    wire N__59119;
    wire N__59116;
    wire N__59109;
    wire N__59106;
    wire N__59105;
    wire N__59102;
    wire N__59099;
    wire N__59096;
    wire N__59093;
    wire N__59088;
    wire N__59085;
    wire N__59082;
    wire N__59081;
    wire N__59078;
    wire N__59075;
    wire N__59072;
    wire N__59069;
    wire N__59064;
    wire N__59061;
    wire N__59058;
    wire N__59057;
    wire N__59054;
    wire N__59053;
    wire N__59050;
    wire N__59047;
    wire N__59044;
    wire N__59039;
    wire N__59034;
    wire N__59031;
    wire N__59028;
    wire N__59025;
    wire N__59022;
    wire N__59019;
    wire N__59018;
    wire N__59015;
    wire N__59012;
    wire N__59011;
    wire N__59010;
    wire N__59005;
    wire N__59002;
    wire N__59001;
    wire N__58998;
    wire N__58995;
    wire N__58990;
    wire N__58983;
    wire N__58980;
    wire N__58979;
    wire N__58974;
    wire N__58971;
    wire N__58968;
    wire N__58967;
    wire N__58966;
    wire N__58963;
    wire N__58960;
    wire N__58957;
    wire N__58952;
    wire N__58949;
    wire N__58946;
    wire N__58943;
    wire N__58938;
    wire N__58937;
    wire N__58934;
    wire N__58931;
    wire N__58930;
    wire N__58927;
    wire N__58924;
    wire N__58921;
    wire N__58918;
    wire N__58915;
    wire N__58912;
    wire N__58907;
    wire N__58902;
    wire N__58899;
    wire N__58896;
    wire N__58893;
    wire N__58892;
    wire N__58891;
    wire N__58890;
    wire N__58887;
    wire N__58884;
    wire N__58879;
    wire N__58872;
    wire N__58871;
    wire N__58868;
    wire N__58865;
    wire N__58862;
    wire N__58859;
    wire N__58854;
    wire N__58851;
    wire N__58848;
    wire N__58847;
    wire N__58844;
    wire N__58843;
    wire N__58836;
    wire N__58833;
    wire N__58830;
    wire N__58829;
    wire N__58828;
    wire N__58825;
    wire N__58822;
    wire N__58821;
    wire N__58818;
    wire N__58815;
    wire N__58810;
    wire N__58803;
    wire N__58800;
    wire N__58797;
    wire N__58794;
    wire N__58791;
    wire N__58788;
    wire N__58785;
    wire N__58782;
    wire N__58779;
    wire N__58778;
    wire N__58777;
    wire N__58776;
    wire N__58775;
    wire N__58768;
    wire N__58767;
    wire N__58764;
    wire N__58761;
    wire N__58758;
    wire N__58755;
    wire N__58752;
    wire N__58751;
    wire N__58748;
    wire N__58743;
    wire N__58740;
    wire N__58737;
    wire N__58732;
    wire N__58725;
    wire N__58722;
    wire N__58719;
    wire N__58716;
    wire N__58715;
    wire N__58712;
    wire N__58709;
    wire N__58704;
    wire N__58701;
    wire N__58700;
    wire N__58697;
    wire N__58694;
    wire N__58689;
    wire N__58686;
    wire N__58683;
    wire N__58680;
    wire N__58677;
    wire N__58674;
    wire N__58671;
    wire N__58670;
    wire N__58669;
    wire N__58666;
    wire N__58663;
    wire N__58662;
    wire N__58659;
    wire N__58656;
    wire N__58651;
    wire N__58646;
    wire N__58643;
    wire N__58638;
    wire N__58635;
    wire N__58632;
    wire N__58629;
    wire N__58626;
    wire N__58623;
    wire N__58620;
    wire N__58619;
    wire N__58618;
    wire N__58615;
    wire N__58614;
    wire N__58611;
    wire N__58608;
    wire N__58605;
    wire N__58602;
    wire N__58599;
    wire N__58594;
    wire N__58587;
    wire N__58584;
    wire N__58581;
    wire N__58578;
    wire N__58575;
    wire N__58572;
    wire N__58569;
    wire N__58566;
    wire N__58563;
    wire N__58560;
    wire N__58557;
    wire N__58554;
    wire N__58551;
    wire N__58548;
    wire N__58545;
    wire N__58544;
    wire N__58541;
    wire N__58538;
    wire N__58535;
    wire N__58532;
    wire N__58527;
    wire N__58524;
    wire N__58523;
    wire N__58520;
    wire N__58517;
    wire N__58514;
    wire N__58511;
    wire N__58506;
    wire N__58503;
    wire N__58500;
    wire N__58497;
    wire N__58496;
    wire N__58493;
    wire N__58490;
    wire N__58485;
    wire N__58482;
    wire N__58479;
    wire N__58476;
    wire N__58473;
    wire N__58472;
    wire N__58469;
    wire N__58466;
    wire N__58461;
    wire N__58458;
    wire N__58455;
    wire N__58452;
    wire N__58451;
    wire N__58448;
    wire N__58447;
    wire N__58444;
    wire N__58441;
    wire N__58438;
    wire N__58435;
    wire N__58430;
    wire N__58425;
    wire N__58422;
    wire N__58419;
    wire N__58416;
    wire N__58413;
    wire N__58410;
    wire N__58407;
    wire N__58404;
    wire N__58403;
    wire N__58400;
    wire N__58399;
    wire N__58396;
    wire N__58395;
    wire N__58392;
    wire N__58387;
    wire N__58384;
    wire N__58377;
    wire N__58374;
    wire N__58373;
    wire N__58372;
    wire N__58369;
    wire N__58366;
    wire N__58363;
    wire N__58360;
    wire N__58355;
    wire N__58350;
    wire N__58347;
    wire N__58344;
    wire N__58341;
    wire N__58338;
    wire N__58335;
    wire N__58332;
    wire N__58331;
    wire N__58326;
    wire N__58323;
    wire N__58320;
    wire N__58317;
    wire N__58314;
    wire N__58313;
    wire N__58308;
    wire N__58305;
    wire N__58304;
    wire N__58301;
    wire N__58298;
    wire N__58295;
    wire N__58292;
    wire N__58289;
    wire N__58284;
    wire N__58281;
    wire N__58280;
    wire N__58279;
    wire N__58274;
    wire N__58271;
    wire N__58268;
    wire N__58263;
    wire N__58260;
    wire N__58257;
    wire N__58254;
    wire N__58253;
    wire N__58250;
    wire N__58247;
    wire N__58242;
    wire N__58239;
    wire N__58236;
    wire N__58233;
    wire N__58230;
    wire N__58227;
    wire N__58224;
    wire N__58221;
    wire N__58218;
    wire N__58215;
    wire N__58212;
    wire N__58209;
    wire N__58206;
    wire N__58203;
    wire N__58200;
    wire N__58199;
    wire N__58196;
    wire N__58193;
    wire N__58190;
    wire N__58187;
    wire N__58184;
    wire N__58181;
    wire N__58178;
    wire N__58173;
    wire N__58170;
    wire N__58169;
    wire N__58166;
    wire N__58163;
    wire N__58162;
    wire N__58159;
    wire N__58156;
    wire N__58155;
    wire N__58152;
    wire N__58147;
    wire N__58144;
    wire N__58137;
    wire N__58136;
    wire N__58133;
    wire N__58132;
    wire N__58129;
    wire N__58128;
    wire N__58125;
    wire N__58122;
    wire N__58119;
    wire N__58116;
    wire N__58113;
    wire N__58108;
    wire N__58101;
    wire N__58098;
    wire N__58097;
    wire N__58094;
    wire N__58091;
    wire N__58090;
    wire N__58087;
    wire N__58084;
    wire N__58081;
    wire N__58080;
    wire N__58079;
    wire N__58078;
    wire N__58075;
    wire N__58072;
    wire N__58063;
    wire N__58056;
    wire N__58055;
    wire N__58054;
    wire N__58053;
    wire N__58052;
    wire N__58051;
    wire N__58050;
    wire N__58049;
    wire N__58048;
    wire N__58047;
    wire N__58044;
    wire N__58043;
    wire N__58040;
    wire N__58037;
    wire N__58026;
    wire N__58021;
    wire N__58018;
    wire N__58015;
    wire N__58014;
    wire N__58013;
    wire N__58012;
    wire N__58009;
    wire N__58002;
    wire N__57999;
    wire N__57996;
    wire N__57993;
    wire N__57988;
    wire N__57983;
    wire N__57972;
    wire N__57969;
    wire N__57966;
    wire N__57963;
    wire N__57960;
    wire N__57959;
    wire N__57958;
    wire N__57957;
    wire N__57952;
    wire N__57951;
    wire N__57950;
    wire N__57949;
    wire N__57946;
    wire N__57943;
    wire N__57942;
    wire N__57939;
    wire N__57934;
    wire N__57931;
    wire N__57930;
    wire N__57925;
    wire N__57922;
    wire N__57917;
    wire N__57912;
    wire N__57909;
    wire N__57900;
    wire N__57897;
    wire N__57894;
    wire N__57891;
    wire N__57888;
    wire N__57887;
    wire N__57886;
    wire N__57883;
    wire N__57878;
    wire N__57875;
    wire N__57872;
    wire N__57869;
    wire N__57864;
    wire N__57861;
    wire N__57858;
    wire N__57855;
    wire N__57852;
    wire N__57849;
    wire N__57846;
    wire N__57843;
    wire N__57840;
    wire N__57837;
    wire N__57834;
    wire N__57831;
    wire N__57828;
    wire N__57825;
    wire N__57822;
    wire N__57819;
    wire N__57816;
    wire N__57813;
    wire N__57810;
    wire N__57807;
    wire N__57804;
    wire N__57801;
    wire N__57800;
    wire N__57797;
    wire N__57794;
    wire N__57791;
    wire N__57788;
    wire N__57783;
    wire N__57782;
    wire N__57779;
    wire N__57776;
    wire N__57773;
    wire N__57768;
    wire N__57765;
    wire N__57762;
    wire N__57759;
    wire N__57756;
    wire N__57753;
    wire N__57750;
    wire N__57747;
    wire N__57744;
    wire N__57741;
    wire N__57738;
    wire N__57735;
    wire N__57732;
    wire N__57731;
    wire N__57730;
    wire N__57729;
    wire N__57728;
    wire N__57725;
    wire N__57722;
    wire N__57721;
    wire N__57714;
    wire N__57711;
    wire N__57708;
    wire N__57705;
    wire N__57702;
    wire N__57699;
    wire N__57694;
    wire N__57691;
    wire N__57684;
    wire N__57683;
    wire N__57678;
    wire N__57675;
    wire N__57672;
    wire N__57671;
    wire N__57668;
    wire N__57667;
    wire N__57664;
    wire N__57663;
    wire N__57662;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57650;
    wire N__57647;
    wire N__57644;
    wire N__57639;
    wire N__57638;
    wire N__57637;
    wire N__57636;
    wire N__57633;
    wire N__57628;
    wire N__57625;
    wire N__57620;
    wire N__57617;
    wire N__57606;
    wire N__57603;
    wire N__57600;
    wire N__57597;
    wire N__57594;
    wire N__57593;
    wire N__57592;
    wire N__57589;
    wire N__57584;
    wire N__57579;
    wire N__57576;
    wire N__57573;
    wire N__57570;
    wire N__57567;
    wire N__57564;
    wire N__57563;
    wire N__57562;
    wire N__57559;
    wire N__57554;
    wire N__57551;
    wire N__57548;
    wire N__57545;
    wire N__57542;
    wire N__57537;
    wire N__57536;
    wire N__57535;
    wire N__57532;
    wire N__57529;
    wire N__57526;
    wire N__57523;
    wire N__57520;
    wire N__57517;
    wire N__57510;
    wire N__57507;
    wire N__57504;
    wire N__57501;
    wire N__57498;
    wire N__57495;
    wire N__57494;
    wire N__57489;
    wire N__57488;
    wire N__57485;
    wire N__57484;
    wire N__57483;
    wire N__57480;
    wire N__57477;
    wire N__57474;
    wire N__57469;
    wire N__57462;
    wire N__57461;
    wire N__57460;
    wire N__57457;
    wire N__57450;
    wire N__57447;
    wire N__57444;
    wire N__57441;
    wire N__57438;
    wire N__57435;
    wire N__57432;
    wire N__57429;
    wire N__57428;
    wire N__57425;
    wire N__57422;
    wire N__57417;
    wire N__57416;
    wire N__57413;
    wire N__57410;
    wire N__57409;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57399;
    wire N__57396;
    wire N__57393;
    wire N__57388;
    wire N__57381;
    wire N__57378;
    wire N__57377;
    wire N__57376;
    wire N__57373;
    wire N__57370;
    wire N__57367;
    wire N__57366;
    wire N__57365;
    wire N__57362;
    wire N__57359;
    wire N__57356;
    wire N__57355;
    wire N__57352;
    wire N__57349;
    wire N__57346;
    wire N__57343;
    wire N__57340;
    wire N__57337;
    wire N__57324;
    wire N__57323;
    wire N__57322;
    wire N__57319;
    wire N__57314;
    wire N__57309;
    wire N__57308;
    wire N__57305;
    wire N__57302;
    wire N__57299;
    wire N__57298;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57286;
    wire N__57283;
    wire N__57280;
    wire N__57277;
    wire N__57270;
    wire N__57267;
    wire N__57264;
    wire N__57263;
    wire N__57260;
    wire N__57257;
    wire N__57254;
    wire N__57251;
    wire N__57246;
    wire N__57245;
    wire N__57244;
    wire N__57243;
    wire N__57240;
    wire N__57237;
    wire N__57236;
    wire N__57235;
    wire N__57234;
    wire N__57233;
    wire N__57232;
    wire N__57229;
    wire N__57228;
    wire N__57225;
    wire N__57220;
    wire N__57213;
    wire N__57208;
    wire N__57203;
    wire N__57192;
    wire N__57189;
    wire N__57186;
    wire N__57183;
    wire N__57180;
    wire N__57177;
    wire N__57174;
    wire N__57171;
    wire N__57168;
    wire N__57165;
    wire N__57162;
    wire N__57159;
    wire N__57156;
    wire N__57155;
    wire N__57152;
    wire N__57149;
    wire N__57146;
    wire N__57143;
    wire N__57140;
    wire N__57137;
    wire N__57134;
    wire N__57129;
    wire N__57126;
    wire N__57123;
    wire N__57120;
    wire N__57117;
    wire N__57114;
    wire N__57113;
    wire N__57112;
    wire N__57109;
    wire N__57106;
    wire N__57103;
    wire N__57102;
    wire N__57099;
    wire N__57096;
    wire N__57091;
    wire N__57088;
    wire N__57081;
    wire N__57080;
    wire N__57077;
    wire N__57076;
    wire N__57073;
    wire N__57072;
    wire N__57069;
    wire N__57066;
    wire N__57063;
    wire N__57060;
    wire N__57053;
    wire N__57048;
    wire N__57045;
    wire N__57042;
    wire N__57039;
    wire N__57036;
    wire N__57033;
    wire N__57030;
    wire N__57027;
    wire N__57024;
    wire N__57021;
    wire N__57018;
    wire N__57017;
    wire N__57016;
    wire N__57015;
    wire N__57014;
    wire N__57011;
    wire N__57002;
    wire N__57001;
    wire N__56998;
    wire N__56995;
    wire N__56994;
    wire N__56991;
    wire N__56988;
    wire N__56985;
    wire N__56980;
    wire N__56973;
    wire N__56970;
    wire N__56967;
    wire N__56964;
    wire N__56961;
    wire N__56958;
    wire N__56955;
    wire N__56952;
    wire N__56949;
    wire N__56946;
    wire N__56943;
    wire N__56940;
    wire N__56937;
    wire N__56934;
    wire N__56931;
    wire N__56928;
    wire N__56925;
    wire N__56922;
    wire N__56919;
    wire N__56916;
    wire N__56913;
    wire N__56910;
    wire N__56907;
    wire N__56904;
    wire N__56903;
    wire N__56898;
    wire N__56895;
    wire N__56894;
    wire N__56893;
    wire N__56890;
    wire N__56887;
    wire N__56886;
    wire N__56883;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56869;
    wire N__56862;
    wire N__56859;
    wire N__56858;
    wire N__56855;
    wire N__56854;
    wire N__56853;
    wire N__56850;
    wire N__56847;
    wire N__56844;
    wire N__56841;
    wire N__56836;
    wire N__56833;
    wire N__56830;
    wire N__56827;
    wire N__56824;
    wire N__56817;
    wire N__56816;
    wire N__56815;
    wire N__56814;
    wire N__56811;
    wire N__56808;
    wire N__56805;
    wire N__56802;
    wire N__56799;
    wire N__56798;
    wire N__56797;
    wire N__56794;
    wire N__56791;
    wire N__56788;
    wire N__56785;
    wire N__56780;
    wire N__56773;
    wire N__56766;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56754;
    wire N__56753;
    wire N__56752;
    wire N__56751;
    wire N__56748;
    wire N__56745;
    wire N__56742;
    wire N__56739;
    wire N__56738;
    wire N__56737;
    wire N__56736;
    wire N__56733;
    wire N__56726;
    wire N__56719;
    wire N__56712;
    wire N__56709;
    wire N__56706;
    wire N__56705;
    wire N__56702;
    wire N__56699;
    wire N__56696;
    wire N__56691;
    wire N__56688;
    wire N__56685;
    wire N__56684;
    wire N__56681;
    wire N__56678;
    wire N__56675;
    wire N__56670;
    wire N__56669;
    wire N__56666;
    wire N__56663;
    wire N__56658;
    wire N__56655;
    wire N__56652;
    wire N__56651;
    wire N__56650;
    wire N__56649;
    wire N__56642;
    wire N__56639;
    wire N__56636;
    wire N__56633;
    wire N__56632;
    wire N__56629;
    wire N__56626;
    wire N__56623;
    wire N__56620;
    wire N__56617;
    wire N__56610;
    wire N__56607;
    wire N__56604;
    wire N__56601;
    wire N__56598;
    wire N__56595;
    wire N__56594;
    wire N__56589;
    wire N__56588;
    wire N__56585;
    wire N__56582;
    wire N__56579;
    wire N__56574;
    wire N__56573;
    wire N__56572;
    wire N__56569;
    wire N__56564;
    wire N__56561;
    wire N__56560;
    wire N__56557;
    wire N__56554;
    wire N__56551;
    wire N__56548;
    wire N__56545;
    wire N__56542;
    wire N__56539;
    wire N__56536;
    wire N__56529;
    wire N__56526;
    wire N__56523;
    wire N__56522;
    wire N__56519;
    wire N__56516;
    wire N__56515;
    wire N__56512;
    wire N__56509;
    wire N__56506;
    wire N__56499;
    wire N__56496;
    wire N__56493;
    wire N__56490;
    wire N__56487;
    wire N__56484;
    wire N__56483;
    wire N__56482;
    wire N__56481;
    wire N__56480;
    wire N__56479;
    wire N__56476;
    wire N__56471;
    wire N__56468;
    wire N__56465;
    wire N__56462;
    wire N__56461;
    wire N__56456;
    wire N__56453;
    wire N__56450;
    wire N__56445;
    wire N__56438;
    wire N__56435;
    wire N__56432;
    wire N__56427;
    wire N__56424;
    wire N__56421;
    wire N__56418;
    wire N__56415;
    wire N__56412;
    wire N__56411;
    wire N__56408;
    wire N__56407;
    wire N__56406;
    wire N__56403;
    wire N__56400;
    wire N__56397;
    wire N__56396;
    wire N__56393;
    wire N__56390;
    wire N__56387;
    wire N__56382;
    wire N__56373;
    wire N__56372;
    wire N__56371;
    wire N__56370;
    wire N__56369;
    wire N__56366;
    wire N__56361;
    wire N__56358;
    wire N__56355;
    wire N__56354;
    wire N__56351;
    wire N__56348;
    wire N__56345;
    wire N__56342;
    wire N__56339;
    wire N__56334;
    wire N__56325;
    wire N__56324;
    wire N__56323;
    wire N__56322;
    wire N__56317;
    wire N__56312;
    wire N__56309;
    wire N__56306;
    wire N__56303;
    wire N__56298;
    wire N__56295;
    wire N__56292;
    wire N__56289;
    wire N__56286;
    wire N__56283;
    wire N__56280;
    wire N__56277;
    wire N__56276;
    wire N__56273;
    wire N__56272;
    wire N__56269;
    wire N__56268;
    wire N__56265;
    wire N__56262;
    wire N__56259;
    wire N__56256;
    wire N__56247;
    wire N__56244;
    wire N__56241;
    wire N__56240;
    wire N__56239;
    wire N__56236;
    wire N__56233;
    wire N__56230;
    wire N__56227;
    wire N__56224;
    wire N__56223;
    wire N__56220;
    wire N__56217;
    wire N__56214;
    wire N__56211;
    wire N__56208;
    wire N__56203;
    wire N__56196;
    wire N__56193;
    wire N__56192;
    wire N__56189;
    wire N__56186;
    wire N__56185;
    wire N__56182;
    wire N__56179;
    wire N__56176;
    wire N__56171;
    wire N__56166;
    wire N__56163;
    wire N__56160;
    wire N__56159;
    wire N__56156;
    wire N__56153;
    wire N__56148;
    wire N__56147;
    wire N__56144;
    wire N__56143;
    wire N__56140;
    wire N__56139;
    wire N__56136;
    wire N__56133;
    wire N__56130;
    wire N__56127;
    wire N__56124;
    wire N__56119;
    wire N__56112;
    wire N__56109;
    wire N__56106;
    wire N__56103;
    wire N__56100;
    wire N__56097;
    wire N__56094;
    wire N__56091;
    wire N__56088;
    wire N__56085;
    wire N__56084;
    wire N__56079;
    wire N__56076;
    wire N__56073;
    wire N__56072;
    wire N__56069;
    wire N__56066;
    wire N__56063;
    wire N__56060;
    wire N__56057;
    wire N__56056;
    wire N__56051;
    wire N__56048;
    wire N__56043;
    wire N__56040;
    wire N__56039;
    wire N__56038;
    wire N__56035;
    wire N__56030;
    wire N__56027;
    wire N__56022;
    wire N__56019;
    wire N__56016;
    wire N__56013;
    wire N__56010;
    wire N__56009;
    wire N__56006;
    wire N__56005;
    wire N__56002;
    wire N__55999;
    wire N__55994;
    wire N__55991;
    wire N__55988;
    wire N__55983;
    wire N__55980;
    wire N__55977;
    wire N__55976;
    wire N__55973;
    wire N__55972;
    wire N__55969;
    wire N__55966;
    wire N__55965;
    wire N__55962;
    wire N__55959;
    wire N__55956;
    wire N__55953;
    wire N__55944;
    wire N__55943;
    wire N__55938;
    wire N__55935;
    wire N__55932;
    wire N__55931;
    wire N__55928;
    wire N__55923;
    wire N__55920;
    wire N__55919;
    wire N__55916;
    wire N__55913;
    wire N__55910;
    wire N__55905;
    wire N__55902;
    wire N__55901;
    wire N__55900;
    wire N__55899;
    wire N__55898;
    wire N__55889;
    wire N__55886;
    wire N__55883;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55873;
    wire N__55866;
    wire N__55863;
    wire N__55860;
    wire N__55857;
    wire N__55854;
    wire N__55851;
    wire N__55848;
    wire N__55845;
    wire N__55842;
    wire N__55839;
    wire N__55838;
    wire N__55835;
    wire N__55832;
    wire N__55827;
    wire N__55824;
    wire N__55823;
    wire N__55820;
    wire N__55817;
    wire N__55814;
    wire N__55811;
    wire N__55808;
    wire N__55803;
    wire N__55800;
    wire N__55799;
    wire N__55798;
    wire N__55797;
    wire N__55790;
    wire N__55787;
    wire N__55782;
    wire N__55779;
    wire N__55776;
    wire N__55775;
    wire N__55770;
    wire N__55767;
    wire N__55766;
    wire N__55761;
    wire N__55760;
    wire N__55757;
    wire N__55754;
    wire N__55751;
    wire N__55746;
    wire N__55743;
    wire N__55742;
    wire N__55741;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55731;
    wire N__55728;
    wire N__55727;
    wire N__55724;
    wire N__55721;
    wire N__55718;
    wire N__55715;
    wire N__55712;
    wire N__55709;
    wire N__55704;
    wire N__55701;
    wire N__55698;
    wire N__55695;
    wire N__55686;
    wire N__55683;
    wire N__55682;
    wire N__55679;
    wire N__55676;
    wire N__55673;
    wire N__55670;
    wire N__55665;
    wire N__55664;
    wire N__55661;
    wire N__55658;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55644;
    wire N__55641;
    wire N__55638;
    wire N__55635;
    wire N__55632;
    wire N__55631;
    wire N__55630;
    wire N__55627;
    wire N__55624;
    wire N__55621;
    wire N__55618;
    wire N__55615;
    wire N__55612;
    wire N__55611;
    wire N__55604;
    wire N__55601;
    wire N__55598;
    wire N__55593;
    wire N__55590;
    wire N__55587;
    wire N__55584;
    wire N__55581;
    wire N__55578;
    wire N__55575;
    wire N__55572;
    wire N__55569;
    wire N__55566;
    wire N__55565;
    wire N__55564;
    wire N__55561;
    wire N__55558;
    wire N__55555;
    wire N__55552;
    wire N__55549;
    wire N__55546;
    wire N__55543;
    wire N__55538;
    wire N__55533;
    wire N__55530;
    wire N__55527;
    wire N__55524;
    wire N__55523;
    wire N__55520;
    wire N__55517;
    wire N__55514;
    wire N__55513;
    wire N__55512;
    wire N__55509;
    wire N__55508;
    wire N__55505;
    wire N__55500;
    wire N__55497;
    wire N__55494;
    wire N__55489;
    wire N__55482;
    wire N__55479;
    wire N__55478;
    wire N__55475;
    wire N__55472;
    wire N__55469;
    wire N__55466;
    wire N__55463;
    wire N__55460;
    wire N__55455;
    wire N__55454;
    wire N__55451;
    wire N__55448;
    wire N__55445;
    wire N__55442;
    wire N__55439;
    wire N__55434;
    wire N__55431;
    wire N__55430;
    wire N__55429;
    wire N__55426;
    wire N__55423;
    wire N__55420;
    wire N__55415;
    wire N__55410;
    wire N__55407;
    wire N__55404;
    wire N__55401;
    wire N__55398;
    wire N__55395;
    wire N__55392;
    wire N__55389;
    wire N__55386;
    wire N__55383;
    wire N__55380;
    wire N__55377;
    wire N__55374;
    wire N__55371;
    wire N__55368;
    wire N__55365;
    wire N__55362;
    wire N__55359;
    wire N__55356;
    wire N__55353;
    wire N__55350;
    wire N__55347;
    wire N__55344;
    wire N__55341;
    wire N__55338;
    wire N__55335;
    wire N__55332;
    wire N__55331;
    wire N__55330;
    wire N__55329;
    wire N__55326;
    wire N__55323;
    wire N__55322;
    wire N__55319;
    wire N__55316;
    wire N__55311;
    wire N__55308;
    wire N__55305;
    wire N__55302;
    wire N__55297;
    wire N__55290;
    wire N__55287;
    wire N__55284;
    wire N__55281;
    wire N__55278;
    wire N__55275;
    wire N__55272;
    wire N__55269;
    wire N__55266;
    wire N__55263;
    wire N__55260;
    wire N__55257;
    wire N__55254;
    wire N__55251;
    wire N__55248;
    wire N__55245;
    wire N__55242;
    wire N__55241;
    wire N__55238;
    wire N__55235;
    wire N__55232;
    wire N__55229;
    wire N__55226;
    wire N__55221;
    wire N__55220;
    wire N__55217;
    wire N__55214;
    wire N__55211;
    wire N__55208;
    wire N__55207;
    wire N__55206;
    wire N__55203;
    wire N__55200;
    wire N__55195;
    wire N__55188;
    wire N__55187;
    wire N__55186;
    wire N__55185;
    wire N__55184;
    wire N__55179;
    wire N__55174;
    wire N__55171;
    wire N__55168;
    wire N__55165;
    wire N__55162;
    wire N__55157;
    wire N__55152;
    wire N__55149;
    wire N__55146;
    wire N__55143;
    wire N__55140;
    wire N__55137;
    wire N__55134;
    wire N__55133;
    wire N__55128;
    wire N__55125;
    wire N__55124;
    wire N__55121;
    wire N__55118;
    wire N__55115;
    wire N__55114;
    wire N__55113;
    wire N__55110;
    wire N__55107;
    wire N__55104;
    wire N__55101;
    wire N__55100;
    wire N__55097;
    wire N__55092;
    wire N__55087;
    wire N__55080;
    wire N__55077;
    wire N__55074;
    wire N__55071;
    wire N__55070;
    wire N__55069;
    wire N__55066;
    wire N__55063;
    wire N__55060;
    wire N__55057;
    wire N__55050;
    wire N__55049;
    wire N__55046;
    wire N__55045;
    wire N__55040;
    wire N__55037;
    wire N__55034;
    wire N__55031;
    wire N__55028;
    wire N__55023;
    wire N__55022;
    wire N__55021;
    wire N__55020;
    wire N__55017;
    wire N__55014;
    wire N__55009;
    wire N__55006;
    wire N__55003;
    wire N__55000;
    wire N__54995;
    wire N__54992;
    wire N__54987;
    wire N__54984;
    wire N__54981;
    wire N__54978;
    wire N__54975;
    wire N__54972;
    wire N__54969;
    wire N__54968;
    wire N__54963;
    wire N__54960;
    wire N__54957;
    wire N__54954;
    wire N__54951;
    wire N__54950;
    wire N__54947;
    wire N__54944;
    wire N__54943;
    wire N__54940;
    wire N__54937;
    wire N__54936;
    wire N__54933;
    wire N__54930;
    wire N__54927;
    wire N__54924;
    wire N__54921;
    wire N__54918;
    wire N__54909;
    wire N__54906;
    wire N__54903;
    wire N__54900;
    wire N__54897;
    wire N__54894;
    wire N__54891;
    wire N__54888;
    wire N__54885;
    wire N__54884;
    wire N__54883;
    wire N__54882;
    wire N__54881;
    wire N__54880;
    wire N__54879;
    wire N__54872;
    wire N__54863;
    wire N__54862;
    wire N__54861;
    wire N__54860;
    wire N__54859;
    wire N__54858;
    wire N__54857;
    wire N__54856;
    wire N__54855;
    wire N__54854;
    wire N__54853;
    wire N__54852;
    wire N__54851;
    wire N__54850;
    wire N__54849;
    wire N__54848;
    wire N__54847;
    wire N__54846;
    wire N__54845;
    wire N__54844;
    wire N__54843;
    wire N__54842;
    wire N__54841;
    wire N__54840;
    wire N__54839;
    wire N__54838;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54834;
    wire N__54833;
    wire N__54832;
    wire N__54831;
    wire N__54830;
    wire N__54829;
    wire N__54828;
    wire N__54827;
    wire N__54822;
    wire N__54815;
    wire N__54806;
    wire N__54799;
    wire N__54790;
    wire N__54783;
    wire N__54774;
    wire N__54767;
    wire N__54758;
    wire N__54755;
    wire N__54754;
    wire N__54751;
    wire N__54750;
    wire N__54747;
    wire N__54746;
    wire N__54743;
    wire N__54742;
    wire N__54741;
    wire N__54740;
    wire N__54739;
    wire N__54738;
    wire N__54737;
    wire N__54736;
    wire N__54733;
    wire N__54732;
    wire N__54729;
    wire N__54728;
    wire N__54725;
    wire N__54724;
    wire N__54721;
    wire N__54720;
    wire N__54719;
    wire N__54718;
    wire N__54717;
    wire N__54716;
    wire N__54715;
    wire N__54714;
    wire N__54695;
    wire N__54680;
    wire N__54673;
    wire N__54664;
    wire N__54649;
    wire N__54642;
    wire N__54633;
    wire N__54632;
    wire N__54631;
    wire N__54630;
    wire N__54615;
    wire N__54614;
    wire N__54613;
    wire N__54612;
    wire N__54611;
    wire N__54610;
    wire N__54609;
    wire N__54608;
    wire N__54607;
    wire N__54606;
    wire N__54605;
    wire N__54604;
    wire N__54603;
    wire N__54602;
    wire N__54601;
    wire N__54600;
    wire N__54599;
    wire N__54598;
    wire N__54597;
    wire N__54596;
    wire N__54595;
    wire N__54594;
    wire N__54593;
    wire N__54590;
    wire N__54589;
    wire N__54586;
    wire N__54585;
    wire N__54582;
    wire N__54581;
    wire N__54580;
    wire N__54579;
    wire N__54578;
    wire N__54577;
    wire N__54576;
    wire N__54575;
    wire N__54574;
    wire N__54573;
    wire N__54572;
    wire N__54571;
    wire N__54570;
    wire N__54569;
    wire N__54566;
    wire N__54559;
    wire N__54550;
    wire N__54543;
    wire N__54534;
    wire N__54527;
    wire N__54518;
    wire N__54517;
    wire N__54516;
    wire N__54515;
    wire N__54514;
    wire N__54513;
    wire N__54512;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54508;
    wire N__54507;
    wire N__54506;
    wire N__54505;
    wire N__54504;
    wire N__54503;
    wire N__54502;
    wire N__54501;
    wire N__54500;
    wire N__54499;
    wire N__54498;
    wire N__54497;
    wire N__54496;
    wire N__54495;
    wire N__54494;
    wire N__54493;
    wire N__54492;
    wire N__54491;
    wire N__54490;
    wire N__54475;
    wire N__54474;
    wire N__54471;
    wire N__54470;
    wire N__54467;
    wire N__54466;
    wire N__54463;
    wire N__54462;
    wire N__54461;
    wire N__54458;
    wire N__54457;
    wire N__54454;
    wire N__54453;
    wire N__54450;
    wire N__54449;
    wire N__54448;
    wire N__54445;
    wire N__54444;
    wire N__54441;
    wire N__54440;
    wire N__54437;
    wire N__54436;
    wire N__54435;
    wire N__54432;
    wire N__54431;
    wire N__54428;
    wire N__54427;
    wire N__54424;
    wire N__54423;
    wire N__54422;
    wire N__54421;
    wire N__54420;
    wire N__54419;
    wire N__54418;
    wire N__54417;
    wire N__54402;
    wire N__54395;
    wire N__54386;
    wire N__54379;
    wire N__54370;
    wire N__54363;
    wire N__54354;
    wire N__54347;
    wire N__54338;
    wire N__54337;
    wire N__54336;
    wire N__54335;
    wire N__54334;
    wire N__54333;
    wire N__54332;
    wire N__54331;
    wire N__54330;
    wire N__54329;
    wire N__54328;
    wire N__54327;
    wire N__54326;
    wire N__54325;
    wire N__54324;
    wire N__54323;
    wire N__54322;
    wire N__54321;
    wire N__54320;
    wire N__54319;
    wire N__54318;
    wire N__54317;
    wire N__54316;
    wire N__54315;
    wire N__54314;
    wire N__54313;
    wire N__54312;
    wire N__54311;
    wire N__54310;
    wire N__54309;
    wire N__54308;
    wire N__54307;
    wire N__54304;
    wire N__54289;
    wire N__54274;
    wire N__54259;
    wire N__54244;
    wire N__54243;
    wire N__54240;
    wire N__54239;
    wire N__54236;
    wire N__54235;
    wire N__54232;
    wire N__54231;
    wire N__54230;
    wire N__54227;
    wire N__54226;
    wire N__54223;
    wire N__54222;
    wire N__54219;
    wire N__54218;
    wire N__54199;
    wire N__54192;
    wire N__54183;
    wire N__54176;
    wire N__54167;
    wire N__54160;
    wire N__54151;
    wire N__54150;
    wire N__54147;
    wire N__54146;
    wire N__54143;
    wire N__54142;
    wire N__54139;
    wire N__54138;
    wire N__54137;
    wire N__54136;
    wire N__54135;
    wire N__54134;
    wire N__54133;
    wire N__54132;
    wire N__54131;
    wire N__54124;
    wire N__54115;
    wire N__54106;
    wire N__54103;
    wire N__54088;
    wire N__54073;
    wire N__54058;
    wire N__54043;
    wire N__54036;
    wire N__54027;
    wire N__54026;
    wire N__54025;
    wire N__54024;
    wire N__54023;
    wire N__54022;
    wire N__54021;
    wire N__54020;
    wire N__54015;
    wire N__54002;
    wire N__54001;
    wire N__54000;
    wire N__53999;
    wire N__53998;
    wire N__53997;
    wire N__53996;
    wire N__53995;
    wire N__53990;
    wire N__53983;
    wire N__53974;
    wire N__53971;
    wire N__53968;
    wire N__53961;
    wire N__53952;
    wire N__53949;
    wire N__53944;
    wire N__53941;
    wire N__53934;
    wire N__53929;
    wire N__53924;
    wire N__53919;
    wire N__53916;
    wire N__53915;
    wire N__53912;
    wire N__53911;
    wire N__53910;
    wire N__53909;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53895;
    wire N__53894;
    wire N__53891;
    wire N__53888;
    wire N__53885;
    wire N__53882;
    wire N__53881;
    wire N__53878;
    wire N__53877;
    wire N__53874;
    wire N__53871;
    wire N__53866;
    wire N__53863;
    wire N__53860;
    wire N__53857;
    wire N__53854;
    wire N__53851;
    wire N__53848;
    wire N__53843;
    wire N__53838;
    wire N__53835;
    wire N__53832;
    wire N__53823;
    wire N__53820;
    wire N__53817;
    wire N__53814;
    wire N__53811;
    wire N__53808;
    wire N__53807;
    wire N__53804;
    wire N__53803;
    wire N__53802;
    wire N__53799;
    wire N__53796;
    wire N__53793;
    wire N__53790;
    wire N__53787;
    wire N__53782;
    wire N__53779;
    wire N__53776;
    wire N__53769;
    wire N__53768;
    wire N__53767;
    wire N__53766;
    wire N__53765;
    wire N__53764;
    wire N__53761;
    wire N__53760;
    wire N__53759;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53749;
    wire N__53748;
    wire N__53747;
    wire N__53746;
    wire N__53745;
    wire N__53744;
    wire N__53743;
    wire N__53742;
    wire N__53741;
    wire N__53740;
    wire N__53737;
    wire N__53734;
    wire N__53731;
    wire N__53728;
    wire N__53725;
    wire N__53724;
    wire N__53717;
    wire N__53714;
    wire N__53713;
    wire N__53712;
    wire N__53709;
    wire N__53706;
    wire N__53703;
    wire N__53700;
    wire N__53699;
    wire N__53698;
    wire N__53697;
    wire N__53696;
    wire N__53695;
    wire N__53694;
    wire N__53693;
    wire N__53692;
    wire N__53689;
    wire N__53686;
    wire N__53683;
    wire N__53680;
    wire N__53677;
    wire N__53666;
    wire N__53665;
    wire N__53662;
    wire N__53657;
    wire N__53654;
    wire N__53651;
    wire N__53642;
    wire N__53641;
    wire N__53640;
    wire N__53637;
    wire N__53634;
    wire N__53631;
    wire N__53628;
    wire N__53625;
    wire N__53622;
    wire N__53619;
    wire N__53616;
    wire N__53603;
    wire N__53600;
    wire N__53589;
    wire N__53586;
    wire N__53583;
    wire N__53580;
    wire N__53563;
    wire N__53558;
    wire N__53547;
    wire N__53544;
    wire N__53543;
    wire N__53542;
    wire N__53539;
    wire N__53536;
    wire N__53533;
    wire N__53530;
    wire N__53523;
    wire N__53520;
    wire N__53517;
    wire N__53514;
    wire N__53511;
    wire N__53510;
    wire N__53509;
    wire N__53506;
    wire N__53503;
    wire N__53500;
    wire N__53497;
    wire N__53490;
    wire N__53487;
    wire N__53484;
    wire N__53481;
    wire N__53480;
    wire N__53479;
    wire N__53476;
    wire N__53473;
    wire N__53470;
    wire N__53467;
    wire N__53460;
    wire N__53457;
    wire N__53454;
    wire N__53451;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53441;
    wire N__53440;
    wire N__53437;
    wire N__53434;
    wire N__53431;
    wire N__53428;
    wire N__53421;
    wire N__53418;
    wire N__53415;
    wire N__53412;
    wire N__53409;
    wire N__53408;
    wire N__53405;
    wire N__53404;
    wire N__53401;
    wire N__53398;
    wire N__53395;
    wire N__53390;
    wire N__53385;
    wire N__53382;
    wire N__53379;
    wire N__53376;
    wire N__53375;
    wire N__53374;
    wire N__53371;
    wire N__53368;
    wire N__53365;
    wire N__53362;
    wire N__53355;
    wire N__53352;
    wire N__53349;
    wire N__53346;
    wire N__53343;
    wire N__53342;
    wire N__53341;
    wire N__53338;
    wire N__53335;
    wire N__53332;
    wire N__53325;
    wire N__53322;
    wire N__53319;
    wire N__53316;
    wire N__53313;
    wire N__53310;
    wire N__53309;
    wire N__53306;
    wire N__53303;
    wire N__53302;
    wire N__53299;
    wire N__53296;
    wire N__53293;
    wire N__53290;
    wire N__53283;
    wire N__53280;
    wire N__53277;
    wire N__53274;
    wire N__53271;
    wire N__53270;
    wire N__53267;
    wire N__53264;
    wire N__53263;
    wire N__53258;
    wire N__53255;
    wire N__53252;
    wire N__53247;
    wire N__53244;
    wire N__53241;
    wire N__53238;
    wire N__53235;
    wire N__53232;
    wire N__53229;
    wire N__53226;
    wire N__53223;
    wire N__53220;
    wire N__53219;
    wire N__53216;
    wire N__53213;
    wire N__53212;
    wire N__53207;
    wire N__53204;
    wire N__53201;
    wire N__53196;
    wire N__53193;
    wire N__53190;
    wire N__53187;
    wire N__53184;
    wire N__53181;
    wire N__53180;
    wire N__53177;
    wire N__53174;
    wire N__53171;
    wire N__53170;
    wire N__53165;
    wire N__53162;
    wire N__53159;
    wire N__53154;
    wire N__53151;
    wire N__53148;
    wire N__53145;
    wire N__53142;
    wire N__53139;
    wire N__53136;
    wire N__53133;
    wire N__53132;
    wire N__53129;
    wire N__53126;
    wire N__53125;
    wire N__53120;
    wire N__53117;
    wire N__53114;
    wire N__53109;
    wire N__53106;
    wire N__53103;
    wire N__53100;
    wire N__53099;
    wire N__53096;
    wire N__53093;
    wire N__53090;
    wire N__53089;
    wire N__53084;
    wire N__53081;
    wire N__53078;
    wire N__53073;
    wire N__53070;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53054;
    wire N__53051;
    wire N__53048;
    wire N__53045;
    wire N__53042;
    wire N__53039;
    wire N__53038;
    wire N__53033;
    wire N__53030;
    wire N__53027;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53013;
    wire N__53010;
    wire N__53007;
    wire N__53006;
    wire N__53003;
    wire N__53000;
    wire N__52997;
    wire N__52996;
    wire N__52993;
    wire N__52990;
    wire N__52987;
    wire N__52982;
    wire N__52977;
    wire N__52974;
    wire N__52971;
    wire N__52968;
    wire N__52965;
    wire N__52962;
    wire N__52959;
    wire N__52956;
    wire N__52955;
    wire N__52952;
    wire N__52949;
    wire N__52946;
    wire N__52943;
    wire N__52942;
    wire N__52939;
    wire N__52936;
    wire N__52933;
    wire N__52930;
    wire N__52923;
    wire N__52920;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52908;
    wire N__52905;
    wire N__52904;
    wire N__52901;
    wire N__52898;
    wire N__52895;
    wire N__52892;
    wire N__52891;
    wire N__52886;
    wire N__52883;
    wire N__52880;
    wire N__52875;
    wire N__52872;
    wire N__52869;
    wire N__52866;
    wire N__52863;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52851;
    wire N__52848;
    wire N__52845;
    wire N__52842;
    wire N__52839;
    wire N__52836;
    wire N__52835;
    wire N__52832;
    wire N__52829;
    wire N__52826;
    wire N__52823;
    wire N__52820;
    wire N__52817;
    wire N__52816;
    wire N__52811;
    wire N__52808;
    wire N__52805;
    wire N__52800;
    wire N__52797;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52776;
    wire N__52773;
    wire N__52770;
    wire N__52769;
    wire N__52766;
    wire N__52763;
    wire N__52760;
    wire N__52757;
    wire N__52756;
    wire N__52751;
    wire N__52748;
    wire N__52745;
    wire N__52740;
    wire N__52737;
    wire N__52734;
    wire N__52731;
    wire N__52728;
    wire N__52725;
    wire N__52722;
    wire N__52721;
    wire N__52716;
    wire N__52713;
    wire N__52712;
    wire N__52709;
    wire N__52706;
    wire N__52703;
    wire N__52698;
    wire N__52695;
    wire N__52694;
    wire N__52691;
    wire N__52688;
    wire N__52685;
    wire N__52682;
    wire N__52679;
    wire N__52676;
    wire N__52673;
    wire N__52670;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52653;
    wire N__52650;
    wire N__52647;
    wire N__52644;
    wire N__52641;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52628;
    wire N__52625;
    wire N__52622;
    wire N__52619;
    wire N__52616;
    wire N__52615;
    wire N__52610;
    wire N__52607;
    wire N__52604;
    wire N__52599;
    wire N__52596;
    wire N__52593;
    wire N__52590;
    wire N__52587;
    wire N__52584;
    wire N__52581;
    wire N__52578;
    wire N__52575;
    wire N__52572;
    wire N__52569;
    wire N__52568;
    wire N__52565;
    wire N__52562;
    wire N__52561;
    wire N__52556;
    wire N__52553;
    wire N__52552;
    wire N__52549;
    wire N__52546;
    wire N__52543;
    wire N__52540;
    wire N__52537;
    wire N__52534;
    wire N__52531;
    wire N__52526;
    wire N__52525;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52500;
    wire N__52497;
    wire N__52494;
    wire N__52491;
    wire N__52488;
    wire N__52485;
    wire N__52482;
    wire N__52481;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52455;
    wire N__52454;
    wire N__52451;
    wire N__52446;
    wire N__52443;
    wire N__52440;
    wire N__52437;
    wire N__52434;
    wire N__52425;
    wire N__52422;
    wire N__52419;
    wire N__52416;
    wire N__52413;
    wire N__52410;
    wire N__52409;
    wire N__52408;
    wire N__52407;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52392;
    wire N__52389;
    wire N__52384;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52374;
    wire N__52371;
    wire N__52366;
    wire N__52363;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52353;
    wire N__52350;
    wire N__52347;
    wire N__52344;
    wire N__52335;
    wire N__52332;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52317;
    wire N__52314;
    wire N__52311;
    wire N__52308;
    wire N__52305;
    wire N__52302;
    wire N__52299;
    wire N__52296;
    wire N__52293;
    wire N__52290;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52278;
    wire N__52275;
    wire N__52272;
    wire N__52269;
    wire N__52266;
    wire N__52263;
    wire N__52260;
    wire N__52257;
    wire N__52254;
    wire N__52251;
    wire N__52248;
    wire N__52245;
    wire N__52242;
    wire N__52241;
    wire N__52238;
    wire N__52235;
    wire N__52232;
    wire N__52229;
    wire N__52226;
    wire N__52223;
    wire N__52220;
    wire N__52215;
    wire N__52212;
    wire N__52209;
    wire N__52206;
    wire N__52205;
    wire N__52204;
    wire N__52201;
    wire N__52198;
    wire N__52195;
    wire N__52192;
    wire N__52191;
    wire N__52188;
    wire N__52185;
    wire N__52182;
    wire N__52179;
    wire N__52176;
    wire N__52167;
    wire N__52166;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52155;
    wire N__52150;
    wire N__52145;
    wire N__52140;
    wire N__52137;
    wire N__52134;
    wire N__52133;
    wire N__52132;
    wire N__52129;
    wire N__52124;
    wire N__52121;
    wire N__52118;
    wire N__52113;
    wire N__52110;
    wire N__52107;
    wire N__52104;
    wire N__52101;
    wire N__52098;
    wire N__52097;
    wire N__52094;
    wire N__52091;
    wire N__52090;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52072;
    wire N__52071;
    wire N__52068;
    wire N__52065;
    wire N__52062;
    wire N__52059;
    wire N__52056;
    wire N__52051;
    wire N__52048;
    wire N__52045;
    wire N__52042;
    wire N__52035;
    wire N__52032;
    wire N__52029;
    wire N__52028;
    wire N__52025;
    wire N__52022;
    wire N__52017;
    wire N__52014;
    wire N__52013;
    wire N__52010;
    wire N__52007;
    wire N__52004;
    wire N__51999;
    wire N__51998;
    wire N__51995;
    wire N__51992;
    wire N__51987;
    wire N__51984;
    wire N__51981;
    wire N__51978;
    wire N__51975;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51960;
    wire N__51957;
    wire N__51954;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51944;
    wire N__51943;
    wire N__51940;
    wire N__51937;
    wire N__51934;
    wire N__51931;
    wire N__51924;
    wire N__51921;
    wire N__51918;
    wire N__51915;
    wire N__51912;
    wire N__51909;
    wire N__51906;
    wire N__51903;
    wire N__51900;
    wire N__51897;
    wire N__51894;
    wire N__51891;
    wire N__51888;
    wire N__51887;
    wire N__51882;
    wire N__51881;
    wire N__51878;
    wire N__51875;
    wire N__51870;
    wire N__51867;
    wire N__51864;
    wire N__51861;
    wire N__51858;
    wire N__51855;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51843;
    wire N__51840;
    wire N__51837;
    wire N__51834;
    wire N__51833;
    wire N__51828;
    wire N__51825;
    wire N__51822;
    wire N__51819;
    wire N__51816;
    wire N__51813;
    wire N__51810;
    wire N__51809;
    wire N__51804;
    wire N__51801;
    wire N__51800;
    wire N__51797;
    wire N__51794;
    wire N__51791;
    wire N__51788;
    wire N__51785;
    wire N__51780;
    wire N__51779;
    wire N__51778;
    wire N__51777;
    wire N__51774;
    wire N__51773;
    wire N__51770;
    wire N__51767;
    wire N__51764;
    wire N__51761;
    wire N__51758;
    wire N__51751;
    wire N__51748;
    wire N__51741;
    wire N__51738;
    wire N__51735;
    wire N__51732;
    wire N__51729;
    wire N__51728;
    wire N__51727;
    wire N__51724;
    wire N__51719;
    wire N__51714;
    wire N__51711;
    wire N__51708;
    wire N__51705;
    wire N__51702;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51687;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51672;
    wire N__51671;
    wire N__51668;
    wire N__51665;
    wire N__51662;
    wire N__51657;
    wire N__51654;
    wire N__51651;
    wire N__51648;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51627;
    wire N__51626;
    wire N__51623;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51597;
    wire N__51594;
    wire N__51591;
    wire N__51588;
    wire N__51585;
    wire N__51582;
    wire N__51581;
    wire N__51578;
    wire N__51575;
    wire N__51574;
    wire N__51573;
    wire N__51568;
    wire N__51565;
    wire N__51564;
    wire N__51563;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51531;
    wire N__51528;
    wire N__51525;
    wire N__51522;
    wire N__51521;
    wire N__51518;
    wire N__51517;
    wire N__51510;
    wire N__51507;
    wire N__51504;
    wire N__51501;
    wire N__51498;
    wire N__51495;
    wire N__51492;
    wire N__51489;
    wire N__51486;
    wire N__51483;
    wire N__51480;
    wire N__51477;
    wire N__51474;
    wire N__51471;
    wire N__51468;
    wire N__51467;
    wire N__51466;
    wire N__51465;
    wire N__51464;
    wire N__51461;
    wire N__51460;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51448;
    wire N__51447;
    wire N__51446;
    wire N__51443;
    wire N__51440;
    wire N__51439;
    wire N__51436;
    wire N__51433;
    wire N__51428;
    wire N__51425;
    wire N__51424;
    wire N__51421;
    wire N__51420;
    wire N__51419;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51402;
    wire N__51397;
    wire N__51390;
    wire N__51387;
    wire N__51372;
    wire N__51369;
    wire N__51366;
    wire N__51363;
    wire N__51360;
    wire N__51357;
    wire N__51354;
    wire N__51351;
    wire N__51348;
    wire N__51345;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51328;
    wire N__51323;
    wire N__51320;
    wire N__51317;
    wire N__51312;
    wire N__51309;
    wire N__51306;
    wire N__51303;
    wire N__51300;
    wire N__51297;
    wire N__51294;
    wire N__51291;
    wire N__51288;
    wire N__51285;
    wire N__51282;
    wire N__51279;
    wire N__51276;
    wire N__51275;
    wire N__51272;
    wire N__51269;
    wire N__51264;
    wire N__51261;
    wire N__51258;
    wire N__51255;
    wire N__51252;
    wire N__51249;
    wire N__51246;
    wire N__51243;
    wire N__51240;
    wire N__51237;
    wire N__51234;
    wire N__51233;
    wire N__51232;
    wire N__51229;
    wire N__51224;
    wire N__51223;
    wire N__51220;
    wire N__51219;
    wire N__51218;
    wire N__51217;
    wire N__51216;
    wire N__51213;
    wire N__51212;
    wire N__51211;
    wire N__51208;
    wire N__51207;
    wire N__51206;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51192;
    wire N__51189;
    wire N__51184;
    wire N__51181;
    wire N__51176;
    wire N__51159;
    wire N__51156;
    wire N__51153;
    wire N__51150;
    wire N__51149;
    wire N__51144;
    wire N__51141;
    wire N__51138;
    wire N__51137;
    wire N__51136;
    wire N__51131;
    wire N__51128;
    wire N__51125;
    wire N__51120;
    wire N__51117;
    wire N__51114;
    wire N__51111;
    wire N__51108;
    wire N__51105;
    wire N__51102;
    wire N__51099;
    wire N__51096;
    wire N__51093;
    wire N__51092;
    wire N__51089;
    wire N__51086;
    wire N__51085;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51069;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51044;
    wire N__51041;
    wire N__51038;
    wire N__51035;
    wire N__51030;
    wire N__51029;
    wire N__51024;
    wire N__51021;
    wire N__51018;
    wire N__51015;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51003;
    wire N__51000;
    wire N__50997;
    wire N__50994;
    wire N__50991;
    wire N__50988;
    wire N__50985;
    wire N__50984;
    wire N__50979;
    wire N__50976;
    wire N__50973;
    wire N__50972;
    wire N__50971;
    wire N__50970;
    wire N__50969;
    wire N__50966;
    wire N__50961;
    wire N__50956;
    wire N__50949;
    wire N__50946;
    wire N__50945;
    wire N__50944;
    wire N__50943;
    wire N__50942;
    wire N__50941;
    wire N__50940;
    wire N__50937;
    wire N__50932;
    wire N__50927;
    wire N__50922;
    wire N__50913;
    wire N__50912;
    wire N__50911;
    wire N__50910;
    wire N__50909;
    wire N__50908;
    wire N__50905;
    wire N__50904;
    wire N__50901;
    wire N__50898;
    wire N__50895;
    wire N__50892;
    wire N__50889;
    wire N__50886;
    wire N__50883;
    wire N__50880;
    wire N__50877;
    wire N__50874;
    wire N__50871;
    wire N__50868;
    wire N__50867;
    wire N__50866;
    wire N__50865;
    wire N__50864;
    wire N__50861;
    wire N__50858;
    wire N__50851;
    wire N__50848;
    wire N__50845;
    wire N__50842;
    wire N__50837;
    wire N__50834;
    wire N__50829;
    wire N__50826;
    wire N__50825;
    wire N__50822;
    wire N__50817;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50805;
    wire N__50802;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50782;
    wire N__50779;
    wire N__50776;
    wire N__50773;
    wire N__50770;
    wire N__50767;
    wire N__50760;
    wire N__50757;
    wire N__50754;
    wire N__50751;
    wire N__50748;
    wire N__50745;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50726;
    wire N__50723;
    wire N__50720;
    wire N__50719;
    wire N__50718;
    wire N__50715;
    wire N__50712;
    wire N__50709;
    wire N__50706;
    wire N__50703;
    wire N__50698;
    wire N__50695;
    wire N__50692;
    wire N__50689;
    wire N__50686;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50670;
    wire N__50667;
    wire N__50664;
    wire N__50661;
    wire N__50658;
    wire N__50655;
    wire N__50652;
    wire N__50651;
    wire N__50650;
    wire N__50647;
    wire N__50644;
    wire N__50641;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50622;
    wire N__50621;
    wire N__50620;
    wire N__50617;
    wire N__50614;
    wire N__50611;
    wire N__50606;
    wire N__50601;
    wire N__50598;
    wire N__50595;
    wire N__50592;
    wire N__50589;
    wire N__50588;
    wire N__50585;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50575;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50556;
    wire N__50553;
    wire N__50550;
    wire N__50541;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50529;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50523;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50480;
    wire N__50477;
    wire N__50474;
    wire N__50473;
    wire N__50472;
    wire N__50467;
    wire N__50466;
    wire N__50465;
    wire N__50464;
    wire N__50463;
    wire N__50462;
    wire N__50461;
    wire N__50460;
    wire N__50459;
    wire N__50458;
    wire N__50455;
    wire N__50454;
    wire N__50453;
    wire N__50448;
    wire N__50445;
    wire N__50442;
    wire N__50439;
    wire N__50438;
    wire N__50437;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50429;
    wire N__50428;
    wire N__50427;
    wire N__50426;
    wire N__50425;
    wire N__50424;
    wire N__50423;
    wire N__50420;
    wire N__50417;
    wire N__50410;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50398;
    wire N__50395;
    wire N__50392;
    wire N__50391;
    wire N__50386;
    wire N__50381;
    wire N__50378;
    wire N__50375;
    wire N__50372;
    wire N__50369;
    wire N__50362;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50348;
    wire N__50339;
    wire N__50334;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50306;
    wire N__50301;
    wire N__50286;
    wire N__50283;
    wire N__50278;
    wire N__50273;
    wire N__50268;
    wire N__50261;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50241;
    wire N__50236;
    wire N__50235;
    wire N__50234;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50217;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50198;
    wire N__50195;
    wire N__50192;
    wire N__50189;
    wire N__50184;
    wire N__50183;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50177;
    wire N__50174;
    wire N__50169;
    wire N__50166;
    wire N__50163;
    wire N__50162;
    wire N__50161;
    wire N__50158;
    wire N__50157;
    wire N__50154;
    wire N__50153;
    wire N__50150;
    wire N__50147;
    wire N__50144;
    wire N__50141;
    wire N__50138;
    wire N__50135;
    wire N__50132;
    wire N__50129;
    wire N__50126;
    wire N__50123;
    wire N__50120;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50103;
    wire N__50100;
    wire N__50095;
    wire N__50090;
    wire N__50087;
    wire N__50084;
    wire N__50079;
    wire N__50076;
    wire N__50071;
    wire N__50066;
    wire N__50055;
    wire N__50052;
    wire N__50049;
    wire N__50048;
    wire N__50045;
    wire N__50044;
    wire N__50043;
    wire N__50042;
    wire N__50039;
    wire N__50036;
    wire N__50035;
    wire N__50034;
    wire N__50031;
    wire N__50026;
    wire N__50025;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50007;
    wire N__50004;
    wire N__50001;
    wire N__50000;
    wire N__49997;
    wire N__49992;
    wire N__49985;
    wire N__49982;
    wire N__49979;
    wire N__49974;
    wire N__49971;
    wire N__49962;
    wire N__49959;
    wire N__49958;
    wire N__49957;
    wire N__49956;
    wire N__49953;
    wire N__49948;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49940;
    wire N__49935;
    wire N__49932;
    wire N__49929;
    wire N__49924;
    wire N__49921;
    wire N__49918;
    wire N__49915;
    wire N__49910;
    wire N__49907;
    wire N__49904;
    wire N__49901;
    wire N__49896;
    wire N__49893;
    wire N__49886;
    wire N__49881;
    wire N__49878;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49866;
    wire N__49863;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49844;
    wire N__49841;
    wire N__49838;
    wire N__49833;
    wire N__49830;
    wire N__49829;
    wire N__49828;
    wire N__49827;
    wire N__49824;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49806;
    wire N__49799;
    wire N__49794;
    wire N__49793;
    wire N__49788;
    wire N__49787;
    wire N__49786;
    wire N__49783;
    wire N__49780;
    wire N__49777;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49765;
    wire N__49762;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49734;
    wire N__49731;
    wire N__49730;
    wire N__49727;
    wire N__49724;
    wire N__49723;
    wire N__49722;
    wire N__49719;
    wire N__49718;
    wire N__49713;
    wire N__49710;
    wire N__49707;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49693;
    wire N__49686;
    wire N__49685;
    wire N__49684;
    wire N__49681;
    wire N__49678;
    wire N__49675;
    wire N__49672;
    wire N__49669;
    wire N__49662;
    wire N__49659;
    wire N__49658;
    wire N__49657;
    wire N__49656;
    wire N__49653;
    wire N__49650;
    wire N__49649;
    wire N__49648;
    wire N__49645;
    wire N__49642;
    wire N__49639;
    wire N__49638;
    wire N__49635;
    wire N__49634;
    wire N__49629;
    wire N__49626;
    wire N__49623;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49611;
    wire N__49608;
    wire N__49603;
    wire N__49600;
    wire N__49597;
    wire N__49592;
    wire N__49589;
    wire N__49586;
    wire N__49583;
    wire N__49572;
    wire N__49569;
    wire N__49566;
    wire N__49563;
    wire N__49560;
    wire N__49557;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49536;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49523;
    wire N__49520;
    wire N__49517;
    wire N__49512;
    wire N__49509;
    wire N__49508;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49479;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49458;
    wire N__49455;
    wire N__49452;
    wire N__49449;
    wire N__49446;
    wire N__49445;
    wire N__49442;
    wire N__49439;
    wire N__49434;
    wire N__49431;
    wire N__49428;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49402;
    wire N__49397;
    wire N__49394;
    wire N__49389;
    wire N__49386;
    wire N__49385;
    wire N__49382;
    wire N__49379;
    wire N__49378;
    wire N__49373;
    wire N__49370;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49353;
    wire N__49350;
    wire N__49349;
    wire N__49344;
    wire N__49341;
    wire N__49338;
    wire N__49335;
    wire N__49332;
    wire N__49329;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49310;
    wire N__49307;
    wire N__49304;
    wire N__49303;
    wire N__49302;
    wire N__49299;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49287;
    wire N__49284;
    wire N__49281;
    wire N__49272;
    wire N__49269;
    wire N__49268;
    wire N__49265;
    wire N__49264;
    wire N__49261;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49249;
    wire N__49242;
    wire N__49239;
    wire N__49238;
    wire N__49237;
    wire N__49234;
    wire N__49231;
    wire N__49228;
    wire N__49225;
    wire N__49222;
    wire N__49215;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49196;
    wire N__49193;
    wire N__49190;
    wire N__49187;
    wire N__49186;
    wire N__49181;
    wire N__49178;
    wire N__49175;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49139;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49107;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49083;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49073;
    wire N__49070;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49054;
    wire N__49047;
    wire N__49044;
    wire N__49043;
    wire N__49040;
    wire N__49037;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49019;
    wire N__49014;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__49003;
    wire N__49000;
    wire N__48999;
    wire N__48996;
    wire N__48993;
    wire N__48992;
    wire N__48991;
    wire N__48990;
    wire N__48989;
    wire N__48988;
    wire N__48987;
    wire N__48986;
    wire N__48985;
    wire N__48984;
    wire N__48981;
    wire N__48980;
    wire N__48979;
    wire N__48978;
    wire N__48975;
    wire N__48970;
    wire N__48969;
    wire N__48966;
    wire N__48963;
    wire N__48962;
    wire N__48961;
    wire N__48960;
    wire N__48957;
    wire N__48954;
    wire N__48951;
    wire N__48948;
    wire N__48945;
    wire N__48942;
    wire N__48941;
    wire N__48938;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48928;
    wire N__48925;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48911;
    wire N__48908;
    wire N__48905;
    wire N__48902;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48882;
    wire N__48879;
    wire N__48874;
    wire N__48871;
    wire N__48870;
    wire N__48867;
    wire N__48860;
    wire N__48853;
    wire N__48850;
    wire N__48845;
    wire N__48842;
    wire N__48839;
    wire N__48838;
    wire N__48837;
    wire N__48834;
    wire N__48829;
    wire N__48826;
    wire N__48825;
    wire N__48824;
    wire N__48821;
    wire N__48814;
    wire N__48811;
    wire N__48806;
    wire N__48803;
    wire N__48800;
    wire N__48793;
    wire N__48790;
    wire N__48787;
    wire N__48768;
    wire N__48767;
    wire N__48766;
    wire N__48763;
    wire N__48758;
    wire N__48753;
    wire N__48750;
    wire N__48747;
    wire N__48744;
    wire N__48743;
    wire N__48740;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48732;
    wire N__48731;
    wire N__48728;
    wire N__48723;
    wire N__48718;
    wire N__48711;
    wire N__48710;
    wire N__48707;
    wire N__48704;
    wire N__48701;
    wire N__48698;
    wire N__48697;
    wire N__48692;
    wire N__48689;
    wire N__48684;
    wire N__48681;
    wire N__48680;
    wire N__48679;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48648;
    wire N__48645;
    wire N__48636;
    wire N__48633;
    wire N__48632;
    wire N__48629;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48606;
    wire N__48603;
    wire N__48600;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48585;
    wire N__48582;
    wire N__48579;
    wire N__48576;
    wire N__48573;
    wire N__48570;
    wire N__48567;
    wire N__48564;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48554;
    wire N__48549;
    wire N__48546;
    wire N__48543;
    wire N__48542;
    wire N__48537;
    wire N__48534;
    wire N__48531;
    wire N__48528;
    wire N__48525;
    wire N__48522;
    wire N__48519;
    wire N__48516;
    wire N__48515;
    wire N__48512;
    wire N__48511;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48496;
    wire N__48493;
    wire N__48486;
    wire N__48483;
    wire N__48482;
    wire N__48479;
    wire N__48476;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48450;
    wire N__48447;
    wire N__48444;
    wire N__48443;
    wire N__48440;
    wire N__48437;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48417;
    wire N__48416;
    wire N__48413;
    wire N__48412;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48390;
    wire N__48387;
    wire N__48384;
    wire N__48381;
    wire N__48380;
    wire N__48379;
    wire N__48378;
    wire N__48377;
    wire N__48376;
    wire N__48375;
    wire N__48374;
    wire N__48373;
    wire N__48372;
    wire N__48369;
    wire N__48366;
    wire N__48365;
    wire N__48364;
    wire N__48363;
    wire N__48362;
    wire N__48359;
    wire N__48356;
    wire N__48353;
    wire N__48350;
    wire N__48349;
    wire N__48348;
    wire N__48347;
    wire N__48346;
    wire N__48345;
    wire N__48338;
    wire N__48335;
    wire N__48330;
    wire N__48325;
    wire N__48324;
    wire N__48323;
    wire N__48322;
    wire N__48321;
    wire N__48320;
    wire N__48319;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48305;
    wire N__48302;
    wire N__48295;
    wire N__48294;
    wire N__48293;
    wire N__48288;
    wire N__48283;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48271;
    wire N__48270;
    wire N__48269;
    wire N__48260;
    wire N__48257;
    wire N__48256;
    wire N__48255;
    wire N__48254;
    wire N__48253;
    wire N__48252;
    wire N__48251;
    wire N__48250;
    wire N__48249;
    wire N__48248;
    wire N__48247;
    wire N__48246;
    wire N__48245;
    wire N__48244;
    wire N__48243;
    wire N__48242;
    wire N__48241;
    wire N__48240;
    wire N__48239;
    wire N__48238;
    wire N__48227;
    wire N__48222;
    wire N__48215;
    wire N__48210;
    wire N__48209;
    wire N__48208;
    wire N__48207;
    wire N__48206;
    wire N__48205;
    wire N__48204;
    wire N__48203;
    wire N__48202;
    wire N__48201;
    wire N__48200;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48169;
    wire N__48162;
    wire N__48159;
    wire N__48154;
    wire N__48143;
    wire N__48142;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48134;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48126;
    wire N__48117;
    wire N__48108;
    wire N__48099;
    wire N__48094;
    wire N__48091;
    wire N__48088;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48078;
    wire N__48077;
    wire N__48072;
    wire N__48069;
    wire N__48068;
    wire N__48067;
    wire N__48064;
    wire N__48047;
    wire N__48036;
    wire N__48029;
    wire N__48024;
    wire N__48013;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47995;
    wire N__47994;
    wire N__47991;
    wire N__47988;
    wire N__47983;
    wire N__47974;
    wire N__47969;
    wire N__47964;
    wire N__47961;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47947;
    wire N__47944;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47927;
    wire N__47922;
    wire N__47919;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47893;
    wire N__47890;
    wire N__47887;
    wire N__47884;
    wire N__47883;
    wire N__47880;
    wire N__47879;
    wire N__47878;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47862;
    wire N__47859;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47824;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47814;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47791;
    wire N__47790;
    wire N__47789;
    wire N__47788;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47770;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47752;
    wire N__47739;
    wire N__47736;
    wire N__47733;
    wire N__47732;
    wire N__47731;
    wire N__47730;
    wire N__47729;
    wire N__47728;
    wire N__47727;
    wire N__47726;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47722;
    wire N__47721;
    wire N__47720;
    wire N__47717;
    wire N__47716;
    wire N__47715;
    wire N__47712;
    wire N__47711;
    wire N__47700;
    wire N__47697;
    wire N__47696;
    wire N__47691;
    wire N__47688;
    wire N__47683;
    wire N__47680;
    wire N__47673;
    wire N__47670;
    wire N__47667;
    wire N__47662;
    wire N__47659;
    wire N__47658;
    wire N__47657;
    wire N__47656;
    wire N__47655;
    wire N__47654;
    wire N__47653;
    wire N__47652;
    wire N__47649;
    wire N__47648;
    wire N__47647;
    wire N__47642;
    wire N__47637;
    wire N__47628;
    wire N__47623;
    wire N__47616;
    wire N__47613;
    wire N__47612;
    wire N__47611;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47599;
    wire N__47598;
    wire N__47597;
    wire N__47594;
    wire N__47585;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47571;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47554;
    wire N__47545;
    wire N__47538;
    wire N__47535;
    wire N__47532;
    wire N__47527;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47501;
    wire N__47498;
    wire N__47497;
    wire N__47494;
    wire N__47489;
    wire N__47486;
    wire N__47485;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47468;
    wire N__47465;
    wire N__47462;
    wire N__47457;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47430;
    wire N__47429;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47415;
    wire N__47412;
    wire N__47409;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47355;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47344;
    wire N__47343;
    wire N__47336;
    wire N__47333;
    wire N__47326;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47298;
    wire N__47295;
    wire N__47294;
    wire N__47293;
    wire N__47290;
    wire N__47287;
    wire N__47278;
    wire N__47277;
    wire N__47276;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47234;
    wire N__47233;
    wire N__47232;
    wire N__47231;
    wire N__47228;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47212;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47191;
    wire N__47188;
    wire N__47183;
    wire N__47180;
    wire N__47179;
    wire N__47174;
    wire N__47167;
    wire N__47164;
    wire N__47159;
    wire N__47154;
    wire N__47151;
    wire N__47150;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47142;
    wire N__47139;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47103;
    wire N__47102;
    wire N__47099;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47077;
    wire N__47072;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47057;
    wire N__47054;
    wire N__47053;
    wire N__47052;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47040;
    wire N__47037;
    wire N__47028;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47014;
    wire N__47013;
    wire N__47012;
    wire N__47011;
    wire N__47008;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46979;
    wire N__46976;
    wire N__46969;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46955;
    wire N__46954;
    wire N__46953;
    wire N__46950;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46929;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46915;
    wire N__46910;
    wire N__46907;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46897;
    wire N__46894;
    wire N__46887;
    wire N__46884;
    wire N__46883;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46874;
    wire N__46873;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46854;
    wire N__46851;
    wire N__46846;
    wire N__46841;
    wire N__46836;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46815;
    wire N__46808;
    wire N__46801;
    wire N__46800;
    wire N__46797;
    wire N__46792;
    wire N__46791;
    wire N__46790;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46762;
    wire N__46759;
    wire N__46752;
    wire N__46749;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46743;
    wire N__46742;
    wire N__46741;
    wire N__46740;
    wire N__46737;
    wire N__46732;
    wire N__46723;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46696;
    wire N__46691;
    wire N__46688;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46670;
    wire N__46667;
    wire N__46664;
    wire N__46661;
    wire N__46656;
    wire N__46653;
    wire N__46652;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46635;
    wire N__46632;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46610;
    wire N__46609;
    wire N__46608;
    wire N__46607;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46599;
    wire N__46594;
    wire N__46591;
    wire N__46590;
    wire N__46587;
    wire N__46582;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46557;
    wire N__46554;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46522;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46505;
    wire N__46500;
    wire N__46499;
    wire N__46498;
    wire N__46493;
    wire N__46490;
    wire N__46485;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46479;
    wire N__46478;
    wire N__46475;
    wire N__46466;
    wire N__46461;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46449;
    wire N__46448;
    wire N__46445;
    wire N__46444;
    wire N__46441;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46395;
    wire N__46392;
    wire N__46391;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46379;
    wire N__46378;
    wire N__46373;
    wire N__46370;
    wire N__46365;
    wire N__46362;
    wire N__46361;
    wire N__46358;
    wire N__46357;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46349;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46315;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46297;
    wire N__46294;
    wire N__46289;
    wire N__46286;
    wire N__46281;
    wire N__46272;
    wire N__46271;
    wire N__46270;
    wire N__46265;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46247;
    wire N__46244;
    wire N__46241;
    wire N__46236;
    wire N__46233;
    wire N__46228;
    wire N__46221;
    wire N__46220;
    wire N__46217;
    wire N__46214;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46204;
    wire N__46199;
    wire N__46196;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46184;
    wire N__46183;
    wire N__46180;
    wire N__46179;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46151;
    wire N__46148;
    wire N__46145;
    wire N__46140;
    wire N__46139;
    wire N__46136;
    wire N__46135;
    wire N__46134;
    wire N__46133;
    wire N__46132;
    wire N__46129;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46106;
    wire N__46101;
    wire N__46098;
    wire N__46097;
    wire N__46096;
    wire N__46095;
    wire N__46094;
    wire N__46093;
    wire N__46092;
    wire N__46091;
    wire N__46090;
    wire N__46089;
    wire N__46088;
    wire N__46087;
    wire N__46086;
    wire N__46085;
    wire N__46084;
    wire N__46083;
    wire N__46080;
    wire N__46079;
    wire N__46078;
    wire N__46071;
    wire N__46064;
    wire N__46063;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46058;
    wire N__46057;
    wire N__46056;
    wire N__46055;
    wire N__46052;
    wire N__46051;
    wire N__46050;
    wire N__46049;
    wire N__46048;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46027;
    wire N__46026;
    wire N__46025;
    wire N__46024;
    wire N__46023;
    wire N__46022;
    wire N__46021;
    wire N__46020;
    wire N__46019;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46011;
    wire N__46010;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45990;
    wire N__45989;
    wire N__45988;
    wire N__45987;
    wire N__45986;
    wire N__45985;
    wire N__45984;
    wire N__45983;
    wire N__45972;
    wire N__45963;
    wire N__45960;
    wire N__45949;
    wire N__45946;
    wire N__45945;
    wire N__45940;
    wire N__45937;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45922;
    wire N__45919;
    wire N__45914;
    wire N__45907;
    wire N__45902;
    wire N__45897;
    wire N__45890;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45882;
    wire N__45881;
    wire N__45880;
    wire N__45879;
    wire N__45878;
    wire N__45877;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45873;
    wire N__45872;
    wire N__45871;
    wire N__45864;
    wire N__45859;
    wire N__45852;
    wire N__45839;
    wire N__45832;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45796;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45775;
    wire N__45766;
    wire N__45755;
    wire N__45752;
    wire N__45741;
    wire N__45734;
    wire N__45723;
    wire N__45718;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45627;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45615;
    wire N__45614;
    wire N__45613;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45602;
    wire N__45599;
    wire N__45598;
    wire N__45595;
    wire N__45592;
    wire N__45591;
    wire N__45588;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45556;
    wire N__45549;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45519;
    wire N__45518;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45508;
    wire N__45507;
    wire N__45506;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45480;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45453;
    wire N__45444;
    wire N__45441;
    wire N__45440;
    wire N__45439;
    wire N__45438;
    wire N__45437;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45411;
    wire N__45408;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45382;
    wire N__45381;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45368;
    wire N__45365;
    wire N__45362;
    wire N__45357;
    wire N__45348;
    wire N__45345;
    wire N__45344;
    wire N__45341;
    wire N__45340;
    wire N__45337;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45323;
    wire N__45322;
    wire N__45321;
    wire N__45316;
    wire N__45311;
    wire N__45308;
    wire N__45305;
    wire N__45302;
    wire N__45297;
    wire N__45294;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45263;
    wire N__45262;
    wire N__45261;
    wire N__45260;
    wire N__45257;
    wire N__45254;
    wire N__45251;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45230;
    wire N__45229;
    wire N__45228;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45185;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45174;
    wire N__45173;
    wire N__45170;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45137;
    wire N__45132;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45059;
    wire N__45056;
    wire N__45055;
    wire N__45054;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45043;
    wire N__45042;
    wire N__45041;
    wire N__45038;
    wire N__45037;
    wire N__45036;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45028;
    wire N__45027;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44996;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44975;
    wire N__44972;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44956;
    wire N__44953;
    wire N__44948;
    wire N__44945;
    wire N__44938;
    wire N__44931;
    wire N__44926;
    wire N__44923;
    wire N__44920;
    wire N__44917;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44896;
    wire N__44891;
    wire N__44888;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44864;
    wire N__44863;
    wire N__44862;
    wire N__44861;
    wire N__44858;
    wire N__44855;
    wire N__44852;
    wire N__44847;
    wire N__44846;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44831;
    wire N__44830;
    wire N__44827;
    wire N__44822;
    wire N__44815;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44798;
    wire N__44793;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44774;
    wire N__44773;
    wire N__44770;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44762;
    wire N__44759;
    wire N__44756;
    wire N__44755;
    wire N__44750;
    wire N__44747;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44732;
    wire N__44727;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44708;
    wire N__44707;
    wire N__44704;
    wire N__44703;
    wire N__44700;
    wire N__44699;
    wire N__44696;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44686;
    wire N__44685;
    wire N__44684;
    wire N__44683;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44668;
    wire N__44665;
    wire N__44660;
    wire N__44657;
    wire N__44652;
    wire N__44645;
    wire N__44642;
    wire N__44631;
    wire N__44628;
    wire N__44627;
    wire N__44626;
    wire N__44623;
    wire N__44618;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44559;
    wire N__44558;
    wire N__44557;
    wire N__44554;
    wire N__44549;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44526;
    wire N__44525;
    wire N__44522;
    wire N__44519;
    wire N__44514;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44492;
    wire N__44489;
    wire N__44486;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44466;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44409;
    wire N__44406;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44331;
    wire N__44328;
    wire N__44327;
    wire N__44326;
    wire N__44325;
    wire N__44322;
    wire N__44315;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44225;
    wire N__44222;
    wire N__44221;
    wire N__44220;
    wire N__44219;
    wire N__44218;
    wire N__44217;
    wire N__44214;
    wire N__44205;
    wire N__44202;
    wire N__44201;
    wire N__44198;
    wire N__44197;
    wire N__44196;
    wire N__44195;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44179;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44159;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44142;
    wire N__44141;
    wire N__44138;
    wire N__44135;
    wire N__44132;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44109;
    wire N__44108;
    wire N__44105;
    wire N__44104;
    wire N__44103;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44067;
    wire N__44058;
    wire N__44057;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44046;
    wire N__44045;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44013;
    wire N__44012;
    wire N__44011;
    wire N__44008;
    wire N__44005;
    wire N__44004;
    wire N__44003;
    wire N__44002;
    wire N__43999;
    wire N__43998;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43969;
    wire N__43968;
    wire N__43967;
    wire N__43964;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43939;
    wire N__43926;
    wire N__43925;
    wire N__43924;
    wire N__43923;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43896;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43880;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43842;
    wire N__43839;
    wire N__43838;
    wire N__43837;
    wire N__43836;
    wire N__43835;
    wire N__43834;
    wire N__43831;
    wire N__43830;
    wire N__43829;
    wire N__43826;
    wire N__43825;
    wire N__43824;
    wire N__43821;
    wire N__43820;
    wire N__43817;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43773;
    wire N__43770;
    wire N__43765;
    wire N__43760;
    wire N__43757;
    wire N__43754;
    wire N__43753;
    wire N__43752;
    wire N__43737;
    wire N__43734;
    wire N__43727;
    wire N__43722;
    wire N__43719;
    wire N__43710;
    wire N__43709;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43698;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43671;
    wire N__43668;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43656;
    wire N__43655;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43610;
    wire N__43609;
    wire N__43606;
    wire N__43605;
    wire N__43604;
    wire N__43599;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43575;
    wire N__43572;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43532;
    wire N__43531;
    wire N__43530;
    wire N__43527;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43516;
    wire N__43515;
    wire N__43514;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43493;
    wire N__43492;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43478;
    wire N__43473;
    wire N__43468;
    wire N__43465;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43408;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43395;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43371;
    wire N__43368;
    wire N__43367;
    wire N__43364;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43347;
    wire N__43346;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43329;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43318;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43308;
    wire N__43305;
    wire N__43296;
    wire N__43293;
    wire N__43292;
    wire N__43289;
    wire N__43286;
    wire N__43285;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43275;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43256;
    wire N__43253;
    wire N__43248;
    wire N__43239;
    wire N__43238;
    wire N__43235;
    wire N__43234;
    wire N__43233;
    wire N__43232;
    wire N__43231;
    wire N__43230;
    wire N__43229;
    wire N__43228;
    wire N__43227;
    wire N__43224;
    wire N__43223;
    wire N__43222;
    wire N__43221;
    wire N__43220;
    wire N__43219;
    wire N__43218;
    wire N__43217;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43206;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43186;
    wire N__43183;
    wire N__43182;
    wire N__43181;
    wire N__43180;
    wire N__43179;
    wire N__43178;
    wire N__43177;
    wire N__43176;
    wire N__43175;
    wire N__43172;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43164;
    wire N__43161;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43114;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43087;
    wire N__43086;
    wire N__43085;
    wire N__43084;
    wire N__43081;
    wire N__43068;
    wire N__43063;
    wire N__43062;
    wire N__43061;
    wire N__43060;
    wire N__43055;
    wire N__43054;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43035;
    wire N__43034;
    wire N__43033;
    wire N__43032;
    wire N__43029;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43009;
    wire N__43006;
    wire N__43001;
    wire N__42998;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42979;
    wire N__42974;
    wire N__42967;
    wire N__42960;
    wire N__42953;
    wire N__42948;
    wire N__42943;
    wire N__42924;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42909;
    wire N__42906;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42856;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42834;
    wire N__42831;
    wire N__42822;
    wire N__42819;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42771;
    wire N__42770;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42738;
    wire N__42733;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42704;
    wire N__42703;
    wire N__42702;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42688;
    wire N__42685;
    wire N__42680;
    wire N__42675;
    wire N__42672;
    wire N__42663;
    wire N__42660;
    wire N__42659;
    wire N__42658;
    wire N__42657;
    wire N__42656;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42632;
    wire N__42629;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42611;
    wire N__42608;
    wire N__42605;
    wire N__42602;
    wire N__42601;
    wire N__42598;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42580;
    wire N__42577;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42560;
    wire N__42559;
    wire N__42556;
    wire N__42553;
    wire N__42552;
    wire N__42549;
    wire N__42544;
    wire N__42541;
    wire N__42538;
    wire N__42537;
    wire N__42536;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42509;
    wire N__42498;
    wire N__42497;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42474;
    wire N__42471;
    wire N__42470;
    wire N__42467;
    wire N__42466;
    wire N__42463;
    wire N__42462;
    wire N__42459;
    wire N__42454;
    wire N__42451;
    wire N__42448;
    wire N__42445;
    wire N__42438;
    wire N__42437;
    wire N__42436;
    wire N__42431;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42418;
    wire N__42415;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42401;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42391;
    wire N__42390;
    wire N__42389;
    wire N__42382;
    wire N__42381;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42366;
    wire N__42363;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42341;
    wire N__42338;
    wire N__42335;
    wire N__42330;
    wire N__42329;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42313;
    wire N__42308;
    wire N__42307;
    wire N__42304;
    wire N__42301;
    wire N__42298;
    wire N__42297;
    wire N__42292;
    wire N__42289;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42267;
    wire N__42264;
    wire N__42263;
    wire N__42262;
    wire N__42261;
    wire N__42258;
    wire N__42257;
    wire N__42254;
    wire N__42251;
    wire N__42248;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42216;
    wire N__42207;
    wire N__42204;
    wire N__42201;
    wire N__42200;
    wire N__42195;
    wire N__42194;
    wire N__42193;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42174;
    wire N__42171;
    wire N__42170;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42123;
    wire N__42122;
    wire N__42121;
    wire N__42118;
    wire N__42115;
    wire N__42114;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42093;
    wire N__42092;
    wire N__42091;
    wire N__42088;
    wire N__42083;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42065;
    wire N__42064;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42049;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42026;
    wire N__42023;
    wire N__42022;
    wire N__42019;
    wire N__42018;
    wire N__42017;
    wire N__42014;
    wire N__42011;
    wire N__42008;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41967;
    wire N__41964;
    wire N__41959;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41945;
    wire N__41944;
    wire N__41943;
    wire N__41940;
    wire N__41935;
    wire N__41932;
    wire N__41925;
    wire N__41922;
    wire N__41921;
    wire N__41916;
    wire N__41913;
    wire N__41912;
    wire N__41911;
    wire N__41908;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41890;
    wire N__41885;
    wire N__41882;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41820;
    wire N__41815;
    wire N__41810;
    wire N__41805;
    wire N__41802;
    wire N__41801;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41789;
    wire N__41786;
    wire N__41781;
    wire N__41780;
    wire N__41779;
    wire N__41776;
    wire N__41773;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41753;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41718;
    wire N__41715;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41705;
    wire N__41700;
    wire N__41699;
    wire N__41698;
    wire N__41695;
    wire N__41692;
    wire N__41689;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41564;
    wire N__41563;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41551;
    wire N__41546;
    wire N__41541;
    wire N__41538;
    wire N__41537;
    wire N__41536;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41524;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41496;
    wire N__41495;
    wire N__41492;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41436;
    wire N__41433;
    wire N__41432;
    wire N__41431;
    wire N__41430;
    wire N__41429;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41413;
    wire N__41412;
    wire N__41409;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41386;
    wire N__41383;
    wire N__41378;
    wire N__41375;
    wire N__41370;
    wire N__41367;
    wire N__41366;
    wire N__41365;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41352;
    wire N__41347;
    wire N__41342;
    wire N__41339;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41327;
    wire N__41326;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41318;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41267;
    wire N__41262;
    wire N__41261;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41231;
    wire N__41230;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41197;
    wire N__41190;
    wire N__41189;
    wire N__41186;
    wire N__41185;
    wire N__41182;
    wire N__41181;
    wire N__41180;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41172;
    wire N__41169;
    wire N__41164;
    wire N__41161;
    wire N__41156;
    wire N__41153;
    wire N__41148;
    wire N__41143;
    wire N__41140;
    wire N__41139;
    wire N__41136;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41108;
    wire N__41107;
    wire N__41106;
    wire N__41105;
    wire N__41104;
    wire N__41103;
    wire N__41102;
    wire N__41099;
    wire N__41094;
    wire N__41089;
    wire N__41086;
    wire N__41081;
    wire N__41074;
    wire N__41067;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41055;
    wire N__41054;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41046;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41038;
    wire N__41035;
    wire N__41034;
    wire N__41033;
    wire N__41030;
    wire N__41027;
    wire N__41026;
    wire N__41025;
    wire N__41024;
    wire N__41023;
    wire N__41022;
    wire N__41021;
    wire N__41020;
    wire N__41019;
    wire N__41018;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41010;
    wire N__41009;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__41001;
    wire N__41000;
    wire N__40997;
    wire N__40996;
    wire N__40995;
    wire N__40994;
    wire N__40991;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40973;
    wire N__40966;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40950;
    wire N__40949;
    wire N__40946;
    wire N__40941;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40920;
    wire N__40913;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40890;
    wire N__40883;
    wire N__40880;
    wire N__40867;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40826;
    wire N__40823;
    wire N__40822;
    wire N__40821;
    wire N__40820;
    wire N__40819;
    wire N__40818;
    wire N__40817;
    wire N__40816;
    wire N__40815;
    wire N__40812;
    wire N__40811;
    wire N__40810;
    wire N__40809;
    wire N__40808;
    wire N__40807;
    wire N__40806;
    wire N__40805;
    wire N__40804;
    wire N__40801;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40782;
    wire N__40781;
    wire N__40780;
    wire N__40779;
    wire N__40778;
    wire N__40777;
    wire N__40776;
    wire N__40775;
    wire N__40774;
    wire N__40773;
    wire N__40772;
    wire N__40771;
    wire N__40770;
    wire N__40769;
    wire N__40768;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40746;
    wire N__40741;
    wire N__40736;
    wire N__40727;
    wire N__40720;
    wire N__40715;
    wire N__40706;
    wire N__40703;
    wire N__40694;
    wire N__40689;
    wire N__40686;
    wire N__40685;
    wire N__40684;
    wire N__40681;
    wire N__40672;
    wire N__40667;
    wire N__40654;
    wire N__40651;
    wire N__40650;
    wire N__40649;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40634;
    wire N__40627;
    wire N__40624;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40570;
    wire N__40569;
    wire N__40568;
    wire N__40567;
    wire N__40566;
    wire N__40565;
    wire N__40564;
    wire N__40563;
    wire N__40562;
    wire N__40559;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40545;
    wire N__40544;
    wire N__40543;
    wire N__40542;
    wire N__40541;
    wire N__40540;
    wire N__40537;
    wire N__40536;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40528;
    wire N__40527;
    wire N__40526;
    wire N__40519;
    wire N__40516;
    wire N__40513;
    wire N__40504;
    wire N__40499;
    wire N__40494;
    wire N__40489;
    wire N__40486;
    wire N__40485;
    wire N__40480;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40468;
    wire N__40467;
    wire N__40464;
    wire N__40457;
    wire N__40452;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40426;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40413;
    wire N__40412;
    wire N__40411;
    wire N__40410;
    wire N__40409;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40391;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40355;
    wire N__40352;
    wire N__40335;
    wire N__40332;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40267;
    wire N__40266;
    wire N__40265;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40241;
    wire N__40236;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40214;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40206;
    wire N__40205;
    wire N__40204;
    wire N__40201;
    wire N__40196;
    wire N__40193;
    wire N__40188;
    wire N__40179;
    wire N__40178;
    wire N__40175;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40148;
    wire N__40145;
    wire N__40144;
    wire N__40143;
    wire N__40138;
    wire N__40133;
    wire N__40128;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40103;
    wire N__40098;
    wire N__40095;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40084;
    wire N__40081;
    wire N__40080;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40070;
    wire N__40065;
    wire N__40064;
    wire N__40059;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40023;
    wire N__40022;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39995;
    wire N__39990;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39944;
    wire N__39939;
    wire N__39936;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39899;
    wire N__39896;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39841;
    wire N__39840;
    wire N__39837;
    wire N__39836;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39798;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39780;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39755;
    wire N__39754;
    wire N__39751;
    wire N__39746;
    wire N__39745;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39626;
    wire N__39625;
    wire N__39624;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39613;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39599;
    wire N__39596;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39581;
    wire N__39578;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39554;
    wire N__39553;
    wire N__39550;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39529;
    wire N__39526;
    wire N__39521;
    wire N__39516;
    wire N__39513;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39441;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39423;
    wire N__39422;
    wire N__39421;
    wire N__39418;
    wire N__39413;
    wire N__39412;
    wire N__39407;
    wire N__39404;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39375;
    wire N__39372;
    wire N__39371;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39353;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39335;
    wire N__39334;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39322;
    wire N__39315;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39301;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39289;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39258;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39206;
    wire N__39203;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39170;
    wire N__39169;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39144;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39113;
    wire N__39112;
    wire N__39111;
    wire N__39110;
    wire N__39109;
    wire N__39108;
    wire N__39103;
    wire N__39098;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39090;
    wire N__39089;
    wire N__39088;
    wire N__39085;
    wire N__39080;
    wire N__39077;
    wire N__39072;
    wire N__39071;
    wire N__39068;
    wire N__39063;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39039;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39021;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39009;
    wire N__39008;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38988;
    wire N__38987;
    wire N__38982;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38967;
    wire N__38966;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38954;
    wire N__38953;
    wire N__38952;
    wire N__38951;
    wire N__38948;
    wire N__38947;
    wire N__38946;
    wire N__38945;
    wire N__38944;
    wire N__38935;
    wire N__38934;
    wire N__38933;
    wire N__38930;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38914;
    wire N__38913;
    wire N__38910;
    wire N__38905;
    wire N__38900;
    wire N__38895;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38879;
    wire N__38876;
    wire N__38875;
    wire N__38872;
    wire N__38869;
    wire N__38868;
    wire N__38865;
    wire N__38860;
    wire N__38857;
    wire N__38852;
    wire N__38847;
    wire N__38846;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38810;
    wire N__38809;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38788;
    wire N__38787;
    wire N__38782;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38763;
    wire N__38762;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38743;
    wire N__38736;
    wire N__38735;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38718;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38697;
    wire N__38694;
    wire N__38693;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38675;
    wire N__38674;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38649;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38631;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38548;
    wire N__38543;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38515;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38483;
    wire N__38482;
    wire N__38479;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38471;
    wire N__38468;
    wire N__38467;
    wire N__38464;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38446;
    wire N__38443;
    wire N__38438;
    wire N__38435;
    wire N__38430;
    wire N__38427;
    wire N__38420;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38393;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38366;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38344;
    wire N__38343;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38319;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38307;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38292;
    wire N__38289;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38264;
    wire N__38263;
    wire N__38262;
    wire N__38259;
    wire N__38258;
    wire N__38255;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38234;
    wire N__38229;
    wire N__38228;
    wire N__38227;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38190;
    wire N__38189;
    wire N__38186;
    wire N__38185;
    wire N__38184;
    wire N__38181;
    wire N__38180;
    wire N__38179;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38175;
    wire N__38174;
    wire N__38169;
    wire N__38166;
    wire N__38165;
    wire N__38164;
    wire N__38155;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38139;
    wire N__38134;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38122;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38101;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38089;
    wire N__38084;
    wire N__38083;
    wire N__38082;
    wire N__38077;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38063;
    wire N__38060;
    wire N__38059;
    wire N__38052;
    wire N__38049;
    wire N__38046;
    wire N__38043;
    wire N__38038;
    wire N__38031;
    wire N__38030;
    wire N__38029;
    wire N__38026;
    wire N__38025;
    wire N__38022;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38011;
    wire N__38010;
    wire N__38007;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37995;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37939;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37927;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37906;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37865;
    wire N__37862;
    wire N__37861;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37826;
    wire N__37823;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37812;
    wire N__37809;
    wire N__37804;
    wire N__37801;
    wire N__37796;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37761;
    wire N__37758;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37743;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37653;
    wire N__37652;
    wire N__37649;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37601;
    wire N__37598;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37581;
    wire N__37578;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37560;
    wire N__37557;
    wire N__37556;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37487;
    wire N__37486;
    wire N__37485;
    wire N__37484;
    wire N__37483;
    wire N__37480;
    wire N__37479;
    wire N__37478;
    wire N__37475;
    wire N__37474;
    wire N__37471;
    wire N__37470;
    wire N__37467;
    wire N__37466;
    wire N__37463;
    wire N__37462;
    wire N__37459;
    wire N__37458;
    wire N__37455;
    wire N__37454;
    wire N__37451;
    wire N__37450;
    wire N__37449;
    wire N__37448;
    wire N__37447;
    wire N__37446;
    wire N__37445;
    wire N__37444;
    wire N__37441;
    wire N__37436;
    wire N__37423;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37384;
    wire N__37383;
    wire N__37382;
    wire N__37381;
    wire N__37380;
    wire N__37371;
    wire N__37362;
    wire N__37353;
    wire N__37350;
    wire N__37349;
    wire N__37346;
    wire N__37345;
    wire N__37342;
    wire N__37341;
    wire N__37338;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37311;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37235;
    wire N__37232;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37188;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37170;
    wire N__37169;
    wire N__37168;
    wire N__37165;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37153;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37139;
    wire N__37138;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37120;
    wire N__37117;
    wire N__37116;
    wire N__37115;
    wire N__37112;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37092;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37035;
    wire N__37034;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37022;
    wire N__37017;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36977;
    wire N__36976;
    wire N__36975;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36957;
    wire N__36952;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36923;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36857;
    wire N__36852;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36788;
    wire N__36785;
    wire N__36784;
    wire N__36781;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36760;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36707;
    wire N__36706;
    wire N__36703;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36693;
    wire N__36690;
    wire N__36689;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36659;
    wire N__36652;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36623;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36599;
    wire N__36598;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36586;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36540;
    wire N__36537;
    wire N__36532;
    wire N__36529;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36490;
    wire N__36489;
    wire N__36488;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36460;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36422;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36414;
    wire N__36413;
    wire N__36410;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36394;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36342;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36266;
    wire N__36265;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36249;
    wire N__36246;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36159;
    wire N__36156;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36144;
    wire N__36141;
    wire N__36138;
    wire N__36133;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36080;
    wire N__36077;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36031;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35964;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35901;
    wire N__35898;
    wire N__35897;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35810;
    wire N__35805;
    wire N__35802;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35770;
    wire N__35761;
    wire N__35758;
    wire N__35757;
    wire N__35756;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35721;
    wire N__35720;
    wire N__35719;
    wire N__35716;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35694;
    wire N__35691;
    wire N__35690;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35669;
    wire N__35664;
    wire N__35663;
    wire N__35662;
    wire N__35659;
    wire N__35654;
    wire N__35653;
    wire N__35652;
    wire N__35651;
    wire N__35646;
    wire N__35641;
    wire N__35638;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35616;
    wire N__35615;
    wire N__35614;
    wire N__35611;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35597;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35554;
    wire N__35551;
    wire N__35546;
    wire N__35545;
    wire N__35544;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35523;
    wire N__35520;
    wire N__35519;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35472;
    wire N__35471;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35453;
    wire N__35450;
    wire N__35443;
    wire N__35438;
    wire N__35435;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35417;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35385;
    wire N__35382;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35353;
    wire N__35348;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35330;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35298;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35287;
    wire N__35286;
    wire N__35285;
    wire N__35284;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35269;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35258;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35240;
    wire N__35235;
    wire N__35226;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35216;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35194;
    wire N__35189;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35148;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35133;
    wire N__35132;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35117;
    wire N__35116;
    wire N__35113;
    wire N__35112;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35096;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35064;
    wire N__35061;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35035;
    wire N__35034;
    wire N__35033;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35018;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__34995;
    wire N__34992;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34977;
    wire N__34976;
    wire N__34975;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34963;
    wire N__34960;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34888;
    wire N__34885;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34860;
    wire N__34857;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34842;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34817;
    wire N__34816;
    wire N__34815;
    wire N__34814;
    wire N__34811;
    wire N__34806;
    wire N__34805;
    wire N__34800;
    wire N__34795;
    wire N__34792;
    wire N__34785;
    wire N__34782;
    wire N__34781;
    wire N__34780;
    wire N__34777;
    wire N__34776;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34746;
    wire N__34741;
    wire N__34738;
    wire N__34737;
    wire N__34734;
    wire N__34729;
    wire N__34726;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34695;
    wire N__34692;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34677;
    wire N__34674;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34659;
    wire N__34656;
    wire N__34655;
    wire N__34654;
    wire N__34651;
    wire N__34650;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34623;
    wire N__34614;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34561;
    wire N__34548;
    wire N__34545;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34437;
    wire N__34434;
    wire N__34433;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34425;
    wire N__34422;
    wire N__34421;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34356;
    wire N__34353;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34345;
    wire N__34344;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34251;
    wire N__34248;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34196;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34154;
    wire N__34151;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34122;
    wire N__34113;
    wire N__34110;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34091;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34083;
    wire N__34080;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34029;
    wire N__34028;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33995;
    wire N__33994;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33954;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33946;
    wire N__33943;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33925;
    wire N__33922;
    wire N__33915;
    wire N__33912;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33870;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33855;
    wire N__33854;
    wire N__33853;
    wire N__33852;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33799;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33781;
    wire N__33778;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33716;
    wire N__33715;
    wire N__33712;
    wire N__33707;
    wire N__33702;
    wire N__33701;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33686;
    wire N__33683;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33645;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33620;
    wire N__33615;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33593;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33552;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33544;
    wire N__33543;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33525;
    wire N__33524;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33501;
    wire N__33500;
    wire N__33499;
    wire N__33496;
    wire N__33491;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33470;
    wire N__33467;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33402;
    wire N__33399;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33342;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33327;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33315;
    wire N__33312;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33258;
    wire N__33255;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33219;
    wire N__33216;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33140;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33134;
    wire N__33133;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33126;
    wire N__33125;
    wire N__33122;
    wire N__33121;
    wire N__33118;
    wire N__33117;
    wire N__33114;
    wire N__33113;
    wire N__33110;
    wire N__33109;
    wire N__33106;
    wire N__33105;
    wire N__33102;
    wire N__33101;
    wire N__33098;
    wire N__33097;
    wire N__33094;
    wire N__33093;
    wire N__33090;
    wire N__33089;
    wire N__33086;
    wire N__33085;
    wire N__33082;
    wire N__33081;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33073;
    wire N__33072;
    wire N__33071;
    wire N__33068;
    wire N__33051;
    wire N__33034;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32995;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32975;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32941;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32888;
    wire N__32885;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32863;
    wire N__32858;
    wire N__32853;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32830;
    wire N__32827;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32707;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32695;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32673;
    wire N__32670;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32459;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32345;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32319;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32301;
    wire N__32298;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32261;
    wire N__32260;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32248;
    wire N__32245;
    wire N__32240;
    wire N__32235;
    wire N__32234;
    wire N__32233;
    wire N__32232;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32200;
    wire N__32197;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32141;
    wire N__32140;
    wire N__32139;
    wire N__32138;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32003;
    wire N__32002;
    wire N__32001;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31980;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31944;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31900;
    wire N__31899;
    wire N__31898;
    wire N__31895;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31871;
    wire N__31868;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31805;
    wire N__31804;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31792;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31775;
    wire N__31774;
    wire N__31773;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31752;
    wire N__31749;
    wire N__31748;
    wire N__31747;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31735;
    wire N__31732;
    wire N__31725;
    wire N__31722;
    wire N__31721;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31702;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31688;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31563;
    wire N__31560;
    wire N__31559;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31546;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31446;
    wire N__31445;
    wire N__31442;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31418;
    wire N__31417;
    wire N__31416;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31396;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31352;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31332;
    wire N__31329;
    wire N__31328;
    wire N__31325;
    wire N__31324;
    wire N__31323;
    wire N__31320;
    wire N__31319;
    wire N__31318;
    wire N__31317;
    wire N__31316;
    wire N__31315;
    wire N__31314;
    wire N__31313;
    wire N__31312;
    wire N__31305;
    wire N__31304;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31286;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31271;
    wire N__31270;
    wire N__31267;
    wire N__31266;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31226;
    wire N__31219;
    wire N__31214;
    wire N__31211;
    wire N__31200;
    wire N__31199;
    wire N__31198;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31190;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31178;
    wire N__31177;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31162;
    wire N__31159;
    wire N__31158;
    wire N__31157;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31120;
    wire N__31115;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30911;
    wire N__30906;
    wire N__30903;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30839;
    wire N__30836;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30824;
    wire N__30823;
    wire N__30820;
    wire N__30815;
    wire N__30810;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30773;
    wire N__30772;
    wire N__30767;
    wire N__30764;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30732;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30656;
    wire N__30653;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30614;
    wire N__30609;
    wire N__30608;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30577;
    wire N__30574;
    wire N__30569;
    wire N__30566;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30555;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30521;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30404;
    wire N__30399;
    wire N__30396;
    wire N__30395;
    wire N__30390;
    wire N__30387;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30359;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30269;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30240;
    wire N__30237;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30222;
    wire N__30221;
    wire N__30218;
    wire N__30217;
    wire N__30214;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30203;
    wire N__30202;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30147;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30139;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30131;
    wire N__30130;
    wire N__30129;
    wire N__30126;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30099;
    wire N__30096;
    wire N__30091;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30018;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29892;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29856;
    wire N__29853;
    wire N__29852;
    wire N__29847;
    wire N__29846;
    wire N__29845;
    wire N__29842;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29817;
    wire N__29816;
    wire N__29815;
    wire N__29810;
    wire N__29807;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29778;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29727;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29715;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29700;
    wire N__29699;
    wire N__29698;
    wire N__29695;
    wire N__29690;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29664;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29652;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29637;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29607;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29595;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29580;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29550;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29538;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29523;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29405;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29277;
    wire N__29274;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29259;
    wire N__29258;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29246;
    wire N__29245;
    wire N__29244;
    wire N__29243;
    wire N__29242;
    wire N__29241;
    wire N__29240;
    wire N__29239;
    wire N__29232;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29220;
    wire N__29215;
    wire N__29214;
    wire N__29213;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29187;
    wire N__29180;
    wire N__29175;
    wire N__29172;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29112;
    wire N__29109;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29088;
    wire N__29085;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29070;
    wire N__29067;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29055;
    wire N__29052;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29040;
    wire N__29037;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28993;
    wire N__28988;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28965;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28952;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28876;
    wire N__28875;
    wire N__28872;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28824;
    wire N__28821;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28802;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28787;
    wire N__28782;
    wire N__28779;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28763;
    wire N__28758;
    wire N__28757;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28735;
    wire N__28728;
    wire N__28727;
    wire N__28726;
    wire N__28723;
    wire N__28722;
    wire N__28721;
    wire N__28720;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28701;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28685;
    wire N__28684;
    wire N__28683;
    wire N__28680;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28669;
    wire N__28668;
    wire N__28667;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28644;
    wire N__28641;
    wire N__28636;
    wire N__28633;
    wire N__28626;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28563;
    wire N__28560;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28532;
    wire N__28531;
    wire N__28530;
    wire N__28527;
    wire N__28520;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28463;
    wire N__28462;
    wire N__28459;
    wire N__28454;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28418;
    wire N__28415;
    wire N__28414;
    wire N__28411;
    wire N__28410;
    wire N__28407;
    wire N__28406;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28374;
    wire N__28373;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28358;
    wire N__28357;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28136;
    wire N__28135;
    wire N__28134;
    wire N__28133;
    wire N__28130;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28114;
    wire N__28111;
    wire N__28106;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28091;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28065;
    wire N__28064;
    wire N__28061;
    wire N__28060;
    wire N__28057;
    wire N__28052;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28029;
    wire N__28026;
    wire N__28025;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28008;
    wire N__28007;
    wire N__28004;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27984;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27969;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27942;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27920;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27909;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27855;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27843;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27831;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27816;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27786;
    wire N__27783;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27771;
    wire N__27768;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27756;
    wire N__27753;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27738;
    wire N__27735;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27723;
    wire N__27720;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27708;
    wire N__27705;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27693;
    wire N__27690;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27678;
    wire N__27675;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27663;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27635;
    wire N__27634;
    wire N__27631;
    wire N__27626;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27597;
    wire N__27594;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27579;
    wire N__27576;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27564;
    wire N__27561;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27546;
    wire N__27543;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27531;
    wire N__27528;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27453;
    wire N__27452;
    wire N__27449;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27417;
    wire N__27416;
    wire N__27413;
    wire N__27412;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27372;
    wire N__27369;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27327;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27282;
    wire N__27279;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27264;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27252;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27240;
    wire N__27237;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27225;
    wire N__27222;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27147;
    wire N__27144;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27096;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27082;
    wire N__27077;
    wire N__27074;
    wire N__27069;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27003;
    wire N__27000;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26943;
    wire N__26940;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26882;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26871;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26852;
    wire N__26849;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26837;
    wire N__26834;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26789;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire tx_enable;
    wire LED_c;
    wire \c0.rx.r_Rx_Data_R ;
    wire \quad_counter0.n22_cascade_ ;
    wire \quad_counter0.n25_adj_4760_cascade_ ;
    wire n12942_cascade_;
    wire \quad_counter0.n28_adj_4754 ;
    wire \quad_counter0.n26_adj_4755 ;
    wire \quad_counter0.n27_adj_4756_cascade_ ;
    wire \quad_counter0.n25_adj_4757 ;
    wire n9809_cascade_;
    wire n9809;
    wire \quad_counter1.n25_adj_4202_cascade_ ;
    wire n12940;
    wire PIN_13_c;
    wire n12940_cascade_;
    wire quadB_delayed_adj_4768;
    wire n14425_cascade_;
    wire \quad_counter1.n26_adj_4200 ;
    wire b_delay_counter_0_adj_4766;
    wire n187_adj_4771;
    wire bfn_5_17_0_;
    wire \quad_counter1.n19686 ;
    wire \quad_counter1.n19687 ;
    wire \quad_counter1.b_delay_counter_3 ;
    wire \quad_counter1.n19688 ;
    wire \quad_counter1.b_delay_counter_4 ;
    wire \quad_counter1.n19689 ;
    wire \quad_counter1.n19690 ;
    wire \quad_counter1.b_delay_counter_6 ;
    wire \quad_counter1.n19691 ;
    wire \quad_counter1.n19692 ;
    wire \quad_counter1.n19693 ;
    wire \quad_counter1.b_delay_counter_8 ;
    wire bfn_5_18_0_;
    wire \quad_counter1.b_delay_counter_9 ;
    wire \quad_counter1.n19694 ;
    wire \quad_counter1.b_delay_counter_10 ;
    wire \quad_counter1.n19695 ;
    wire \quad_counter1.b_delay_counter_11 ;
    wire \quad_counter1.n19696 ;
    wire \quad_counter1.n19697 ;
    wire \quad_counter1.n19698 ;
    wire \quad_counter1.n19699 ;
    wire \quad_counter1.n19700 ;
    wire n14425;
    wire b_delay_counter_15__N_4140_adj_4773;
    wire b_delay_counter_0;
    wire n187;
    wire bfn_6_10_0_;
    wire \quad_counter0.b_delay_counter_1 ;
    wire \quad_counter0.n19656 ;
    wire \quad_counter0.b_delay_counter_2 ;
    wire \quad_counter0.n19657 ;
    wire \quad_counter0.b_delay_counter_3 ;
    wire \quad_counter0.n19658 ;
    wire \quad_counter0.b_delay_counter_4 ;
    wire \quad_counter0.n19659 ;
    wire \quad_counter0.n19660 ;
    wire \quad_counter0.b_delay_counter_6 ;
    wire \quad_counter0.n19661 ;
    wire \quad_counter0.n19662 ;
    wire \quad_counter0.n19663 ;
    wire bfn_6_11_0_;
    wire \quad_counter0.b_delay_counter_9 ;
    wire \quad_counter0.n19664 ;
    wire \quad_counter0.n19665 ;
    wire \quad_counter0.n19666 ;
    wire \quad_counter0.n19667 ;
    wire \quad_counter0.b_delay_counter_13 ;
    wire \quad_counter0.n19668 ;
    wire \quad_counter0.n19669 ;
    wire \quad_counter0.n19670 ;
    wire n14315;
    wire b_delay_counter_15__N_4140;
    wire PIN_8_c;
    wire quadB_delayed;
    wire n12942;
    wire \quad_counter0.b_delay_counter_15 ;
    wire \quad_counter0.b_delay_counter_8 ;
    wire \quad_counter0.A_delayed ;
    wire \quad_counter0.b_delay_counter_7 ;
    wire \quad_counter0.b_delay_counter_12 ;
    wire \quad_counter0.b_delay_counter_5 ;
    wire \quad_counter0.b_delay_counter_14 ;
    wire \quad_counter0.b_delay_counter_10 ;
    wire \quad_counter0.b_delay_counter_11 ;
    wire \quad_counter0.n24_adj_4758_cascade_ ;
    wire \quad_counter0.n18 ;
    wire \quad_counter0.n26_adj_4759 ;
    wire a_delay_counter_0;
    wire n39;
    wire bfn_6_13_0_;
    wire \quad_counter0.a_delay_counter_1 ;
    wire \quad_counter0.n19671 ;
    wire \quad_counter0.a_delay_counter_2 ;
    wire \quad_counter0.n19672 ;
    wire \quad_counter0.a_delay_counter_3 ;
    wire \quad_counter0.n19673 ;
    wire \quad_counter0.a_delay_counter_4 ;
    wire \quad_counter0.n19674 ;
    wire \quad_counter0.a_delay_counter_5 ;
    wire \quad_counter0.n19675 ;
    wire \quad_counter0.a_delay_counter_6 ;
    wire \quad_counter0.n19676 ;
    wire \quad_counter0.a_delay_counter_7 ;
    wire \quad_counter0.n19677 ;
    wire \quad_counter0.n19678 ;
    wire \quad_counter0.a_delay_counter_8 ;
    wire bfn_6_14_0_;
    wire \quad_counter0.a_delay_counter_9 ;
    wire \quad_counter0.n19679 ;
    wire \quad_counter0.a_delay_counter_10 ;
    wire \quad_counter0.n19680 ;
    wire \quad_counter0.a_delay_counter_11 ;
    wire \quad_counter0.n19681 ;
    wire \quad_counter0.a_delay_counter_12 ;
    wire \quad_counter0.n19682 ;
    wire \quad_counter0.a_delay_counter_13 ;
    wire \quad_counter0.n19683 ;
    wire \quad_counter0.a_delay_counter_14 ;
    wire \quad_counter0.n19684 ;
    wire \quad_counter0.n19685 ;
    wire \quad_counter0.a_delay_counter_15 ;
    wire n14469;
    wire a_delay_counter_15__N_4123;
    wire \quad_counter1.b_delay_counter_13 ;
    wire \quad_counter1.b_delay_counter_1 ;
    wire \quad_counter1.b_delay_counter_2 ;
    wire \quad_counter1.b_delay_counter_5 ;
    wire \quad_counter1.n28_adj_4199 ;
    wire PIN_7_c;
    wire quadA_delayed;
    wire \quad_counter1.b_delay_counter_14 ;
    wire \quad_counter1.b_delay_counter_7 ;
    wire \quad_counter1.b_delay_counter_12 ;
    wire \quad_counter1.b_delay_counter_15 ;
    wire \quad_counter1.n27_adj_4201 ;
    wire A_filtered;
    wire n8628;
    wire n9603_cascade_;
    wire B_filtered;
    wire \quad_counter0.B_delayed ;
    wire n10_adj_4777;
    wire \c0.n25086_cascade_ ;
    wire data_out_frame_9_3;
    wire n24802_cascade_;
    wire \c0.n11_adj_4715_cascade_ ;
    wire n25010;
    wire \c0.tx.n6_cascade_ ;
    wire \c0.n25089 ;
    wire n25018;
    wire \c0.tx.n23980 ;
    wire \c0.n5_adj_4712_cascade_ ;
    wire \c0.n24800 ;
    wire \c0.tx.n5_adj_4207 ;
    wire \c0.n24949 ;
    wire \c0.n25104_cascade_ ;
    wire \c0.n25107 ;
    wire data_out_frame_5_7;
    wire n25071;
    wire n3821_cascade_;
    wire data_out_frame_9_7;
    wire \c0.rx.n24875 ;
    wire \c0.rx.n25068 ;
    wire bfn_9_7_0_;
    wire \quad_counter1.n19701 ;
    wire \quad_counter1.n19702 ;
    wire \quad_counter1.n19703 ;
    wire \quad_counter1.n19704 ;
    wire \quad_counter1.n19705 ;
    wire \quad_counter1.n19706 ;
    wire \quad_counter1.n19707 ;
    wire \quad_counter1.n19708 ;
    wire bfn_9_8_0_;
    wire \quad_counter1.n19709 ;
    wire \quad_counter1.n19710 ;
    wire \quad_counter1.n19711 ;
    wire \quad_counter1.n19712 ;
    wire \quad_counter1.n19713 ;
    wire \quad_counter1.n19714 ;
    wire \quad_counter1.n19715 ;
    wire \c0.tx.r_SM_Main_2 ;
    wire r_SM_Main_2_N_3751_1;
    wire \c0.tx.n3843 ;
    wire n3_cascade_;
    wire tx_o;
    wire r_Tx_Data_3;
    wire \c0.tx.n19492 ;
    wire \c0.tx.n22949 ;
    wire \c0.tx.n19492_cascade_ ;
    wire r_Tx_Data_1;
    wire \c0.tx.n25080 ;
    wire \c0.tx.n25083_cascade_ ;
    wire \c0.tx.o_Tx_Serial_N_3782 ;
    wire n10;
    wire \c0.tx.r_Bit_Index_2 ;
    wire \c0.tx.n17832 ;
    wire n10_adj_4776_cascade_;
    wire r_Tx_Data_5;
    wire \c0.tx.n25077 ;
    wire r_Tx_Data_7;
    wire \c0.tx.r_Bit_Index_0 ;
    wire \c0.tx.r_Bit_Index_1 ;
    wire \c0.tx.n25074 ;
    wire r_SM_Main_0;
    wire \c0.n24960_cascade_ ;
    wire \c0.n24806_cascade_ ;
    wire n24757;
    wire \c0.n26_adj_4645 ;
    wire n24808;
    wire n10_adj_4779;
    wire \c0.tx.n5_cascade_ ;
    wire \c0.tx.n17904 ;
    wire \c0.tx.n25051 ;
    wire bfn_9_16_0_;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.tx.n19723 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n19724 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.n19725 ;
    wire \c0.tx.r_Clock_Count_4 ;
    wire \c0.tx.n19726 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire \c0.tx.n19727 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire \c0.tx.n19728 ;
    wire \c0.tx.r_Clock_Count_7 ;
    wire \c0.tx.n19729 ;
    wire \c0.tx.n19730 ;
    wire bfn_9_17_0_;
    wire \c0.tx.r_Clock_Count_8 ;
    wire \c0.tx.n17199 ;
    wire \c0.tx.n4 ;
    wire \c0.tx.n14290_cascade_ ;
    wire data_out_frame_6_7;
    wire r_Tx_Data_6;
    wire data_out_frame_5_2;
    wire n17951;
    wire r_SM_Main_1_adj_4774;
    wire n25006;
    wire \c0.n11_adj_4663 ;
    wire data_out_frame_5_1;
    wire data_out_frame_13_3;
    wire data_out_frame_8_7;
    wire data_out_frame_12_6;
    wire \c0.n5_adj_4334 ;
    wire \c0.n4_adj_4332 ;
    wire \c0.n26_adj_4662 ;
    wire bfn_9_21_0_;
    wire \c0.n19795 ;
    wire \c0.n19796 ;
    wire \c0.n19797 ;
    wire \c0.n19798 ;
    wire \c0.n19799 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.n19800 ;
    wire \c0.n19801 ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.n21611 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.n21573 ;
    wire \c0.n21581 ;
    wire \c0.n21575 ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.n21577 ;
    wire n9806_cascade_;
    wire PIN_12_c;
    wire quadA_delayed_adj_4767;
    wire n9806;
    wire n14345;
    wire a_delay_counter_15__N_4123_adj_4772;
    wire n14345_cascade_;
    wire n39_adj_4770;
    wire \quad_counter1.a_delay_counter_5 ;
    wire \quad_counter1.a_delay_counter_11 ;
    wire \quad_counter1.a_delay_counter_4 ;
    wire a_delay_counter_0_adj_4765;
    wire \quad_counter1.n25 ;
    wire \quad_counter1.a_delay_counter_9 ;
    wire \quad_counter1.a_delay_counter_6 ;
    wire \quad_counter1.a_delay_counter_12 ;
    wire \quad_counter1.a_delay_counter_13 ;
    wire \quad_counter1.n26 ;
    wire \quad_counter1.a_delay_counter_8 ;
    wire \quad_counter1.a_delay_counter_1 ;
    wire \quad_counter1.a_delay_counter_2 ;
    wire \quad_counter1.a_delay_counter_3 ;
    wire \quad_counter1.n28 ;
    wire \quad_counter1.a_delay_counter_14 ;
    wire \quad_counter1.a_delay_counter_7 ;
    wire \quad_counter1.a_delay_counter_10 ;
    wire \quad_counter1.a_delay_counter_15 ;
    wire \quad_counter1.n27 ;
    wire B_filtered_adj_4764;
    wire \quad_counter1.A_delayed ;
    wire r_Tx_Data_4;
    wire \c0.n21391_cascade_ ;
    wire \c0.n21362_cascade_ ;
    wire \c0.n21244_cascade_ ;
    wire \c0.n22163 ;
    wire \c0.n6_adj_4297_cascade_ ;
    wire \c0.data_out_frame_28_4 ;
    wire n26_cascade_;
    wire n25021;
    wire n25022;
    wire \c0.n24033_cascade_ ;
    wire n21307_cascade_;
    wire \c0.n7_cascade_ ;
    wire \c0.n23918 ;
    wire r_Tx_Data_2;
    wire \c0.n20341_cascade_ ;
    wire data_out_frame_13_7;
    wire data_out_frame_10_7;
    wire n9603;
    wire byte_transmit_counter_5;
    wire r_Tx_Data_0;
    wire data_out_frame_13_6;
    wire data_out_frame_8_3;
    wire n24796;
    wire data_out_frame_7_7;
    wire n24805_cascade_;
    wire n10_adj_4780;
    wire data_out_frame_11_5;
    wire \c0.n25092_cascade_ ;
    wire \c0.n25095_cascade_ ;
    wire n25014;
    wire data_out_frame_9_5;
    wire n25008;
    wire \c0.n11_adj_4681 ;
    wire \c0.n24897 ;
    wire data_out_frame_5_0;
    wire data_out_frame_0_2;
    wire data_out_frame_12_5;
    wire \c0.n24900 ;
    wire n14247_cascade_;
    wire data_out_frame_0_3;
    wire \c0.n8_adj_4740_cascade_ ;
    wire \c0.n22952_cascade_ ;
    wire \c0.n14380 ;
    wire \c0.n14380_cascade_ ;
    wire \c0.n14942 ;
    wire \c0.n4728 ;
    wire \c0.n4728_cascade_ ;
    wire \c0.n58_adj_4742 ;
    wire \c0.n22952 ;
    wire \c0.r_SM_Main_2_N_3754_0 ;
    wire \c0.tx_active ;
    wire \c0.n5_cascade_ ;
    wire \c0.n21585 ;
    wire \c0.n3 ;
    wire \c0.n21597 ;
    wire \c0.n21587 ;
    wire \c0.n10_adj_4303_cascade_ ;
    wire \c0.data_out_frame_29__7__N_849 ;
    wire \c0.n22246_cascade_ ;
    wire \c0.n22846 ;
    wire \c0.n20379_cascade_ ;
    wire A_filtered_adj_4763;
    wire \quad_counter1.B_delayed ;
    wire \c0.n6_adj_4456 ;
    wire n21484_cascade_;
    wire \c0.n22246 ;
    wire data_out_frame_7_3;
    wire \c0.n10_adj_4313 ;
    wire data_out_frame_11_3;
    wire \c0.n22534 ;
    wire \c0.n22534_cascade_ ;
    wire \c0.n20415_cascade_ ;
    wire \c0.n20384 ;
    wire \c0.n22544 ;
    wire \c0.data_out_frame_28_5 ;
    wire \c0.n26_adj_4680 ;
    wire \c0.n22478 ;
    wire n22735;
    wire n22735_cascade_;
    wire \c0.n22757 ;
    wire \c0.n20_adj_4699_cascade_ ;
    wire n22285;
    wire \c0.n6_adj_4210 ;
    wire \c0.n13683 ;
    wire data_out_frame_10_3;
    wire \c0.n21362 ;
    wire \c0.n11_adj_4572 ;
    wire data_out_frame_13_0;
    wire data_out_frame_6_2;
    wire \c0.n5_adj_4650_cascade_ ;
    wire \c0.n6_adj_4649 ;
    wire \c0.n24953 ;
    wire \c0.n24803 ;
    wire data_out_frame_8_2;
    wire \c0.n25059_cascade_ ;
    wire n25004_cascade_;
    wire n10_adj_4778;
    wire \c0.n24809 ;
    wire n24811;
    wire n24904;
    wire data_out_frame_28_3;
    wire \c0.n25110_cascade_ ;
    wire \c0.n25113 ;
    wire \c0.n25056 ;
    wire data_out_frame_10_2;
    wire data_out_frame_11_0;
    wire \c0.n11_adj_4703 ;
    wire \c0.n24945_cascade_ ;
    wire n24682;
    wire \c0.n24797_cascade_ ;
    wire byte_transmit_counter_4;
    wire byte_transmit_counter_3;
    wire n24799_cascade_;
    wire n25012;
    wire n10_adj_4775;
    wire data_out_frame_11_6;
    wire \c0.n25098_cascade_ ;
    wire \c0.n25101 ;
    wire data_out_frame_6_5;
    wire data_out_frame_5_5;
    wire \c0.n5_adj_4679 ;
    wire \c0.n25016_cascade_ ;
    wire \c0.n24794 ;
    wire \c0.n5_adj_4700 ;
    wire \c0.n24255 ;
    wire \c0.n21583 ;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.n14530_cascade_ ;
    wire \c0.rx.n9_cascade_ ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.rx.n17531_cascade_ ;
    wire \c0.rx.n17590 ;
    wire \c0.rx.n17848 ;
    wire \c0.rx.n14 ;
    wire \c0.rx.n24697_cascade_ ;
    wire \c0.rx.n24914_cascade_ ;
    wire n14895_cascade_;
    wire n24921_cascade_;
    wire n24922;
    wire \c0.rx.n24916 ;
    wire \c0.rx.n8 ;
    wire r_Clock_Count_0;
    wire n226;
    wire bfn_11_26_0_;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n19716 ;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.n19717 ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.n19718 ;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.n19719 ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.n19720 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.n19721 ;
    wire \c0.rx.n19722 ;
    wire \c0.rx.r_Clock_Count_7 ;
    wire n14895;
    wire \c0.n21645 ;
    wire \c0.n22638_cascade_ ;
    wire \c0.n21323_cascade_ ;
    wire \c0.n14_adj_4368 ;
    wire \c0.n12488_cascade_ ;
    wire \c0.n20379 ;
    wire \c0.n13531_cascade_ ;
    wire \c0.n22294 ;
    wire \c0.n13741 ;
    wire \c0.n14_adj_4317_cascade_ ;
    wire \c0.n15_adj_4318 ;
    wire \c0.n6_adj_4330 ;
    wire \c0.n20367 ;
    wire \c0.n6_adj_4336 ;
    wire \c0.n22531 ;
    wire n25065;
    wire \c0.n13531 ;
    wire \c0.n20415 ;
    wire \c0.n22452 ;
    wire \c0.n9_adj_4562 ;
    wire \c0.n10_adj_4690_cascade_ ;
    wire \c0.n22710 ;
    wire \c0.n22710_cascade_ ;
    wire \c0.n12539 ;
    wire \c0.n21309 ;
    wire \c0.n6_adj_4683_cascade_ ;
    wire \c0.n13938 ;
    wire \c0.n12_adj_4688 ;
    wire \c0.n20360 ;
    wire \c0.n22668 ;
    wire \c0.n20360_cascade_ ;
    wire \c0.data_out_frame_29_7 ;
    wire \c0.n26_adj_4713 ;
    wire data_out_frame_7_0;
    wire \c0.n5_adj_4567 ;
    wire data_out_frame_13_1;
    wire \c0.n11_adj_4646 ;
    wire \c0.n5_adj_4644 ;
    wire \c0.n11_adj_4652 ;
    wire \c0.data_out_frame_28_2 ;
    wire \c0.n26_adj_4651 ;
    wire bfn_12_15_0_;
    wire \quad_counter1.count_direction ;
    wire n2291;
    wire \quad_counter1.n19731 ;
    wire n2290;
    wire \quad_counter1.n19732 ;
    wire n2289;
    wire \quad_counter1.n19733 ;
    wire n2288;
    wire \quad_counter1.n19734 ;
    wire n2287;
    wire \quad_counter1.n19735 ;
    wire n2286;
    wire \quad_counter1.n19736 ;
    wire n2285;
    wire \quad_counter1.n19737 ;
    wire \quad_counter1.n19738 ;
    wire n2284;
    wire bfn_12_16_0_;
    wire \quad_counter1.n19739 ;
    wire n2282;
    wire \quad_counter1.n19740 ;
    wire \quad_counter1.n19741 ;
    wire n2280;
    wire \quad_counter1.n19742 ;
    wire n2279;
    wire \quad_counter1.n19743 ;
    wire encoder1_position_13;
    wire n2278;
    wire \quad_counter1.n19744 ;
    wire n2277;
    wire \quad_counter1.n19745 ;
    wire \quad_counter1.n19746 ;
    wire n2276;
    wire bfn_12_17_0_;
    wire \quad_counter1.n19747 ;
    wire \quad_counter1.n19748 ;
    wire \quad_counter1.n19749 ;
    wire encoder1_position_19;
    wire n2272;
    wire \quad_counter1.n19750 ;
    wire n2271;
    wire \quad_counter1.n19751 ;
    wire \quad_counter1.n19752 ;
    wire n2269;
    wire \quad_counter1.n19753 ;
    wire \quad_counter1.n19754 ;
    wire bfn_12_18_0_;
    wire \quad_counter1.n19755 ;
    wire n2266;
    wire \quad_counter1.n19756 ;
    wire \quad_counter1.n19757 ;
    wire \quad_counter1.n19758 ;
    wire \quad_counter1.n19759 ;
    wire \quad_counter1.n19760 ;
    wire \quad_counter1.n19761 ;
    wire \quad_counter1.n19762 ;
    wire \quad_counter1.n2226 ;
    wire bfn_12_19_0_;
    wire \c0.n24784_cascade_ ;
    wire n25019;
    wire data_out_frame_11_2;
    wire n2273;
    wire encoder1_position_18;
    wire n2275;
    wire data_out_frame_10_0;
    wire data_out_frame_10_4;
    wire \c0.n24783 ;
    wire data_out_frame_6_0;
    wire \c0.tx_transmit_N_3650 ;
    wire \c0.n24888 ;
    wire data_out_frame_12_0;
    wire data_out_frame_12_1;
    wire data_out_frame_9_6;
    wire data_out_frame_6_6;
    wire n14247;
    wire data_out_frame_0_4;
    wire data_out_frame_9_2;
    wire data_out_frame_11_4;
    wire data_out_frame_13_2;
    wire \c0.n12976 ;
    wire \c0.n12976_cascade_ ;
    wire \c0.data_out_frame_29_7_N_1482_0_cascade_ ;
    wire \c0.n6_adj_4495 ;
    wire \c0.n14784 ;
    wire \c0.n9706_cascade_ ;
    wire \c0.n6_cascade_ ;
    wire \c0.n21579 ;
    wire \c0.n4_adj_4678 ;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n22131 ;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire \c0.n21625 ;
    wire \c0.n8_adj_4561 ;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.n8_adj_4558 ;
    wire \c0.n21637 ;
    wire \c0.n22638 ;
    wire \c0.n22831_cascade_ ;
    wire \c0.n20_adj_4321 ;
    wire \c0.n13_adj_4320_cascade_ ;
    wire \c0.n14_adj_4319 ;
    wire \c0.n28_adj_4322_cascade_ ;
    wire \c0.n12488 ;
    wire encoder1_position_14;
    wire \c0.n20318_cascade_ ;
    wire encoder1_position_16;
    wire \c0.n20449 ;
    wire \c0.n10_adj_4374 ;
    wire \c0.data_out_frame_29__7__N_855 ;
    wire \c0.n13384 ;
    wire encoder1_position_0;
    wire \c0.n22611 ;
    wire \c0.n10_adj_4274 ;
    wire \c0.n22791 ;
    wire \c0.n22466 ;
    wire \c0.n13121 ;
    wire \c0.n34_adj_4328 ;
    wire \c0.n30_adj_4326_cascade_ ;
    wire \c0.n29_adj_4329 ;
    wire encoder1_position_20;
    wire \c0.n22788 ;
    wire \c0.n22788_cascade_ ;
    wire n2274;
    wire n2283;
    wire \c0.n22656 ;
    wire \c0.n22800 ;
    wire \c0.n10_adj_4339 ;
    wire \c0.n14_adj_4338_cascade_ ;
    wire \c0.n20461_cascade_ ;
    wire \c0.n20388 ;
    wire \c0.n22408 ;
    wire \c0.n22268 ;
    wire \c0.n5_adj_4660 ;
    wire \c0.n6_adj_4659 ;
    wire \c0.n24755 ;
    wire \c0.n22330 ;
    wire \c0.n19_adj_4693_cascade_ ;
    wire \c0.n6_adj_4691_cascade_ ;
    wire \c0.n21_adj_4692 ;
    wire \c0.n21457 ;
    wire \c0.n21489 ;
    wire encoder1_position_6;
    wire \c0.n20461 ;
    wire \c0.n21330_cascade_ ;
    wire \c0.n6_adj_4331 ;
    wire \c0.n22414 ;
    wire n21307;
    wire \c0.n6_adj_4215_cascade_ ;
    wire \c0.data_out_frame_29_0 ;
    wire \c0.data_out_frame_28_0 ;
    wire \c0.n26_adj_4570 ;
    wire \c0.n10529_cascade_ ;
    wire \c0.n22489_cascade_ ;
    wire \c0.n21416_cascade_ ;
    wire \c0.n24530 ;
    wire \c0.n22671_cascade_ ;
    wire \c0.n20230 ;
    wire \c0.n20230_cascade_ ;
    wire \c0.data_out_frame_29_5 ;
    wire data_out_frame_7_1;
    wire n2270;
    wire \c0.n13395 ;
    wire encoder1_position_1;
    wire data_out_frame_9_0;
    wire data_out_frame_5_4;
    wire encoder1_position_22;
    wire encoder1_position_7;
    wire data_out_frame_7_2;
    wire encoder1_position_11;
    wire data_out_frame_12_3;
    wire data_out_frame_12_2;
    wire n2281;
    wire encoder1_position_10;
    wire data_out_frame_5_6;
    wire encoder1_position_15;
    wire data_out_frame_12_7;
    wire n2263;
    wire n2264;
    wire encoder1_position_27;
    wire data_out_frame_5_3;
    wire n2262;
    wire data_out_frame_10_6;
    wire encoder1_position_4;
    wire data_out_frame_8_0;
    wire encoder1_position_17;
    wire \c0.n16_adj_4233 ;
    wire data_out_frame_11_7;
    wire data_out_frame_13_5;
    wire data_out_frame_13_4;
    wire \c0.n11_adj_4669 ;
    wire data_out_frame_8_5;
    wire data_out_frame_7_5;
    wire encoder1_position_25;
    wire \c0.n7570_cascade_ ;
    wire data_out_frame_6_4;
    wire data_out_frame_7_4;
    wire \c0.n13055_cascade_ ;
    wire n13058_cascade_;
    wire data_out_frame_7_6;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.n5_adj_4477 ;
    wire \c0.data_out_frame_29_7_N_1482_2 ;
    wire \c0.n14_adj_4727_cascade_ ;
    wire \c0.n13056 ;
    wire \c0.n63_adj_4235 ;
    wire \c0.n63_adj_4238 ;
    wire \c0.n2004_cascade_ ;
    wire \c0.n28_adj_4565 ;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.n6_adj_4583 ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.n14_adj_4520 ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.n9_adj_4522 ;
    wire \c0.n20_adj_4265 ;
    wire \c0.n16919 ;
    wire \c0.n20_adj_4265_cascade_ ;
    wire \c0.n22148 ;
    wire \c0.n22145 ;
    wire \c0.n6_adj_4264 ;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n14721 ;
    wire \c0.n14530 ;
    wire \c0.n7_adj_4741 ;
    wire \c0.n9683 ;
    wire \c0.n9587 ;
    wire \c0.n9683_cascade_ ;
    wire \c0.n10 ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.n21653 ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.n21649 ;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.n21595 ;
    wire \c0.n21643 ;
    wire bfn_14_9_0_;
    wire encoder0_position_0;
    wire \quad_counter0.count_direction ;
    wire n2357;
    wire \quad_counter0.n19763 ;
    wire encoder0_position_1;
    wire n2356;
    wire \quad_counter0.n19764 ;
    wire n2355;
    wire \quad_counter0.n19765 ;
    wire n2354;
    wire \quad_counter0.n19766 ;
    wire n2353;
    wire \quad_counter0.n19767 ;
    wire \quad_counter0.n19768 ;
    wire n2351;
    wire \quad_counter0.n19769 ;
    wire \quad_counter0.n19770 ;
    wire encoder0_position_7;
    wire n2350;
    wire bfn_14_10_0_;
    wire \quad_counter0.n19771 ;
    wire \quad_counter0.n19772 ;
    wire encoder0_position_10;
    wire n2347;
    wire \quad_counter0.n19773 ;
    wire encoder0_position_11;
    wire n2346;
    wire \quad_counter0.n19774 ;
    wire encoder0_position_12;
    wire n2345;
    wire \quad_counter0.n19775 ;
    wire \quad_counter0.n19776 ;
    wire \quad_counter0.n19777 ;
    wire \quad_counter0.n19778 ;
    wire bfn_14_11_0_;
    wire encoder0_position_16;
    wire n2341;
    wire \quad_counter0.n19779 ;
    wire \quad_counter0.n19780 ;
    wire \quad_counter0.n19781 ;
    wire \quad_counter0.n19782 ;
    wire \quad_counter0.n19783 ;
    wire \quad_counter0.n19784 ;
    wire \quad_counter0.n19785 ;
    wire \quad_counter0.n19786 ;
    wire bfn_14_12_0_;
    wire n2333;
    wire \quad_counter0.n19787 ;
    wire n2332;
    wire \quad_counter0.n19788 ;
    wire encoder0_position_26;
    wire n2331;
    wire \quad_counter0.n19789 ;
    wire n2330;
    wire \quad_counter0.n19790 ;
    wire encoder0_position_28;
    wire n2329;
    wire \quad_counter0.n19791 ;
    wire encoder0_position_29;
    wire n2328;
    wire \quad_counter0.n19792 ;
    wire n2327;
    wire \quad_counter0.n19793 ;
    wire \quad_counter0.n19794 ;
    wire \quad_counter0.n2313 ;
    wire bfn_14_13_0_;
    wire n2326_cascade_;
    wire \c0.n22218 ;
    wire \c0.n21323 ;
    wire \c0.n22671 ;
    wire \c0.n20_adj_4694 ;
    wire \c0.n20348 ;
    wire \c0.n21330 ;
    wire \c0.n21355_cascade_ ;
    wire \c0.n12464 ;
    wire \c0.n20404 ;
    wire \c0.n20766 ;
    wire n2335;
    wire \c0.n10427 ;
    wire \c0.n21360_cascade_ ;
    wire \c0.n10504 ;
    wire \c0.n22366 ;
    wire \c0.n10504_cascade_ ;
    wire \c0.n22327 ;
    wire n21484;
    wire \c0.n28_adj_4698 ;
    wire \c0.n25_adj_4695_cascade_ ;
    wire \c0.data_out_frame_29_1 ;
    wire \c0.n22489 ;
    wire \c0.n21393 ;
    wire \c0.n22797 ;
    wire \c0.n26_adj_4697 ;
    wire \c0.n22475 ;
    wire \c0.data_out_frame_29__7__N_1143 ;
    wire \c0.n10_adj_4214 ;
    wire \c0.data_out_frame_28_1 ;
    wire \c0.n24033 ;
    wire \c0.n27_adj_4696 ;
    wire data_in_0_0;
    wire data_in_0_4;
    wire \c0.n15_adj_4242_cascade_ ;
    wire \c0.n22291 ;
    wire \c0.n20333 ;
    wire \c0.data_out_frame_29__7__N_1148 ;
    wire \c0.n21464 ;
    wire n2267;
    wire encoder1_position_24;
    wire \c0.n10_adj_4367 ;
    wire \c0.n10_adj_4239 ;
    wire \c0.n13049 ;
    wire data_in_2_4;
    wire \c0.n13049_cascade_ ;
    wire \c0.n18_adj_4236_cascade_ ;
    wire \c0.n20_adj_4237 ;
    wire data_in_1_4;
    wire \c0.n14_adj_4241 ;
    wire \c0.n17_adj_4234 ;
    wire n2268;
    wire encoder1_position_23;
    wire n2344;
    wire \c0.n10_adj_4240 ;
    wire n14374;
    wire \c0.tx.n24889 ;
    wire \c0.tx.r_Clock_Count_0 ;
    wire n2265;
    wire encoder1_position_26;
    wire data_out_frame_10_1;
    wire data_out_frame_11_1;
    wire \c0.n25116_cascade_ ;
    wire data_out_frame_9_1;
    wire \c0.n25119 ;
    wire data_in_2_2;
    wire data_out_frame_8_1;
    wire encoder1_position_29;
    wire data_out_frame_10_5;
    wire \c0.n13046 ;
    wire \c0.n12898 ;
    wire \c0.n20_adj_4308_cascade_ ;
    wire \c0.n19_adj_4307 ;
    wire \c0.n16_adj_4231_cascade_ ;
    wire \c0.n12986 ;
    wire \c0.n24745 ;
    wire data_in_2_6;
    wire data_in_0_5;
    wire \c0.n17_adj_4232 ;
    wire n2261;
    wire encoder1_position_30;
    wire data_in_3_7;
    wire data_in_3_5;
    wire \c0.n13063 ;
    wire \c0.n13063_cascade_ ;
    wire \c0.n6_adj_4263 ;
    wire \c0.n9706 ;
    wire \c0.n3325 ;
    wire data_in_2_7;
    wire data_in_1_7;
    wire \c0.n17682 ;
    wire \c0.n1 ;
    wire \c0.n17846 ;
    wire \c0.n4_adj_4654 ;
    wire \c0.n17533 ;
    wire \c0.n22907 ;
    wire \c0.n24422 ;
    wire \c0.n24596_cascade_ ;
    wire \c0.n2004 ;
    wire \c0.rx.r_SM_Main_2_N_3686_0 ;
    wire \c0.rx.n6_cascade_ ;
    wire n14439;
    wire \c0.n7570 ;
    wire \c0.n24386 ;
    wire \c0.n24302_cascade_ ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.n8_adj_4556 ;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.n21639 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n8_adj_4555 ;
    wire \c0.n21641 ;
    wire encoder0_position_30;
    wire n2342;
    wire encoder0_position_15;
    wire n2352;
    wire \c0.n30_adj_4730_cascade_ ;
    wire \c0.n17539 ;
    wire \c0.n22372 ;
    wire encoder1_position_28;
    wire \c0.n31_adj_4325 ;
    wire \c0.n22775 ;
    wire n2348;
    wire n2336;
    wire \c0.n22608 ;
    wire encoder0_position_2;
    wire \c0.n22785 ;
    wire \c0.n13630 ;
    wire n2340;
    wire \c0.byte_transmit_counter_2 ;
    wire \c0.n5_adj_4217 ;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n24901 ;
    wire \c0.n25062 ;
    wire n2260;
    wire count_enable_adj_4769;
    wire encoder1_position_31;
    wire n2338;
    wire encoder1_position_21;
    wire encoder0_position_17;
    wire encoder1_position_8;
    wire \c0.n22593 ;
    wire encoder1_position_9;
    wire \c0.n6_adj_4276 ;
    wire \c0.n21441 ;
    wire encoder0_position_25;
    wire data_out_frame_6_1;
    wire data_out_frame_29_2;
    wire \c0.n12_adj_4312 ;
    wire \c0.n24113_cascade_ ;
    wire \c0.n10529 ;
    wire encoder1_position_5;
    wire \c0.n21364 ;
    wire \c0.n24113 ;
    wire \c0.n21311_cascade_ ;
    wire \c0.n21244 ;
    wire \c0.n21496 ;
    wire \c0.n21273_cascade_ ;
    wire \c0.data_out_frame_29_6 ;
    wire \c0.data_out_frame_28_6 ;
    wire \c0.n26_adj_4702 ;
    wire \c0.n22617 ;
    wire \c0.n20341 ;
    wire \c0.n18_adj_4684_cascade_ ;
    wire \c0.n13268 ;
    wire \c0.n15_adj_4686 ;
    wire \c0.n20_adj_4685_cascade_ ;
    wire \c0.n21475 ;
    wire \c0.data_out_frame_28_7 ;
    wire \c0.n22461 ;
    wire \c0.n21358 ;
    wire \c0.n22461_cascade_ ;
    wire \c0.n21406 ;
    wire \c0.n24028 ;
    wire \c0.n14_adj_4478_cascade_ ;
    wire \c0.n22193 ;
    wire \c0.n13422 ;
    wire \c0.n22722 ;
    wire data_out_frame_29__2__N_1748;
    wire \c0.n19_adj_4720 ;
    wire data_in_2_1;
    wire data_out_frame_29_3;
    wire encoder1_position_12;
    wire data_out_frame_12_4;
    wire data_in_0_3;
    wire \c0.n15 ;
    wire data_in_3_4;
    wire n2334;
    wire data_in_1_0;
    wire n2349;
    wire \c0.rx.r_SM_Main_2_N_3680_2 ;
    wire encoder0_position_19;
    wire \c0.n22199_cascade_ ;
    wire \c0.n22834 ;
    wire encoder0_position_13;
    wire encoder0_position_22;
    wire \c0.n6_adj_4366 ;
    wire data_in_2_0;
    wire \c0.n22635 ;
    wire \c0.n22256_cascade_ ;
    wire \c0.n22772 ;
    wire data_in_1_3;
    wire control_mode_4;
    wire \c0.byte_transmit_counter_0 ;
    wire data_out_frame_9_4;
    wire data_out_frame_8_4;
    wire \c0.n24782 ;
    wire encoder0_position_8;
    wire \c0.n22423 ;
    wire encoder0_position_6;
    wire \c0.n6_adj_4293 ;
    wire encoder0_position_23;
    wire encoder0_position_9;
    wire control_mode_7;
    wire \c0.n22385_cascade_ ;
    wire encoder0_position_24;
    wire \c0.n20325 ;
    wire data_in_2_5;
    wire data_in_1_5;
    wire control_mode_6;
    wire data_in_1_1;
    wire data_in_0_1;
    wire data_in_3_2;
    wire \c0.n74_adj_4525 ;
    wire \c0.n4_adj_4212 ;
    wire \c0.n22098_cascade_ ;
    wire \c0.n4_adj_4306 ;
    wire \c0.n63_adj_4305_cascade_ ;
    wire \c0.n13001 ;
    wire \c0.FRAME_MATCHER_state_0 ;
    wire \c0.n9248 ;
    wire \c0.n13055 ;
    wire \c0.data_out_frame_29_7_N_1482_0 ;
    wire data_out_frame_29_7_N_2878_2;
    wire \c0.n9_adj_4549 ;
    wire n63;
    wire \c0.n3844 ;
    wire \c0.n58_adj_4706 ;
    wire \c0.n24591_cascade_ ;
    wire \c0.n6_adj_4728 ;
    wire \c0.FRAME_MATCHER_state_2 ;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.n21659 ;
    wire \c0.n4_adj_4721 ;
    wire \c0.n937 ;
    wire \c0.data_out_frame_29_7_N_1482_1 ;
    wire \c0.FRAME_MATCHER_state_1 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire \c0.n8_adj_4553 ;
    wire data_in_1_6;
    wire data_in_0_6;
    wire data_in_3_6;
    wire \c0.n20_adj_4726 ;
    wire \c0.n27_adj_4735 ;
    wire \c0.data_out_frame_29__7__N_735 ;
    wire \c0.n13665 ;
    wire \c0.n22754 ;
    wire \c0.n13558 ;
    wire \c0.n22754_cascade_ ;
    wire \c0.n22243 ;
    wire \c0.n22580 ;
    wire \c0.n10477 ;
    wire n2339;
    wire encoder0_position_18;
    wire \c0.n22583 ;
    wire \c0.n22149 ;
    wire encoder0_position_3;
    wire \c0.n22583_cascade_ ;
    wire encoder0_position_31;
    wire \c0.n13872 ;
    wire n2337;
    wire n17571;
    wire encoder0_position_21;
    wire \c0.n22252 ;
    wire encoder0_position_27;
    wire data_out_frame_6_3;
    wire encoder1_position_3;
    wire \c0.n20455 ;
    wire encoder0_position_5;
    wire encoder0_position_20;
    wire \c0.n22689 ;
    wire \c0.n22641 ;
    wire encoder0_position_4;
    wire \c0.n22689_cascade_ ;
    wire control_mode_0;
    wire \c0.n10455 ;
    wire \c0.n20312 ;
    wire \c0.n20312_cascade_ ;
    wire \c0.n22522 ;
    wire \c0.n6_adj_4674_cascade_ ;
    wire \c0.data_out_frame_29_4 ;
    wire \c0.n8162 ;
    wire \c0.n21355 ;
    wire \c0.n12604 ;
    wire \c0.n20786 ;
    wire \c0.n20786_cascade_ ;
    wire \c0.n9_adj_4494 ;
    wire \c0.n10497 ;
    wire \c0.n21433 ;
    wire \c0.n21311 ;
    wire \c0.n12590 ;
    wire \c0.n21399 ;
    wire \c0.n22553 ;
    wire encoder1_position_2;
    wire \c0.n21416 ;
    wire \c0.n10531 ;
    wire \c0.n20511 ;
    wire \c0.n10531_cascade_ ;
    wire \c0.n21451 ;
    wire \c0.n21437 ;
    wire \c0.n21451_cascade_ ;
    wire n13058;
    wire data_out_frame_8_6;
    wire \c0.n10467 ;
    wire \c0.n10500 ;
    wire \c0.n21349 ;
    wire \c0.n4_adj_4271 ;
    wire \c0.data_out_frame_29__6__N_1538 ;
    wire \c0.n21327 ;
    wire \c0.n4_adj_4271_cascade_ ;
    wire \c0.data_out_frame_29__3__N_1730 ;
    wire data_out_frame_29__3__N_1661;
    wire \c0.rx.n12909 ;
    wire \c0.n22112_cascade_ ;
    wire data_in_2_3;
    wire \c0.n82_cascade_ ;
    wire r_Bit_Index_0;
    wire \c0.rx.n17834_cascade_ ;
    wire n14484;
    wire n14988;
    wire control_mode_5;
    wire control_mode_1;
    wire control_mode_3;
    wire count_enable;
    wire n2343;
    wire encoder0_position_14;
    wire n4_adj_4761;
    wire \c0.data_in_frame_29_3 ;
    wire \c0.n17_adj_4483 ;
    wire \c0.n26_adj_4480_cascade_ ;
    wire \c0.n63_adj_4249 ;
    wire \c0.n34_adj_4546_cascade_ ;
    wire n24622;
    wire n24622_cascade_;
    wire control_mode_2;
    wire \c0.n24539 ;
    wire \c0.n24733 ;
    wire \c0.n18_adj_4485 ;
    wire \c0.n22134_cascade_ ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n21633 ;
    wire \c0.n6 ;
    wire \c0.n4_adj_4266 ;
    wire \c0.n5024 ;
    wire \c0.n12992 ;
    wire \c0.n13052 ;
    wire \c0.n24736 ;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n21651 ;
    wire FRAME_MATCHER_state_31_N_2975_2;
    wire \c0.n22_adj_4643_cascade_ ;
    wire \c0.n10_adj_4639_cascade_ ;
    wire \c0.n13_adj_4640 ;
    wire \c0.n20_adj_4642 ;
    wire \c0.n14_adj_4607_cascade_ ;
    wire \c0.n22626 ;
    wire \c0.data_out_frame_0__7__N_2626_cascade_ ;
    wire \c0.n30_adj_4585 ;
    wire \c0.n6_adj_4254_cascade_ ;
    wire \c0.n28_adj_4731 ;
    wire data_in_3_3;
    wire data_in_0_7;
    wire \c0.n14 ;
    wire \c0.n20_adj_4729 ;
    wire \c0.n6_adj_4704 ;
    wire \c0.n14016_cascade_ ;
    wire \c0.n20_cascade_ ;
    wire data_in_frame_5_6;
    wire \c0.data_in_frame_7_7 ;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n21629 ;
    wire \c0.n25_adj_4723 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n22049 ;
    wire \c0.n5 ;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.n21647 ;
    wire data_in_1_2;
    wire data_in_0_2;
    wire \c0.n10_adj_4732 ;
    wire \c0.n26_adj_4733_cascade_ ;
    wire \c0.n20409_cascade_ ;
    wire \c0.n22716_cascade_ ;
    wire \c0.n8_adj_4248 ;
    wire data_in_3_1;
    wire data_in_3_0;
    wire n12981;
    wire n4_adj_4762;
    wire \c0.n22716 ;
    wire \c0.n5_adj_4302 ;
    wire \c0.n12_adj_4348_cascade_ ;
    wire \c0.n8_adj_4526 ;
    wire \c0.n8_adj_4526_cascade_ ;
    wire \c0.n9_adj_4536 ;
    wire \c0.n14_adj_4528 ;
    wire \c0.n14_adj_4576 ;
    wire \c0.data_in_frame_29_5 ;
    wire \c0.n24098_cascade_ ;
    wire \c0.n10_adj_4484 ;
    wire \c0.n52_cascade_ ;
    wire \c0.n47_adj_4537_cascade_ ;
    wire \c0.n24581 ;
    wire \c0.data_in_frame_29_1 ;
    wire \c0.data_in_frame_29_6 ;
    wire \c0.n20793 ;
    wire \c0.n20793_cascade_ ;
    wire \c0.n12927 ;
    wire \c0.n39_adj_4295 ;
    wire \c0.n13043 ;
    wire \c0.n23912 ;
    wire \c0.n35 ;
    wire \c0.n22885 ;
    wire r_Bit_Index_2;
    wire r_Bit_Index_1;
    wire n4;
    wire r_Rx_Data;
    wire n4_cascade_;
    wire n12904;
    wire \c0.rx.n14277 ;
    wire \c0.n12514 ;
    wire \c0.n20641 ;
    wire \c0.n21391 ;
    wire \c0.n21360 ;
    wire \c0.n21_adj_4719 ;
    wire rx_data_ready;
    wire \c0.FRAME_MATCHER_rx_data_ready_prev ;
    wire r_SM_Main_1;
    wire \c0.rx.r_SM_Main_0 ;
    wire r_SM_Main_2;
    wire \c0.rx.n22094 ;
    wire \c0.n46_adj_4739 ;
    wire \c0.n39_adj_4737 ;
    wire \c0.n38_adj_4736 ;
    wire \c0.n23562 ;
    wire \c0.n23562_cascade_ ;
    wire data_in_frame_5_5;
    wire \c0.data_in_frame_3_4 ;
    wire \c0.n12_adj_4657 ;
    wire \c0.n23_adj_4648 ;
    wire \c0.n38_adj_4285_cascade_ ;
    wire \c0.n26_adj_4289 ;
    wire \c0.n26_adj_4289_cascade_ ;
    wire \c0.data_out_frame_0__7__N_2626 ;
    wire \c0.n20_adj_4290 ;
    wire \c0.n20_adj_4290_cascade_ ;
    wire data_in_frame_1_1;
    wire \c0.n51 ;
    wire \c0.n29 ;
    wire \c0.n51_cascade_ ;
    wire \c0.n22_adj_4647 ;
    wire \c0.n102_cascade_ ;
    wire \c0.n32 ;
    wire \c0.n16_adj_4256_cascade_ ;
    wire \c0.n9_adj_4279 ;
    wire \c0.n13141 ;
    wire \c0.n9_adj_4279_cascade_ ;
    wire \c0.n23574_cascade_ ;
    wire \c0.n11_adj_4257 ;
    wire \c0.n7_adj_4337 ;
    wire \c0.n38_adj_4573_cascade_ ;
    wire \c0.n44_adj_4744 ;
    wire \c0.n43_adj_4574_cascade_ ;
    wire \c0.n41_adj_4745 ;
    wire \c0.n24048 ;
    wire \c0.n24048_cascade_ ;
    wire \c0.n109 ;
    wire \c0.n23_adj_4590 ;
    wire \c0.n29_adj_4734 ;
    wire \c0.n7_adj_4221 ;
    wire \c0.n16_adj_4641 ;
    wire \c0.n23116_cascade_ ;
    wire \c0.n23116 ;
    wire \c0.n128 ;
    wire \c0.n129_cascade_ ;
    wire \c0.n11_adj_4614 ;
    wire \c0.n16_adj_4613_cascade_ ;
    wire data_in_frame_1_3;
    wire \c0.n126 ;
    wire \c0.n123 ;
    wire \c0.n144_cascade_ ;
    wire \c0.n154 ;
    wire \c0.n15_adj_4301 ;
    wire \c0.n21_adj_4605 ;
    wire \c0.n19_adj_4604 ;
    wire \c0.n16_adj_4256 ;
    wire \c0.n22 ;
    wire \c0.n13280 ;
    wire \c0.n13_cascade_ ;
    wire \c0.n20_adj_4222 ;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.n22_adj_4223_cascade_ ;
    wire \c0.n21_adj_4225_cascade_ ;
    wire \c0.n10_adj_4277_cascade_ ;
    wire \c0.n10_adj_4591_cascade_ ;
    wire \c0.n10_adj_4591 ;
    wire data_in_frame_21_2;
    wire \c0.n12_adj_4606_cascade_ ;
    wire \c0.n21325_cascade_ ;
    wire \c0.n24384 ;
    wire \c0.n4_adj_4464_cascade_ ;
    wire \c0.n21428_cascade_ ;
    wire \c0.n24_adj_4593 ;
    wire \c0.n23_adj_4598 ;
    wire \c0.n4_adj_4352 ;
    wire \c0.n23_adj_4353 ;
    wire \c0.n23_adj_4353_cascade_ ;
    wire \c0.n15_adj_4344 ;
    wire \c0.n21428 ;
    wire \c0.n11_adj_4438_cascade_ ;
    wire \c0.n16_adj_4437 ;
    wire \c0.n22420 ;
    wire \c0.data_in_frame_28_0 ;
    wire \c0.n21491 ;
    wire \c0.n23187_cascade_ ;
    wire \c0.n10_adj_4439_cascade_ ;
    wire \c0.n20_adj_4441 ;
    wire \c0.n13_adj_4442_cascade_ ;
    wire \c0.n24528_cascade_ ;
    wire \c0.n23718 ;
    wire \c0.n12_adj_4506 ;
    wire \c0.n20_adj_4512 ;
    wire \c0.n24_adj_4509 ;
    wire \c0.n22_adj_4507 ;
    wire \c0.n23627 ;
    wire \c0.n23627_cascade_ ;
    wire \c0.n24528 ;
    wire \c0.n10_adj_4575 ;
    wire \c0.data_in_frame_24_7 ;
    wire \c0.n25467 ;
    wire \c0.n24098 ;
    wire \c0.data_in_frame_29_4 ;
    wire \c0.n23533 ;
    wire \c0.n5_adj_4370 ;
    wire \c0.n10_adj_4371 ;
    wire \c0.n5_adj_4349 ;
    wire \c0.n10_adj_4371_cascade_ ;
    wire \c0.n12_adj_4372 ;
    wire \c0.n12_adj_4671_cascade_ ;
    wire \c0.data_in_frame_28_7 ;
    wire \c0.n45_adj_4298 ;
    wire \c0.data_in_frame_25_3 ;
    wire \c0.data_in_frame_25_2 ;
    wire \c0.n40_adj_4294 ;
    wire \c0.n41_adj_4292 ;
    wire \c0.n42_adj_4272_cascade_ ;
    wire \c0.n44_adj_4270 ;
    wire \c0.n50_adj_4296 ;
    wire \c0.n43_adj_4275 ;
    wire \c0.n161 ;
    wire bfn_19_1_0_;
    wire \c0.n19625 ;
    wire \c0.n19625_THRU_CRY_0_THRU_CO ;
    wire \c0.n19625_THRU_CRY_1_THRU_CO ;
    wire \c0.n19625_THRU_CRY_2_THRU_CO ;
    wire \c0.n19625_THRU_CRY_3_THRU_CO ;
    wire \c0.n19625_THRU_CRY_4_THRU_CO ;
    wire \c0.n19625_THRU_CRY_5_THRU_CO ;
    wire \c0.n19625_THRU_CRY_6_THRU_CO ;
    wire bfn_19_2_0_;
    wire \c0.n3_adj_4434 ;
    wire \c0.n19626 ;
    wire \c0.n19626_THRU_CRY_0_THRU_CO ;
    wire \c0.n19626_THRU_CRY_1_THRU_CO ;
    wire \c0.n19626_THRU_CRY_2_THRU_CO ;
    wire \c0.n19626_THRU_CRY_3_THRU_CO ;
    wire \c0.n19626_THRU_CRY_4_THRU_CO ;
    wire \c0.n19626_THRU_CRY_5_THRU_CO ;
    wire \c0.n19626_THRU_CRY_6_THRU_CO ;
    wire bfn_19_3_0_;
    wire \c0.n3_adj_4432 ;
    wire \c0.n19627 ;
    wire \c0.n19627_THRU_CRY_0_THRU_CO ;
    wire \c0.n19627_THRU_CRY_1_THRU_CO ;
    wire \c0.n19627_THRU_CRY_2_THRU_CO ;
    wire \c0.n19627_THRU_CRY_3_THRU_CO ;
    wire \c0.n19627_THRU_CRY_4_THRU_CO ;
    wire \c0.n19627_THRU_CRY_5_THRU_CO ;
    wire \c0.n19627_THRU_CRY_6_THRU_CO ;
    wire bfn_19_4_0_;
    wire \c0.n19628 ;
    wire \c0.n19628_THRU_CRY_0_THRU_CO ;
    wire \c0.n19628_THRU_CRY_1_THRU_CO ;
    wire \c0.n19628_THRU_CRY_2_THRU_CO ;
    wire \c0.n19628_THRU_CRY_3_THRU_CO ;
    wire \c0.n19628_THRU_CRY_4_THRU_CO ;
    wire \c0.n19628_THRU_CRY_5_THRU_CO ;
    wire \c0.n19628_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire bfn_19_5_0_;
    wire \c0.n3_adj_4428 ;
    wire \c0.n19629 ;
    wire \c0.n19629_THRU_CRY_0_THRU_CO ;
    wire \c0.n19629_THRU_CRY_1_THRU_CO ;
    wire \c0.n19629_THRU_CRY_2_THRU_CO ;
    wire \c0.n19629_THRU_CRY_3_THRU_CO ;
    wire \c0.n19629_THRU_CRY_4_THRU_CO ;
    wire \c0.n19629_THRU_CRY_5_THRU_CO ;
    wire \c0.n19629_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire bfn_19_6_0_;
    wire \c0.n3_adj_4426 ;
    wire \c0.n19630 ;
    wire \c0.n19630_THRU_CRY_0_THRU_CO ;
    wire \c0.n19630_THRU_CRY_1_THRU_CO ;
    wire \c0.n19630_THRU_CRY_2_THRU_CO ;
    wire \c0.n19630_THRU_CRY_3_THRU_CO ;
    wire \c0.n19630_THRU_CRY_4_THRU_CO ;
    wire \c0.n19630_THRU_CRY_5_THRU_CO ;
    wire \c0.n19630_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire bfn_19_7_0_;
    wire \c0.n3_adj_4424 ;
    wire \c0.n19631 ;
    wire \c0.n19631_THRU_CRY_0_THRU_CO ;
    wire \c0.n19631_THRU_CRY_1_THRU_CO ;
    wire \c0.n19631_THRU_CRY_2_THRU_CO ;
    wire \c0.n19631_THRU_CRY_3_THRU_CO ;
    wire \c0.n19631_THRU_CRY_4_THRU_CO ;
    wire \c0.n19631_THRU_CRY_5_THRU_CO ;
    wire \c0.n19631_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire bfn_19_8_0_;
    wire \c0.n3_adj_4422 ;
    wire \c0.n19632 ;
    wire \c0.n19632_THRU_CRY_0_THRU_CO ;
    wire \c0.n19632_THRU_CRY_1_THRU_CO ;
    wire \c0.n19632_THRU_CRY_2_THRU_CO ;
    wire \c0.n19632_THRU_CRY_3_THRU_CO ;
    wire \c0.n19632_THRU_CRY_4_THRU_CO ;
    wire \c0.n19632_THRU_CRY_5_THRU_CO ;
    wire \c0.n19632_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire bfn_19_9_0_;
    wire \c0.n3_adj_4420 ;
    wire \c0.n19633 ;
    wire \c0.n19633_THRU_CRY_0_THRU_CO ;
    wire \c0.n19633_THRU_CRY_1_THRU_CO ;
    wire \c0.n19633_THRU_CRY_2_THRU_CO ;
    wire \c0.n19633_THRU_CRY_3_THRU_CO ;
    wire \c0.n19633_THRU_CRY_4_THRU_CO ;
    wire \c0.n19633_THRU_CRY_5_THRU_CO ;
    wire \c0.n19633_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire bfn_19_10_0_;
    wire \c0.n3_adj_4418 ;
    wire \c0.n19634 ;
    wire \c0.n19634_THRU_CRY_0_THRU_CO ;
    wire \c0.n19634_THRU_CRY_1_THRU_CO ;
    wire \c0.n19634_THRU_CRY_2_THRU_CO ;
    wire \c0.n19634_THRU_CRY_3_THRU_CO ;
    wire \c0.n19634_THRU_CRY_4_THRU_CO ;
    wire \c0.n19634_THRU_CRY_5_THRU_CO ;
    wire \c0.n19634_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire bfn_19_11_0_;
    wire \c0.n3_adj_4416 ;
    wire \c0.n19635 ;
    wire \c0.n19635_THRU_CRY_0_THRU_CO ;
    wire \c0.n19635_THRU_CRY_1_THRU_CO ;
    wire \c0.n19635_THRU_CRY_2_THRU_CO ;
    wire \c0.n19635_THRU_CRY_3_THRU_CO ;
    wire \c0.n19635_THRU_CRY_4_THRU_CO ;
    wire \c0.n19635_THRU_CRY_5_THRU_CO ;
    wire \c0.n19635_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire bfn_19_12_0_;
    wire \c0.n3_adj_4414 ;
    wire \c0.n19636 ;
    wire \c0.n19636_THRU_CRY_0_THRU_CO ;
    wire \c0.n19636_THRU_CRY_1_THRU_CO ;
    wire \c0.n19636_THRU_CRY_2_THRU_CO ;
    wire \c0.n19636_THRU_CRY_3_THRU_CO ;
    wire \c0.n19636_THRU_CRY_4_THRU_CO ;
    wire \c0.n19636_THRU_CRY_5_THRU_CO ;
    wire \c0.n19636_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire bfn_19_13_0_;
    wire \c0.n3_adj_4412 ;
    wire \c0.n19637 ;
    wire \c0.n19637_THRU_CRY_0_THRU_CO ;
    wire \c0.n19637_THRU_CRY_1_THRU_CO ;
    wire \c0.n19637_THRU_CRY_2_THRU_CO ;
    wire \c0.n19637_THRU_CRY_3_THRU_CO ;
    wire \c0.n19637_THRU_CRY_4_THRU_CO ;
    wire \c0.n19637_THRU_CRY_5_THRU_CO ;
    wire \c0.n19637_THRU_CRY_6_THRU_CO ;
    wire bfn_19_14_0_;
    wire \c0.n19638 ;
    wire \c0.n19638_THRU_CRY_0_THRU_CO ;
    wire \c0.n19638_THRU_CRY_1_THRU_CO ;
    wire \c0.n19638_THRU_CRY_2_THRU_CO ;
    wire \c0.n19638_THRU_CRY_3_THRU_CO ;
    wire \c0.n19638_THRU_CRY_4_THRU_CO ;
    wire \c0.n19638_THRU_CRY_5_THRU_CO ;
    wire \c0.n19638_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire bfn_19_15_0_;
    wire \c0.n3_adj_4408 ;
    wire \c0.n19639 ;
    wire \c0.n19639_THRU_CRY_0_THRU_CO ;
    wire \c0.n19639_THRU_CRY_1_THRU_CO ;
    wire \c0.n19639_THRU_CRY_2_THRU_CO ;
    wire \c0.n19639_THRU_CRY_3_THRU_CO ;
    wire \c0.n19639_THRU_CRY_4_THRU_CO ;
    wire \c0.n19639_THRU_CRY_5_THRU_CO ;
    wire \c0.n19639_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire bfn_19_16_0_;
    wire \c0.n3_adj_4406 ;
    wire \c0.n19640 ;
    wire \c0.n19640_THRU_CRY_0_THRU_CO ;
    wire \c0.n19640_THRU_CRY_1_THRU_CO ;
    wire \c0.n19640_THRU_CRY_2_THRU_CO ;
    wire \c0.n19640_THRU_CRY_3_THRU_CO ;
    wire \c0.n19640_THRU_CRY_4_THRU_CO ;
    wire \c0.n19640_THRU_CRY_5_THRU_CO ;
    wire \c0.n19640_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire bfn_19_17_0_;
    wire \c0.n3_adj_4404 ;
    wire \c0.n19641 ;
    wire \c0.n19641_THRU_CRY_0_THRU_CO ;
    wire \c0.n19641_THRU_CRY_1_THRU_CO ;
    wire \c0.n19641_THRU_CRY_2_THRU_CO ;
    wire \c0.n19641_THRU_CRY_3_THRU_CO ;
    wire \c0.n19641_THRU_CRY_4_THRU_CO ;
    wire \c0.n19641_THRU_CRY_5_THRU_CO ;
    wire \c0.n19641_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire bfn_19_18_0_;
    wire \c0.n3_adj_4402 ;
    wire \c0.n19642 ;
    wire \c0.n19642_THRU_CRY_0_THRU_CO ;
    wire \c0.n19642_THRU_CRY_1_THRU_CO ;
    wire \c0.n19642_THRU_CRY_2_THRU_CO ;
    wire \c0.n19642_THRU_CRY_3_THRU_CO ;
    wire \c0.n19642_THRU_CRY_4_THRU_CO ;
    wire \c0.n19642_THRU_CRY_5_THRU_CO ;
    wire \c0.n19642_THRU_CRY_6_THRU_CO ;
    wire bfn_19_19_0_;
    wire \c0.n19643 ;
    wire \c0.n19643_THRU_CRY_0_THRU_CO ;
    wire \c0.n19643_THRU_CRY_1_THRU_CO ;
    wire \c0.n19643_THRU_CRY_2_THRU_CO ;
    wire \c0.n19643_THRU_CRY_3_THRU_CO ;
    wire \c0.n19643_THRU_CRY_4_THRU_CO ;
    wire \c0.n19643_THRU_CRY_5_THRU_CO ;
    wire \c0.n19643_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire bfn_19_20_0_;
    wire \c0.n3_adj_4398 ;
    wire \c0.n19644 ;
    wire \c0.n19644_THRU_CRY_0_THRU_CO ;
    wire \c0.n19644_THRU_CRY_1_THRU_CO ;
    wire \c0.n19644_THRU_CRY_2_THRU_CO ;
    wire \c0.n19644_THRU_CRY_3_THRU_CO ;
    wire \c0.n19644_THRU_CRY_4_THRU_CO ;
    wire \c0.n19644_THRU_CRY_5_THRU_CO ;
    wire \c0.n19644_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire bfn_19_21_0_;
    wire \c0.n3_adj_4396 ;
    wire \c0.n19645 ;
    wire \c0.n19645_THRU_CRY_0_THRU_CO ;
    wire \c0.n19645_THRU_CRY_1_THRU_CO ;
    wire \c0.n19645_THRU_CRY_2_THRU_CO ;
    wire \c0.n19645_THRU_CRY_3_THRU_CO ;
    wire \c0.n19645_THRU_CRY_4_THRU_CO ;
    wire \c0.n19645_THRU_CRY_5_THRU_CO ;
    wire \c0.n19645_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire bfn_19_22_0_;
    wire \c0.n3_adj_4394 ;
    wire \c0.n19646 ;
    wire \c0.n19646_THRU_CRY_0_THRU_CO ;
    wire \c0.n19646_THRU_CRY_1_THRU_CO ;
    wire \c0.n19646_THRU_CRY_2_THRU_CO ;
    wire \c0.n19646_THRU_CRY_3_THRU_CO ;
    wire \c0.n19646_THRU_CRY_4_THRU_CO ;
    wire \c0.n19646_THRU_CRY_5_THRU_CO ;
    wire \c0.n19646_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire bfn_19_23_0_;
    wire \c0.n3_adj_4392 ;
    wire \c0.n19647 ;
    wire \c0.n19647_THRU_CRY_0_THRU_CO ;
    wire \c0.n19647_THRU_CRY_1_THRU_CO ;
    wire \c0.n19647_THRU_CRY_2_THRU_CO ;
    wire \c0.n19647_THRU_CRY_3_THRU_CO ;
    wire \c0.n19647_THRU_CRY_4_THRU_CO ;
    wire \c0.n19647_THRU_CRY_5_THRU_CO ;
    wire \c0.n19647_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire bfn_19_24_0_;
    wire \c0.n3_adj_4390 ;
    wire \c0.n19648 ;
    wire \c0.n19648_THRU_CRY_0_THRU_CO ;
    wire \c0.n19648_THRU_CRY_1_THRU_CO ;
    wire \c0.n19648_THRU_CRY_2_THRU_CO ;
    wire \c0.n19648_THRU_CRY_3_THRU_CO ;
    wire \c0.n19648_THRU_CRY_4_THRU_CO ;
    wire \c0.n19648_THRU_CRY_5_THRU_CO ;
    wire \c0.n19648_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire bfn_19_25_0_;
    wire \c0.n3_adj_4388 ;
    wire \c0.n19649 ;
    wire \c0.n19649_THRU_CRY_0_THRU_CO ;
    wire \c0.n19649_THRU_CRY_1_THRU_CO ;
    wire \c0.n19649_THRU_CRY_2_THRU_CO ;
    wire \c0.n19649_THRU_CRY_3_THRU_CO ;
    wire \c0.n19649_THRU_CRY_4_THRU_CO ;
    wire \c0.n19649_THRU_CRY_5_THRU_CO ;
    wire \c0.n19649_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire bfn_19_26_0_;
    wire \c0.n3_adj_4386 ;
    wire \c0.n19650 ;
    wire \c0.n19650_THRU_CRY_0_THRU_CO ;
    wire \c0.n19650_THRU_CRY_1_THRU_CO ;
    wire \c0.n19650_THRU_CRY_2_THRU_CO ;
    wire \c0.n19650_THRU_CRY_3_THRU_CO ;
    wire \c0.n19650_THRU_CRY_4_THRU_CO ;
    wire \c0.n19650_THRU_CRY_5_THRU_CO ;
    wire \c0.n19650_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire bfn_19_27_0_;
    wire \c0.n3_adj_4384 ;
    wire \c0.n19651 ;
    wire \c0.n19651_THRU_CRY_0_THRU_CO ;
    wire \c0.n19651_THRU_CRY_1_THRU_CO ;
    wire \c0.n19651_THRU_CRY_2_THRU_CO ;
    wire \c0.n19651_THRU_CRY_3_THRU_CO ;
    wire \c0.n19651_THRU_CRY_4_THRU_CO ;
    wire \c0.n19651_THRU_CRY_5_THRU_CO ;
    wire \c0.n19651_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire bfn_19_28_0_;
    wire \c0.n3_adj_4382 ;
    wire \c0.n19652 ;
    wire \c0.n19652_THRU_CRY_0_THRU_CO ;
    wire \c0.n19652_THRU_CRY_1_THRU_CO ;
    wire \c0.n19652_THRU_CRY_2_THRU_CO ;
    wire \c0.n19652_THRU_CRY_3_THRU_CO ;
    wire \c0.n19652_THRU_CRY_4_THRU_CO ;
    wire \c0.n19652_THRU_CRY_5_THRU_CO ;
    wire \c0.n19652_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire bfn_19_29_0_;
    wire \c0.n3_adj_4380 ;
    wire \c0.n19653 ;
    wire \c0.n19653_THRU_CRY_0_THRU_CO ;
    wire \c0.n19653_THRU_CRY_1_THRU_CO ;
    wire \c0.n19653_THRU_CRY_2_THRU_CO ;
    wire \c0.n19653_THRU_CRY_3_THRU_CO ;
    wire \c0.n19653_THRU_CRY_4_THRU_CO ;
    wire \c0.n19653_THRU_CRY_5_THRU_CO ;
    wire \c0.n19653_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire bfn_19_30_0_;
    wire \c0.n3_adj_4378 ;
    wire \c0.n19654 ;
    wire \c0.n19654_THRU_CRY_0_THRU_CO ;
    wire \c0.n19654_THRU_CRY_1_THRU_CO ;
    wire \c0.n19654_THRU_CRY_2_THRU_CO ;
    wire \c0.n19654_THRU_CRY_3_THRU_CO ;
    wire \c0.n19654_THRU_CRY_4_THRU_CO ;
    wire \c0.n19654_THRU_CRY_5_THRU_CO ;
    wire \c0.n19654_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire bfn_19_31_0_;
    wire \c0.n3_adj_4376 ;
    wire \c0.n19655 ;
    wire \c0.n19655_THRU_CRY_0_THRU_CO ;
    wire \c0.n19655_THRU_CRY_1_THRU_CO ;
    wire \c0.n19655_THRU_CRY_2_THRU_CO ;
    wire \c0.n19655_THRU_CRY_3_THRU_CO ;
    wire \c0.n19655_THRU_CRY_4_THRU_CO ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \c0.n19655_THRU_CRY_5_THRU_CO ;
    wire \c0.n19655_THRU_CRY_6_THRU_CO ;
    wire bfn_19_32_0_;
    wire \c0.FRAME_MATCHER_i_31 ;
    wire \c0.n3_adj_4373 ;
    wire \c0.n17856 ;
    wire \c0.n1306 ;
    wire \c0.n3_adj_4436 ;
    wire \c0.n22196_cascade_ ;
    wire \c0.n12_adj_4258 ;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.n10_adj_4615 ;
    wire \c0.data_in_frame_3_1 ;
    wire \c0.n7_adj_4300 ;
    wire \c0.n12_adj_4299 ;
    wire \c0.n7_adj_4300_cascade_ ;
    wire \c0.n11_adj_4280 ;
    wire \c0.n23251 ;
    wire \c0.n23305 ;
    wire \c0.n23251_cascade_ ;
    wire \c0.n23574 ;
    wire \c0.n7_adj_4282_cascade_ ;
    wire \c0.n10_adj_4283 ;
    wire \c0.data_in_frame_8_1 ;
    wire \c0.n13_adj_4638_cascade_ ;
    wire \c0.data_in_frame_10_1 ;
    wire \c0.data_in_frame_10_2 ;
    wire \c0.data_in_frame_9_7 ;
    wire \c0.n5_adj_4268 ;
    wire \c0.n4_adj_4267 ;
    wire \c0.n4_adj_4269 ;
    wire \c0.n22196 ;
    wire \c0.n4_adj_4269_cascade_ ;
    wire \c0.n68 ;
    wire \c0.n89_cascade_ ;
    wire \c0.n23_cascade_ ;
    wire \c0.n26 ;
    wire \c0.n13075_cascade_ ;
    wire \c0.n93_cascade_ ;
    wire data_in_frame_14_1;
    wire \c0.n102 ;
    wire \c0.n147_cascade_ ;
    wire \c0.n134 ;
    wire \c0.n131 ;
    wire \c0.n31_adj_4284 ;
    wire \c0.n36_adj_4447 ;
    wire \c0.n41_adj_4452_cascade_ ;
    wire \c0.data_in_frame_11_7 ;
    wire \c0.n39_adj_4453 ;
    wire \c0.n40_adj_4451 ;
    wire \c0.n14016 ;
    wire \c0.n13223 ;
    wire \c0.n16_adj_4608 ;
    wire \c0.n21 ;
    wire \c0.n20 ;
    wire \c0.n13_adj_4610 ;
    wire \c0.data_in_frame_4_1 ;
    wire \c0.data_in_frame_10_4 ;
    wire \c0.n22455 ;
    wire \c0.data_in_frame_12_5 ;
    wire \c0.n42 ;
    wire \c0.n58 ;
    wire \c0.n127 ;
    wire \c0.n5_adj_4311 ;
    wire \c0.n5_adj_4311_cascade_ ;
    wire \c0.data_in_frame_10_3 ;
    wire \c0.n23677 ;
    wire data_in_frame_14_4;
    wire \c0.data_in_frame_8_2 ;
    wire \c0.n120_cascade_ ;
    wire \c0.n142 ;
    wire \c0.n152_cascade_ ;
    wire \c0.n158 ;
    wire \c0.n22472 ;
    wire data_in_frame_14_3;
    wire \c0.n30_adj_4571_cascade_ ;
    wire \c0.n33 ;
    wire \c0.n34_adj_4600_cascade_ ;
    wire \c0.n38_adj_4573 ;
    wire \c0.n24333_cascade_ ;
    wire \c0.n23661 ;
    wire \c0.data_in_frame_18_5 ;
    wire \c0.data_in_frame_16_3 ;
    wire \c0.n155 ;
    wire \c0.n160 ;
    wire \c0.n12989 ;
    wire \c0.n22104_cascade_ ;
    wire \c0.data_in_frame_19_4 ;
    wire \c0.n22347_cascade_ ;
    wire \c0.n24520 ;
    wire \c0.data_in_frame_20_5 ;
    wire \c0.n22_adj_4350 ;
    wire \c0.n22_adj_4350_cascade_ ;
    wire \c0.data_in_frame_20_6 ;
    wire \c0.data_in_frame_20_7 ;
    wire \c0.n21_adj_4225 ;
    wire \c0.n22227 ;
    wire \c0.n23863 ;
    wire \c0.n9_adj_4521 ;
    wire \c0.n20_adj_4596 ;
    wire \c0.n23733_cascade_ ;
    wire \c0.data_in_frame_26_0 ;
    wire \c0.data_in_frame_27_7 ;
    wire \c0.n20314_cascade_ ;
    wire \c0.n21325 ;
    wire \c0.n20314 ;
    wire \c0.n22_adj_4597 ;
    wire \c0.n12_adj_4671 ;
    wire \c0.data_in_frame_29_7 ;
    wire \c0.data_in_frame_27_5 ;
    wire \c0.data_in_frame_27_6 ;
    wire \c0.data_in_frame_25_5 ;
    wire \c0.n12_adj_4466 ;
    wire \c0.n11_adj_4474_cascade_ ;
    wire \c0.n21280 ;
    wire \c0.data_in_frame_29_2 ;
    wire \c0.n25446 ;
    wire \c0.data_in_frame_29_0 ;
    wire \c0.n10874 ;
    wire \c0.n43_adj_4463_cascade_ ;
    wire \c0.n21389 ;
    wire \c0.data_in_frame_25_0 ;
    wire \c0.n64_adj_4539 ;
    wire \c0.n10_adj_4544 ;
    wire \c0.n13911 ;
    wire \c0.n23921_cascade_ ;
    wire \c0.n21_adj_4547 ;
    wire \c0.n23975 ;
    wire \c0.n32_adj_4533 ;
    wire \c0.n74 ;
    wire \c0.n70_adj_4514 ;
    wire \c0.n71_cascade_ ;
    wire \c0.n17537 ;
    wire \c0.n81_cascade_ ;
    wire \c0.n82_adj_4517 ;
    wire \c0.n28_adj_4523 ;
    wire \c0.data_in_frame_27_3 ;
    wire \c0.data_in_frame_27_4 ;
    wire \c0.n23_adj_4532_cascade_ ;
    wire \c0.n31_adj_4542 ;
    wire \c0.n38_adj_4535_cascade_ ;
    wire \c0.n32_adj_4534 ;
    wire \c0.n8_adj_4677 ;
    wire \c0.data_in_frame_9_6 ;
    wire data_in_frame_5_3;
    wire data_in_frame_5_2;
    wire \c0.data_in_frame_7_6 ;
    wire data_in_frame_1_2;
    wire \c0.n12_adj_4612 ;
    wire \c0.n15_adj_4444 ;
    wire \c0.n15_adj_4444_cascade_ ;
    wire \c0.n11_adj_4656 ;
    wire \c0.data_in_frame_3_2 ;
    wire data_in_frame_5_4;
    wire \c0.n6_adj_4611 ;
    wire \c0.n6_adj_4611_cascade_ ;
    wire \c0.n91 ;
    wire \c0.n13453 ;
    wire \c0.n13_adj_4584 ;
    wire \c0.n102_adj_4445 ;
    wire \c0.n101 ;
    wire \c0.n103 ;
    wire \c0.n98 ;
    wire \c0.n97 ;
    wire \c0.n110_cascade_ ;
    wire \c0.n24465 ;
    wire \c0.data_out_frame_0__7__N_2579 ;
    wire \c0.n15_adj_4450 ;
    wire \c0.n87 ;
    wire \c0.n85 ;
    wire \c0.n88 ;
    wire \c0.n87_cascade_ ;
    wire \c0.n106 ;
    wire \c0.n22160 ;
    wire \c0.n7_adj_4304 ;
    wire \c0.n7_adj_4304_cascade_ ;
    wire data_in_frame_5_7;
    wire data_in_frame_6_0;
    wire \c0.n27_adj_4725 ;
    wire \c0.n17_adj_4224 ;
    wire \c0.n130 ;
    wire \c0.n14_adj_4707 ;
    wire \c0.n15_adj_4710 ;
    wire \c0.n22511 ;
    wire \c0.n22_adj_4259 ;
    wire data_in_frame_6_1;
    wire \c0.n18_adj_4314_cascade_ ;
    wire \c0.data_in_frame_3_7 ;
    wire data_in_frame_1_6;
    wire \c0.n38_adj_4448 ;
    wire \c0.n42_adj_4449 ;
    wire \c0.data_in_frame_3_3 ;
    wire \c0.n24_adj_4689 ;
    wire \c0.n13_adj_4281 ;
    wire \c0.n31 ;
    wire \c0.n31_cascade_ ;
    wire \c0.data_in_frame_10_0 ;
    wire \c0.n28 ;
    wire \c0.n24 ;
    wire \c0.n16 ;
    wire data_in_frame_14_2;
    wire \c0.n8_adj_4673 ;
    wire data_in_frame_6_2;
    wire \c0.data_in_frame_13_0 ;
    wire \c0.n22205_cascade_ ;
    wire \c0.n23491 ;
    wire \c0.n23598_cascade_ ;
    wire \c0.n23611 ;
    wire \c0.n9_adj_4208_cascade_ ;
    wire \c0.n22304 ;
    wire \c0.n13892_cascade_ ;
    wire \c0.data_in_frame_11_6 ;
    wire \c0.n13892 ;
    wire \c0.data_in_frame_17_2 ;
    wire \c0.n22_adj_4622 ;
    wire \c0.n22825_cascade_ ;
    wire data_in_frame_14_0;
    wire \c0.n136 ;
    wire \c0.n22751_cascade_ ;
    wire \c0.n107 ;
    wire \c0.n149 ;
    wire \c0.n140 ;
    wire \c0.n22843 ;
    wire \c0.n22_adj_4245 ;
    wire \c0.n22514_cascade_ ;
    wire \c0.data_in_frame_16_1 ;
    wire \c0.n14_adj_4566 ;
    wire \c0.n14165_cascade_ ;
    wire \c0.data_in_frame_12_4 ;
    wire \c0.n4_adj_4658_cascade_ ;
    wire \c0.n24433 ;
    wire \c0.data_in_frame_16_6 ;
    wire \c0.n12_adj_4682_cascade_ ;
    wire \c0.n23390 ;
    wire \c0.n22249 ;
    wire \c0.n10_adj_4315 ;
    wire \c0.n24534 ;
    wire \c0.data_in_frame_17_3 ;
    wire \c0.n4_adj_4345 ;
    wire \c0.n24534_cascade_ ;
    wire \c0.n12_adj_4346 ;
    wire \c0.n13329 ;
    wire \c0.n4_adj_4621 ;
    wire \c0.n12_adj_4500 ;
    wire \c0.n9_adj_4208 ;
    wire \c0.n6_adj_4587_cascade_ ;
    wire \c0.n13461 ;
    wire \c0.n13756 ;
    wire \c0.n13461_cascade_ ;
    wire \c0.n6227_cascade_ ;
    wire \c0.n22173 ;
    wire \c0.n19_adj_4291 ;
    wire data_in_frame_14_6;
    wire n22118;
    wire \c0.data_in_frame_19_3 ;
    wire \c0.n14088 ;
    wire \c0.n23300 ;
    wire \c0.n6_adj_4577 ;
    wire \c0.n22662 ;
    wire \c0.n23300_cascade_ ;
    wire \c0.n21_adj_4594 ;
    wire \c0.n4_adj_4347 ;
    wire \c0.data_in_frame_23_4 ;
    wire \c0.n4_adj_4347_cascade_ ;
    wire \c0.data_in_frame_23_1 ;
    wire \c0.n30_adj_4357_cascade_ ;
    wire \c0.n14_adj_4356 ;
    wire \c0.n40_adj_4359 ;
    wire \c0.n42_adj_4358_cascade_ ;
    wire \c0.n41_adj_4360 ;
    wire \c0.n37_adj_4458 ;
    wire \c0.n34_adj_4361_cascade_ ;
    wire \c0.n14148 ;
    wire \c0.data_in_frame_20_4 ;
    wire \c0.n30_adj_4357 ;
    wire \c0.n22334 ;
    wire \c0.data_in_frame_25_6 ;
    wire \c0.data_in_frame_24_3 ;
    wire \c0.n24547 ;
    wire \c0.n21353 ;
    wire \c0.n66_cascade_ ;
    wire \c0.n75 ;
    wire \c0.n46_adj_4461 ;
    wire \c0.n10_adj_4513 ;
    wire \c0.n15_adj_4497 ;
    wire \c0.data_in_frame_25_4 ;
    wire \c0.n23_adj_4551 ;
    wire \c0.n26_adj_4548 ;
    wire \c0.n24_adj_4550_cascade_ ;
    wire \c0.n21010_cascade_ ;
    wire \c0.n53_adj_4538 ;
    wire \c0.n61_adj_4543 ;
    wire \c0.n42_adj_4540 ;
    wire \c0.n62_adj_4541 ;
    wire \c0.n13_adj_4492 ;
    wire \c0.n18_adj_4493 ;
    wire \c0.n22_adj_4498 ;
    wire \c0.n26_adj_4499_cascade_ ;
    wire \c0.n24441_cascade_ ;
    wire \c0.n30_adj_4545 ;
    wire \c0.n72 ;
    wire \c0.n24559 ;
    wire \c0.n42_adj_4510 ;
    wire \c0.n20_adj_4518 ;
    wire \c0.n24751 ;
    wire \c0.n14_adj_4676_cascade_ ;
    wire \c0.data_out_frame_0__7__N_2777 ;
    wire \c0.data_in_frame_0_6 ;
    wire \c0.n24016 ;
    wire \c0.n24749 ;
    wire data_in_frame_1_4;
    wire data_in_frame_1_5;
    wire \c0.n37_adj_4738 ;
    wire \c0.data_in_frame_0_5 ;
    wire \c0.data_in_frame_0_7 ;
    wire \c0.n22316 ;
    wire \c0.n23554 ;
    wire \c0.n34_cascade_ ;
    wire \c0.n23655 ;
    wire \c0.n53 ;
    wire \c0.n54_cascade_ ;
    wire \c0.n56 ;
    wire \c0.n13821 ;
    wire \c0.n48 ;
    wire \c0.n37_cascade_ ;
    wire \c0.n22647_cascade_ ;
    wire \c0.data_in_frame_2_6 ;
    wire \c0.n24747 ;
    wire \c0.n10_adj_4722 ;
    wire \c0.n14_adj_4616_cascade_ ;
    wire \c0.n23666 ;
    wire \c0.n37 ;
    wire \c0.n55 ;
    wire \c0.n18_adj_4314 ;
    wire \c0.n24_adj_4724 ;
    wire data_in_frame_1_0;
    wire \c0.n5_adj_4711 ;
    wire \c0.n16_adj_4716 ;
    wire \c0.n28_adj_4718_cascade_ ;
    wire \c0.n24_adj_4717 ;
    wire \c0.n23_adj_4599 ;
    wire \c0.n4_adj_4446 ;
    wire \c0.n4_adj_4446_cascade_ ;
    wire \c0.n26_adj_4714 ;
    wire \c0.data_in_frame_4_0 ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.n23597 ;
    wire \c0.data_in_frame_2_0 ;
    wire \c0.n22230 ;
    wire \c0.data_in_frame_9_4 ;
    wire \c0.n150 ;
    wire \c0.n13651 ;
    wire \c0.n18_adj_4228 ;
    wire \c0.n27_cascade_ ;
    wire \c0.n19 ;
    wire \c0.n23528_cascade_ ;
    wire \c0.n34_adj_4278_cascade_ ;
    wire \c0.n36 ;
    wire \c0.n48_adj_4227 ;
    wire \c0.n30_adj_4705_cascade_ ;
    wire \c0.n23523_cascade_ ;
    wire \c0.n30 ;
    wire \c0.n13075 ;
    wire \c0.n7_adj_4634_cascade_ ;
    wire \c0.data_in_frame_10_5 ;
    wire \c0.n96_cascade_ ;
    wire \c0.data_in_frame_8_0 ;
    wire \c0.n104 ;
    wire \c0.n7_adj_4253 ;
    wire \c0.n5_adj_4252 ;
    wire \c0.n5_adj_4443 ;
    wire \c0.n13734_cascade_ ;
    wire \c0.n17734 ;
    wire \c0.n12973 ;
    wire \c0.n13128 ;
    wire \c0.n7_adj_4603 ;
    wire \c0.n22589 ;
    wire \c0.n13738_cascade_ ;
    wire \c0.data_in_frame_10_6 ;
    wire \c0.data_in_frame_10_7 ;
    wire \c0.n13734 ;
    wire \c0.n39_adj_4708_cascade_ ;
    wire \c0.n63 ;
    wire \c0.n64_cascade_ ;
    wire \c0.n13721 ;
    wire \c0.n55_adj_4709 ;
    wire \c0.n13186 ;
    wire \c0.n124 ;
    wire \c0.n10_adj_4247 ;
    wire \c0.n22547 ;
    wire \c0.n13998 ;
    wire \c0.n23156 ;
    wire \c0.n65 ;
    wire \c0.n60 ;
    wire \c0.n59_cascade_ ;
    wire \c0.n70 ;
    wire \c0.n24444_cascade_ ;
    wire \c0.n21282 ;
    wire \c0.data_in_frame_15_7 ;
    wire \c0.n22514 ;
    wire \c0.n23224_cascade_ ;
    wire \c0.n21409 ;
    wire \c0.data_in_frame_18_6 ;
    wire \c0.n22540 ;
    wire \c0.n24333 ;
    wire \c0.n22822 ;
    wire data_in_frame_14_7;
    wire \c0.n12_adj_4246_cascade_ ;
    wire \c0.n23691_cascade_ ;
    wire \c0.n20543 ;
    wire \c0.data_in_frame_16_5 ;
    wire \c0.n10_adj_4602 ;
    wire \c0.n22644 ;
    wire \c0.data_in_frame_15_1 ;
    wire \c0.n14165 ;
    wire data_in_frame_14_5;
    wire \c0.n24444 ;
    wire \c0.n7_adj_4581 ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire \c0.n3_adj_4430 ;
    wire \c0.n20467 ;
    wire \c0.n20467_cascade_ ;
    wire \c0.n6404 ;
    wire \c0.n17_adj_4354_cascade_ ;
    wire \c0.n10_adj_4630 ;
    wire \c0.n23523 ;
    wire \c0.n6_adj_4209 ;
    wire \c0.data_in_frame_13_7 ;
    wire \c0.data_in_frame_12_6 ;
    wire \c0.n22782 ;
    wire \c0.n12_adj_4246 ;
    wire \c0.n23453 ;
    wire \c0.data_in_frame_12_7 ;
    wire \c0.n25_adj_4579 ;
    wire \c0.n25_adj_4579_cascade_ ;
    wire \c0.n23433_cascade_ ;
    wire \c0.n18_adj_4580 ;
    wire \c0.n24_adj_4655 ;
    wire \c0.n41_adj_4592 ;
    wire \c0.n43_adj_4661 ;
    wire \c0.n44_adj_4588 ;
    wire \c0.n39_adj_4341 ;
    wire \c0.n22205 ;
    wire \c0.n50_adj_4340_cascade_ ;
    wire \c0.n5_adj_4486 ;
    wire \c0.n12559_cascade_ ;
    wire \c0.n22375 ;
    wire \c0.n24451 ;
    wire \c0.data_in_frame_19_1 ;
    wire \c0.n6215 ;
    wire \c0.data_in_frame_19_2 ;
    wire \c0.n21275 ;
    wire \c0.n21275_cascade_ ;
    wire \c0.n14_adj_4440 ;
    wire \c0.n63_adj_4516 ;
    wire \c0.n14189 ;
    wire \c0.n46 ;
    wire \c0.n46_cascade_ ;
    wire \c0.n34_adj_4361 ;
    wire \c0.n57_cascade_ ;
    wire \c0.n48_adj_4365 ;
    wire \c0.n21426_cascade_ ;
    wire \c0.n23032 ;
    wire \c0.n23032_cascade_ ;
    wire \c0.n25456 ;
    wire \c0.n23209_cascade_ ;
    wire \c0.n56_adj_4479 ;
    wire \c0.n21299 ;
    wire data_in_frame_22_6;
    wire data_in_frame_22_0;
    wire \c0.data_in_frame_23_7 ;
    wire \c0.n7_adj_4364_cascade_ ;
    wire \c0.n21426 ;
    wire \c0.n23031_cascade_ ;
    wire \c0.data_in_frame_25_7 ;
    wire \c0.data_in_frame_26_5 ;
    wire \c0.n24482 ;
    wire \c0.n23031 ;
    wire \c0.data_in_frame_28_2 ;
    wire \c0.n36_adj_4460_cascade_ ;
    wire \c0.n41_adj_4511 ;
    wire \c0.n6_adj_4459 ;
    wire \c0.n22426 ;
    wire \c0.data_in_frame_26_1 ;
    wire \c0.n22340 ;
    wire \c0.n5_adj_4472_cascade_ ;
    wire \c0.n21010 ;
    wire \c0.n24_adj_4496 ;
    wire \c0.data_in_frame_24_1 ;
    wire \c0.data_in_frame_27_1 ;
    wire \c0.n39_adj_4515 ;
    wire \c0.n10_adj_4675 ;
    wire \c0.data_in_frame_11_0 ;
    wire \c0.data_in_frame_4_6 ;
    wire \c0.n4_adj_4211 ;
    wire \c0.n22647 ;
    wire \c0.n13904_cascade_ ;
    wire \c0.n21_adj_4327 ;
    wire \c0.n19_adj_4324_cascade_ ;
    wire \c0.n22417 ;
    wire \c0.data_in_frame_7_5 ;
    wire \c0.n22417_cascade_ ;
    wire \c0.n4_adj_4333 ;
    wire \c0.n86 ;
    wire \c0.n13085 ;
    wire \c0.n7_adj_4282 ;
    wire \c0.n50 ;
    wire n22121_cascade_;
    wire data_in_frame_6_6;
    wire \c0.data_in_frame_2_2 ;
    wire data_in_frame_6_7;
    wire \c0.data_in_frame_4_7 ;
    wire \c0.data_in_frame_2_7 ;
    wire \c0.n49 ;
    wire \c0.n23528 ;
    wire \c0.n7_adj_4229 ;
    wire \c0.data_out_frame_0__7__N_2743 ;
    wire \c0.n13523 ;
    wire \c0.n47 ;
    wire \c0.n10_adj_4664 ;
    wire \c0.data_in_frame_9_2 ;
    wire \c0.data_in_frame_7_0 ;
    wire \c0.n23406 ;
    wire data_in_frame_6_4;
    wire \c0.n14_adj_4609_cascade_ ;
    wire \c0.n10_adj_4617 ;
    wire \c0.n17 ;
    wire \c0.n8_adj_4216 ;
    wire \c0.n12_cascade_ ;
    wire \c0.data_in_frame_4_2 ;
    wire \c0.data_in_frame_12_2 ;
    wire \c0.n13809 ;
    wire \c0.data_in_frame_11_5 ;
    wire \c0.n22751 ;
    wire \c0.n23_adj_4665 ;
    wire \c0.data_in_frame_15_2 ;
    wire \c0.data_in_frame_8_5 ;
    wire \c0.data_in_frame_11_1 ;
    wire \c0.n22176 ;
    wire \c0.n28_adj_4637_cascade_ ;
    wire \c0.n24_adj_4636 ;
    wire \c0.n7_adj_4634 ;
    wire \c0.n16_adj_4635 ;
    wire \c0.data_in_frame_4_5 ;
    wire \c0.n23283 ;
    wire \c0.data_in_frame_8_7 ;
    wire \c0.n20_adj_4260 ;
    wire \c0.n22803 ;
    wire \c0.n4_adj_4261 ;
    wire \c0.n31_adj_4743 ;
    wire \c0.n5813 ;
    wire \c0.n22602 ;
    wire \c0.n11 ;
    wire \c0.n17_adj_4219 ;
    wire \c0.n16_adj_4218_cascade_ ;
    wire \c0.n13767_cascade_ ;
    wire \c0.n5965 ;
    wire \c0.n6_adj_4454 ;
    wire \c0.data_in_frame_15_3 ;
    wire \c0.n12_adj_4455 ;
    wire \c0.n22463 ;
    wire \c0.n24540 ;
    wire \c0.n23507 ;
    wire data_in_frame_21_0;
    wire \c0.data_in_frame_17_0 ;
    wire \c0.n23313 ;
    wire \c0.n26_adj_4578 ;
    wire \c0.data_in_frame_13_5 ;
    wire \c0.data_in_frame_17_7 ;
    wire \c0.data_in_frame_16_2 ;
    wire \c0.n24527 ;
    wire data_in_frame_21_3;
    wire \c0.n21344 ;
    wire \c0.n42_adj_4589 ;
    wire \c0.n22_adj_4243 ;
    wire \c0.n13738 ;
    wire \c0.n10_adj_4230 ;
    wire \c0.n5_adj_4310 ;
    wire \c0.n13604 ;
    wire \c0.n7_adj_4251_cascade_ ;
    wire \c0.n23224 ;
    wire \c0.n7_adj_4251 ;
    wire data_in_frame_22_7;
    wire \c0.n22825 ;
    wire \c0.data_in_frame_15_4 ;
    wire \c0.data_in_frame_18_2 ;
    wire \c0.data_in_frame_18_4 ;
    wire \c0.data_in_frame_18_3 ;
    wire \c0.n5_adj_4335 ;
    wire \c0.n4_adj_4568 ;
    wire \c0.n15_adj_4569 ;
    wire \c0.data_in_frame_18_7 ;
    wire data_in_frame_22_5;
    wire \c0.data_in_frame_17_5 ;
    wire \c0.n22748 ;
    wire \c0.n14_adj_4623_cascade_ ;
    wire \c0.n15_adj_4624 ;
    wire data_in_frame_21_1;
    wire \c0.n13963_cascade_ ;
    wire \c0.n22508 ;
    wire \c0.n40_adj_4342 ;
    wire \c0.data_in_frame_24_6 ;
    wire \c0.n22495 ;
    wire \c0.data_in_frame_20_1 ;
    wire \c0.n58_adj_4355 ;
    wire \c0.n59_adj_4351 ;
    wire \c0.n28_adj_4363 ;
    wire \c0.n23691 ;
    wire \c0.n22577 ;
    wire \c0.n21414 ;
    wire \c0.n10_adj_4524_cascade_ ;
    wire \c0.n13797 ;
    wire \c0.n24576 ;
    wire \c0.data_in_frame_26_2 ;
    wire \c0.n24576_cascade_ ;
    wire \c0.n14_adj_4519 ;
    wire data_in_frame_21_4;
    wire \c0.n23733 ;
    wire \c0.n22686 ;
    wire \c0.n5_adj_4472 ;
    wire \c0.n22686_cascade_ ;
    wire \c0.n21316 ;
    wire \c0.n39_adj_4487 ;
    wire \c0.n30_adj_4489_cascade_ ;
    wire \c0.n23209 ;
    wire \c0.n45_adj_4490_cascade_ ;
    wire \c0.n44_adj_4501 ;
    wire \c0.n11_adj_4505 ;
    wire \c0.n48_adj_4503_cascade_ ;
    wire \c0.n28_adj_4504 ;
    wire \c0.n24573 ;
    wire \c0.n41_adj_4488 ;
    wire \c0.n17_adj_4354 ;
    wire \c0.n28_adj_4343 ;
    wire \c0.n27_adj_4502 ;
    wire \c0.data_in_frame_26_7 ;
    wire \c0.data_in_frame_24_4 ;
    wire data_in_frame_21_6;
    wire \c0.n21301 ;
    wire \c0.n23_adj_4582 ;
    wire \c0.data_in_frame_27_2 ;
    wire \c0.n25_adj_4469 ;
    wire \c0.n26_adj_4470 ;
    wire \c0.n39_adj_4467 ;
    wire \c0.n38_adj_4468 ;
    wire \c0.n37_adj_4473 ;
    wire \c0.n44_adj_4471_cascade_ ;
    wire \c0.n45_adj_4476 ;
    wire \c0.n14_adj_4529 ;
    wire \c0.n15_adj_4508 ;
    wire \c0.n24362_cascade_ ;
    wire \c0.n18_adj_4475 ;
    wire \c0.n26_adj_4530 ;
    wire n22103;
    wire \c0.n22632 ;
    wire \c0.n22632_cascade_ ;
    wire \c0.data_in_frame_24_2 ;
    wire \c0.data_in_frame_26_3 ;
    wire \c0.n22362_cascade_ ;
    wire \c0.n12559 ;
    wire \c0.n13_adj_4527 ;
    wire \c0.n20802 ;
    wire \c0.n20358 ;
    wire \c0.n12_adj_4491 ;
    wire \c0.data_in_frame_28_6 ;
    wire \c0.data_in_frame_28_4 ;
    wire \c0.n13904 ;
    wire \c0.n28_adj_4286 ;
    wire data_in_frame_5_0;
    wire \c0.n23302 ;
    wire \c0.data_in_frame_0_3 ;
    wire \c0.data_in_frame_2_4 ;
    wire \c0.n42_adj_4746 ;
    wire \c0.data_in_frame_7_1 ;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.data_in_frame_4_3 ;
    wire \c0.n6_adj_4687_cascade_ ;
    wire \c0.n23274 ;
    wire \c0.n23282 ;
    wire \c0.n23274_cascade_ ;
    wire \c0.n20_adj_4316 ;
    wire \c0.n29_adj_4287 ;
    wire \c0.data_in_frame_0_2 ;
    wire \c0.data_in_frame_2_3 ;
    wire \c0.data_in_frame_0_1 ;
    wire \c0.data_in_frame_4_4 ;
    wire \c0.n23276 ;
    wire \c0.n22322 ;
    wire \c0.n23276_cascade_ ;
    wire \c0.n25 ;
    wire \c0.n24_adj_4213 ;
    wire \c0.n8_cascade_ ;
    wire \c0.data_in_frame_0_4 ;
    wire n22121;
    wire \c0.data_in_frame_0_0 ;
    wire \c0.n22701 ;
    wire \c0.n5_adj_4323 ;
    wire n22101;
    wire \c0.n9_cascade_ ;
    wire \c0.data_in_frame_9_1 ;
    wire \c0.data_in_frame_8_6 ;
    wire \c0.data_in_frame_18_0 ;
    wire data_in_frame_6_5;
    wire \c0.n19_adj_4620 ;
    wire \c0.n9 ;
    wire \c0.n22392 ;
    wire \c0.data_in_frame_9_5 ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire \c0.n3_adj_4410 ;
    wire \c0.data_in_frame_7_4 ;
    wire data_in_frame_5_1;
    wire \c0.n40_adj_4288 ;
    wire \c0.n22120 ;
    wire \c0.data_in_frame_7_3 ;
    wire \c0.data_in_frame_12_0 ;
    wire \c0.data_in_frame_12_1 ;
    wire \c0.n39 ;
    wire \c0.n61 ;
    wire \c0.n13253 ;
    wire \c0.n13253_cascade_ ;
    wire \c0.n22518 ;
    wire \c0.n22828 ;
    wire \c0.data_in_frame_11_4 ;
    wire \c0.data_in_frame_7_2 ;
    wire \c0.n9_adj_4220 ;
    wire \c0.n7_adj_4226 ;
    wire \c0.n27_adj_4748 ;
    wire \c0.data_in_frame_11_3 ;
    wire \c0.data_in_frame_9_0 ;
    wire \c0.n4 ;
    wire \c0.data_in_frame_28_3 ;
    wire \c0.data_in_frame_12_3 ;
    wire \c0.data_in_frame_15_6 ;
    wire \c0.n22379 ;
    wire \c0.n6_adj_4559 ;
    wire \c0.data_in_frame_17_6 ;
    wire \c0.data_in_frame_15_5 ;
    wire \c0.n31_adj_4701 ;
    wire \c0.n13474 ;
    wire \c0.n22650 ;
    wire data_in_frame_1_7;
    wire \c0.n30_adj_4747 ;
    wire \c0.n6_adj_4632 ;
    wire \c0.n5_adj_4631 ;
    wire \c0.n23343 ;
    wire \c0.n25_adj_4633 ;
    wire \c0.data_in_frame_9_3 ;
    wire \c0.data_in_frame_11_2 ;
    wire \c0.data_in_frame_28_1 ;
    wire \c0.data_in_frame_8_3 ;
    wire \c0.data_in_frame_17_4 ;
    wire \c0.data_in_frame_13_3 ;
    wire \c0.n22319 ;
    wire \c0.n4_adj_4586 ;
    wire \c0.data_in_frame_16_0 ;
    wire \c0.data_in_frame_13_6 ;
    wire \c0.data_in_frame_18_1 ;
    wire \c0.n14081 ;
    wire \c0.n10_adj_4250 ;
    wire \c0.data_in_frame_16_4 ;
    wire rx_data_4;
    wire \c0.data_in_frame_13_4 ;
    wire \c0.data_in_frame_19_5 ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire \c0.n2119 ;
    wire \c0.n3_adj_4400 ;
    wire \c0.n22112 ;
    wire \c0.data_in_frame_15_0 ;
    wire rx_data_6;
    wire data_in_frame_22_1;
    wire \c0.data_in_frame_20_2 ;
    wire \c0.data_in_frame_23_5 ;
    wire \c0.n9_adj_4563 ;
    wire \c0.data_in_frame_16_7 ;
    wire \c0.n22_adj_4244 ;
    wire \c0.n24_adj_4618 ;
    wire \c0.n14_adj_4619 ;
    wire \c0.data_in_frame_2_1 ;
    wire \c0.n22288 ;
    wire \c0.data_in_frame_13_2 ;
    wire \c0.n22288_cascade_ ;
    wire \c0.n5807 ;
    wire \c0.n14160 ;
    wire \c0.data_in_frame_17_1 ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire \c0.FRAME_MATCHER_i_0 ;
    wire \c0.n9_adj_4601 ;
    wire \c0.data_in_frame_25_1 ;
    wire \c0.data_in_frame_20_0 ;
    wire \c0.data_in_frame_19_0 ;
    wire \c0.n12_adj_4564 ;
    wire \c0.n21404 ;
    wire \c0.n6_adj_4462_cascade_ ;
    wire \c0.n22562 ;
    wire data_in_frame_22_3;
    wire \c0.data_in_frame_26_6 ;
    wire \c0.n22769 ;
    wire data_in_frame_21_5;
    wire \c0.n22698 ;
    wire \c0.data_in_frame_23_6 ;
    wire \c0.n4_adj_4464 ;
    wire \c0.n14_adj_4465 ;
    wire \c0.data_in_frame_20_3 ;
    wire \c0.n21412 ;
    wire \c0.n4_adj_4369 ;
    wire \c0.data_in_frame_27_0 ;
    wire \c0.n73 ;
    wire \c0.n20409 ;
    wire data_in_frame_22_4;
    wire \c0.n12_adj_4672 ;
    wire \c0.n22099 ;
    wire rx_data_1;
    wire \c0.data_in_frame_13_1 ;
    wire \c0.n13490 ;
    wire \c0.data_in_frame_24_5 ;
    wire \c0.n22505 ;
    wire \c0.n6718 ;
    wire \c0.n13963 ;
    wire \c0.n21295 ;
    wire \c0.n20239 ;
    wire \c0.n13468 ;
    wire \c0.n20239_cascade_ ;
    wire \c0.data_in_frame_26_4 ;
    wire \c0.n10_adj_4457 ;
    wire \c0.n6_adj_4668 ;
    wire \c0.data_in_frame_23_2 ;
    wire \c0.n13314 ;
    wire \c0.n6227 ;
    wire data_in_frame_21_7;
    wire \c0.n20350 ;
    wire rx_data_3;
    wire \c0.data_in_frame_23_3 ;
    wire \c0.n25484 ;
    wire \c0.n62 ;
    wire \c0.n21_adj_4481 ;
    wire \c0.n6_adj_4462 ;
    wire \c0.n30_adj_4482 ;
    wire \c0.n9_adj_4273 ;
    wire rx_data_7;
    wire \c0.n23598 ;
    wire \c0.data_in_frame_8_4 ;
    wire data_in_frame_6_3;
    wire \c0.n23267 ;
    wire \c0.n18_cascade_ ;
    wire \c0.n16_adj_4666 ;
    wire \c0.n28_adj_4667 ;
    wire \c0.n24_adj_4653_cascade_ ;
    wire \c0.n22369 ;
    wire \c0.n6_adj_4587 ;
    wire \c0.n22586 ;
    wire \c0.data_in_frame_19_6 ;
    wire \c0.data_in_frame_19_7 ;
    wire \c0.n23433 ;
    wire \c0.n15_adj_4625 ;
    wire \c0.n17_adj_4626 ;
    wire \c0.n16_adj_4627 ;
    wire \c0.n15_adj_4625_cascade_ ;
    wire \c0.n18 ;
    wire \c0.n22605 ;
    wire \c0.n13767 ;
    wire \c0.n19_adj_4595 ;
    wire \c0.n24_adj_4628 ;
    wire \c0.n14_adj_4629_cascade_ ;
    wire \c0.n23178 ;
    wire \c0.n22234 ;
    wire \c0.n17830 ;
    wire rx_data_0;
    wire \c0.n22104 ;
    wire \c0.data_in_frame_23_0 ;
    wire \c0.n9_adj_4552 ;
    wire rx_data_5;
    wire \c0.n22134 ;
    wire \c0.data_in_frame_28_5 ;
    wire rx_data_2;
    wire n22110;
    wire data_in_frame_22_2;
    wire CLK_c;
    wire \c0.data_in_frame_24_0 ;
    wire \c0.n29_adj_4362 ;
    wire \c0.n24_adj_4531 ;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__81286),
            .DIN(N__81285),
            .DOUT(N__81284),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__81286),
            .PADOUT(N__81285),
            .PADIN(N__81284),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26751),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_12_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_12_pad_iopad (
            .OE(N__81277),
            .DIN(N__81276),
            .DOUT(N__81275),
            .PACKAGEPIN(PIN_12));
    defparam PIN_12_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_12_pad_preio (
            .PADOEN(N__81277),
            .PADOUT(N__81276),
            .PADIN(N__81275),
            .CLOCKENABLE(),
            .DIN0(PIN_12_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_13_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_13_pad_iopad (
            .OE(N__81268),
            .DIN(N__81267),
            .DOUT(N__81266),
            .PACKAGEPIN(PIN_13));
    defparam PIN_13_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_13_pad_preio (
            .PADOEN(N__81268),
            .PADOUT(N__81267),
            .PADIN(N__81266),
            .CLOCKENABLE(),
            .DIN0(PIN_13_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_1_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_1_pad_iopad (
            .OE(N__81259),
            .DIN(N__81258),
            .DOUT(N__81257),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_1_pad_preio (
            .PADOEN(N__81259),
            .PADOUT(N__81258),
            .PADIN(N__81257),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_22_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_22_pad_iopad (
            .OE(N__81250),
            .DIN(N__81249),
            .DOUT(N__81248),
            .PACKAGEPIN(PIN_22));
    defparam PIN_22_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_22_pad_preio (
            .PADOEN(N__81250),
            .PADOUT(N__81249),
            .PADIN(N__81248),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_23_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_23_pad_iopad (
            .OE(N__81241),
            .DIN(N__81240),
            .DOUT(N__81239),
            .PACKAGEPIN(PIN_23));
    defparam PIN_23_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_23_pad_preio (
            .PADOEN(N__81241),
            .PADOUT(N__81240),
            .PADIN(N__81239),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_24_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_24_pad_iopad (
            .OE(N__81232),
            .DIN(N__81231),
            .DOUT(N__81230),
            .PACKAGEPIN(PIN_24));
    defparam PIN_24_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_24_pad_preio (
            .PADOEN(N__81232),
            .PADOUT(N__81231),
            .PADIN(N__81230),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__81223),
            .DIN(N__81222),
            .DOUT(N__81221),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__81223),
            .PADOUT(N__81222),
            .PADIN(N__81221),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_3_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_3_pad_iopad (
            .OE(N__81214),
            .DIN(N__81213),
            .DOUT(N__81212),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_3_pad_preio (
            .PADOEN(N__81214),
            .PADOUT(N__81213),
            .PADIN(N__81212),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_7_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_7_pad_iopad (
            .OE(N__81205),
            .DIN(N__81204),
            .DOUT(N__81203),
            .PACKAGEPIN(PIN_7));
    defparam PIN_7_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_7_pad_preio (
            .PADOEN(N__81205),
            .PADOUT(N__81204),
            .PADIN(N__81203),
            .CLOCKENABLE(),
            .DIN0(PIN_7_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_8_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_8_pad_iopad (
            .OE(N__81196),
            .DIN(N__81195),
            .DOUT(N__81194),
            .PACKAGEPIN(PIN_8));
    defparam PIN_8_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_8_pad_preio (
            .PADOEN(N__81196),
            .PADOUT(N__81195),
            .PADIN(N__81194),
            .CLOCKENABLE(),
            .DIN0(PIN_8_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__81187),
            .DIN(N__81186),
            .DOUT(N__81185),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__81187),
            .PADOUT(N__81186),
            .PADIN(N__81185),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__81178),
            .DIN(N__81177),
            .DOUT(N__81176),
            .PACKAGEPIN(PIN_4));
    defparam hall1_input_preio.PIN_TYPE=6'b000001;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__81178),
            .PADOUT(N__81177),
            .PADIN(N__81176),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__81169),
            .DIN(N__81168),
            .DOUT(N__81167),
            .PACKAGEPIN(PIN_5));
    defparam hall2_input_preio.PIN_TYPE=6'b000001;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__81169),
            .PADOUT(N__81168),
            .PADIN(N__81167),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__81160),
            .DIN(N__81159),
            .DOUT(N__81158),
            .PACKAGEPIN(PIN_6));
    defparam hall3_input_preio.PIN_TYPE=6'b000001;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__81160),
            .PADOUT(N__81159),
            .PADIN(N__81158),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__81151),
            .DIN(N__81150),
            .DOUT(N__81149),
            .PACKAGEPIN(PIN_11));
    defparam rx_input_preio.PIN_TYPE=6'b000001;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__81151),
            .PADOUT(N__81150),
            .PADIN(N__81149),
            .CLOCKENABLE(),
            .DIN0(LED_c),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__81142),
            .DIN(N__81141),
            .DOUT(N__81140),
            .PACKAGEPIN(PIN_10));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__81142),
            .PADOUT(N__81141),
            .PADIN(N__81140),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__28599),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__26757));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__81133),
            .DIN(N__81132),
            .DOUT(N__81131),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__81133),
            .PADOUT(N__81132),
            .PADIN(N__81131),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__20379 (
            .O(N__81114),
            .I(N__81111));
    InMux I__20378 (
            .O(N__81111),
            .I(N__81108));
    LocalMux I__20377 (
            .O(N__81108),
            .I(N__81105));
    Span4Mux_h I__20376 (
            .O(N__81105),
            .I(N__81100));
    InMux I__20375 (
            .O(N__81104),
            .I(N__81097));
    InMux I__20374 (
            .O(N__81103),
            .I(N__81094));
    Span4Mux_v I__20373 (
            .O(N__81100),
            .I(N__81091));
    LocalMux I__20372 (
            .O(N__81097),
            .I(N__81086));
    LocalMux I__20371 (
            .O(N__81094),
            .I(N__81086));
    Odrv4 I__20370 (
            .O(N__81091),
            .I(\c0.n19_adj_4595 ));
    Odrv12 I__20369 (
            .O(N__81086),
            .I(\c0.n19_adj_4595 ));
    InMux I__20368 (
            .O(N__81081),
            .I(N__81078));
    LocalMux I__20367 (
            .O(N__81078),
            .I(\c0.n24_adj_4628 ));
    CascadeMux I__20366 (
            .O(N__81075),
            .I(\c0.n14_adj_4629_cascade_ ));
    InMux I__20365 (
            .O(N__81072),
            .I(N__81068));
    InMux I__20364 (
            .O(N__81071),
            .I(N__81065));
    LocalMux I__20363 (
            .O(N__81068),
            .I(N__81062));
    LocalMux I__20362 (
            .O(N__81065),
            .I(N__81059));
    Span4Mux_v I__20361 (
            .O(N__81062),
            .I(N__81054));
    Span4Mux_h I__20360 (
            .O(N__81059),
            .I(N__81051));
    InMux I__20359 (
            .O(N__81058),
            .I(N__81048));
    InMux I__20358 (
            .O(N__81057),
            .I(N__81045));
    Span4Mux_h I__20357 (
            .O(N__81054),
            .I(N__81042));
    Span4Mux_h I__20356 (
            .O(N__81051),
            .I(N__81039));
    LocalMux I__20355 (
            .O(N__81048),
            .I(N__81036));
    LocalMux I__20354 (
            .O(N__81045),
            .I(N__81033));
    Span4Mux_v I__20353 (
            .O(N__81042),
            .I(N__81028));
    Span4Mux_v I__20352 (
            .O(N__81039),
            .I(N__81025));
    Span4Mux_v I__20351 (
            .O(N__81036),
            .I(N__81020));
    Span4Mux_h I__20350 (
            .O(N__81033),
            .I(N__81020));
    InMux I__20349 (
            .O(N__81032),
            .I(N__81015));
    InMux I__20348 (
            .O(N__81031),
            .I(N__81015));
    Odrv4 I__20347 (
            .O(N__81028),
            .I(\c0.n23178 ));
    Odrv4 I__20346 (
            .O(N__81025),
            .I(\c0.n23178 ));
    Odrv4 I__20345 (
            .O(N__81020),
            .I(\c0.n23178 ));
    LocalMux I__20344 (
            .O(N__81015),
            .I(\c0.n23178 ));
    InMux I__20343 (
            .O(N__81006),
            .I(N__81003));
    LocalMux I__20342 (
            .O(N__81003),
            .I(N__80999));
    InMux I__20341 (
            .O(N__81002),
            .I(N__80996));
    Span4Mux_v I__20340 (
            .O(N__80999),
            .I(N__80991));
    LocalMux I__20339 (
            .O(N__80996),
            .I(N__80991));
    Odrv4 I__20338 (
            .O(N__80991),
            .I(\c0.n22234 ));
    InMux I__20337 (
            .O(N__80988),
            .I(N__80983));
    InMux I__20336 (
            .O(N__80987),
            .I(N__80979));
    CascadeMux I__20335 (
            .O(N__80986),
            .I(N__80976));
    LocalMux I__20334 (
            .O(N__80983),
            .I(N__80970));
    CascadeMux I__20333 (
            .O(N__80982),
            .I(N__80967));
    LocalMux I__20332 (
            .O(N__80979),
            .I(N__80963));
    InMux I__20331 (
            .O(N__80976),
            .I(N__80960));
    InMux I__20330 (
            .O(N__80975),
            .I(N__80957));
    InMux I__20329 (
            .O(N__80974),
            .I(N__80952));
    InMux I__20328 (
            .O(N__80973),
            .I(N__80952));
    Span4Mux_v I__20327 (
            .O(N__80970),
            .I(N__80948));
    InMux I__20326 (
            .O(N__80967),
            .I(N__80945));
    InMux I__20325 (
            .O(N__80966),
            .I(N__80937));
    Span4Mux_v I__20324 (
            .O(N__80963),
            .I(N__80928));
    LocalMux I__20323 (
            .O(N__80960),
            .I(N__80928));
    LocalMux I__20322 (
            .O(N__80957),
            .I(N__80928));
    LocalMux I__20321 (
            .O(N__80952),
            .I(N__80928));
    CascadeMux I__20320 (
            .O(N__80951),
            .I(N__80925));
    Span4Mux_h I__20319 (
            .O(N__80948),
            .I(N__80913));
    LocalMux I__20318 (
            .O(N__80945),
            .I(N__80913));
    InMux I__20317 (
            .O(N__80944),
            .I(N__80908));
    InMux I__20316 (
            .O(N__80943),
            .I(N__80908));
    InMux I__20315 (
            .O(N__80942),
            .I(N__80905));
    InMux I__20314 (
            .O(N__80941),
            .I(N__80900));
    InMux I__20313 (
            .O(N__80940),
            .I(N__80900));
    LocalMux I__20312 (
            .O(N__80937),
            .I(N__80894));
    Span4Mux_v I__20311 (
            .O(N__80928),
            .I(N__80894));
    InMux I__20310 (
            .O(N__80925),
            .I(N__80889));
    InMux I__20309 (
            .O(N__80924),
            .I(N__80889));
    InMux I__20308 (
            .O(N__80923),
            .I(N__80885));
    InMux I__20307 (
            .O(N__80922),
            .I(N__80882));
    InMux I__20306 (
            .O(N__80921),
            .I(N__80875));
    InMux I__20305 (
            .O(N__80920),
            .I(N__80875));
    InMux I__20304 (
            .O(N__80919),
            .I(N__80875));
    InMux I__20303 (
            .O(N__80918),
            .I(N__80872));
    Span4Mux_v I__20302 (
            .O(N__80913),
            .I(N__80868));
    LocalMux I__20301 (
            .O(N__80908),
            .I(N__80864));
    LocalMux I__20300 (
            .O(N__80905),
            .I(N__80859));
    LocalMux I__20299 (
            .O(N__80900),
            .I(N__80859));
    InMux I__20298 (
            .O(N__80899),
            .I(N__80856));
    Span4Mux_h I__20297 (
            .O(N__80894),
            .I(N__80853));
    LocalMux I__20296 (
            .O(N__80889),
            .I(N__80850));
    InMux I__20295 (
            .O(N__80888),
            .I(N__80847));
    LocalMux I__20294 (
            .O(N__80885),
            .I(N__80844));
    LocalMux I__20293 (
            .O(N__80882),
            .I(N__80840));
    LocalMux I__20292 (
            .O(N__80875),
            .I(N__80837));
    LocalMux I__20291 (
            .O(N__80872),
            .I(N__80834));
    InMux I__20290 (
            .O(N__80871),
            .I(N__80831));
    Span4Mux_v I__20289 (
            .O(N__80868),
            .I(N__80828));
    InMux I__20288 (
            .O(N__80867),
            .I(N__80825));
    Span4Mux_h I__20287 (
            .O(N__80864),
            .I(N__80820));
    Span4Mux_v I__20286 (
            .O(N__80859),
            .I(N__80820));
    LocalMux I__20285 (
            .O(N__80856),
            .I(N__80813));
    Span4Mux_h I__20284 (
            .O(N__80853),
            .I(N__80813));
    Span4Mux_v I__20283 (
            .O(N__80850),
            .I(N__80813));
    LocalMux I__20282 (
            .O(N__80847),
            .I(N__80810));
    Span4Mux_v I__20281 (
            .O(N__80844),
            .I(N__80807));
    InMux I__20280 (
            .O(N__80843),
            .I(N__80804));
    Span4Mux_h I__20279 (
            .O(N__80840),
            .I(N__80799));
    Span4Mux_v I__20278 (
            .O(N__80837),
            .I(N__80799));
    Sp12to4 I__20277 (
            .O(N__80834),
            .I(N__80796));
    LocalMux I__20276 (
            .O(N__80831),
            .I(N__80793));
    Span4Mux_h I__20275 (
            .O(N__80828),
            .I(N__80790));
    LocalMux I__20274 (
            .O(N__80825),
            .I(N__80787));
    Span4Mux_h I__20273 (
            .O(N__80820),
            .I(N__80784));
    Span4Mux_v I__20272 (
            .O(N__80813),
            .I(N__80781));
    Span4Mux_v I__20271 (
            .O(N__80810),
            .I(N__80776));
    Span4Mux_h I__20270 (
            .O(N__80807),
            .I(N__80776));
    LocalMux I__20269 (
            .O(N__80804),
            .I(N__80769));
    Sp12to4 I__20268 (
            .O(N__80799),
            .I(N__80769));
    Span12Mux_v I__20267 (
            .O(N__80796),
            .I(N__80769));
    Span4Mux_h I__20266 (
            .O(N__80793),
            .I(N__80764));
    Span4Mux_h I__20265 (
            .O(N__80790),
            .I(N__80764));
    Span4Mux_v I__20264 (
            .O(N__80787),
            .I(N__80757));
    Span4Mux_h I__20263 (
            .O(N__80784),
            .I(N__80757));
    Span4Mux_v I__20262 (
            .O(N__80781),
            .I(N__80757));
    Odrv4 I__20261 (
            .O(N__80776),
            .I(\c0.n17830 ));
    Odrv12 I__20260 (
            .O(N__80769),
            .I(\c0.n17830 ));
    Odrv4 I__20259 (
            .O(N__80764),
            .I(\c0.n17830 ));
    Odrv4 I__20258 (
            .O(N__80757),
            .I(\c0.n17830 ));
    InMux I__20257 (
            .O(N__80748),
            .I(N__80743));
    CascadeMux I__20256 (
            .O(N__80747),
            .I(N__80730));
    InMux I__20255 (
            .O(N__80746),
            .I(N__80726));
    LocalMux I__20254 (
            .O(N__80743),
            .I(N__80723));
    InMux I__20253 (
            .O(N__80742),
            .I(N__80720));
    InMux I__20252 (
            .O(N__80741),
            .I(N__80715));
    InMux I__20251 (
            .O(N__80740),
            .I(N__80712));
    CascadeMux I__20250 (
            .O(N__80739),
            .I(N__80708));
    InMux I__20249 (
            .O(N__80738),
            .I(N__80704));
    InMux I__20248 (
            .O(N__80737),
            .I(N__80700));
    CascadeMux I__20247 (
            .O(N__80736),
            .I(N__80697));
    CascadeMux I__20246 (
            .O(N__80735),
            .I(N__80693));
    InMux I__20245 (
            .O(N__80734),
            .I(N__80688));
    InMux I__20244 (
            .O(N__80733),
            .I(N__80688));
    InMux I__20243 (
            .O(N__80730),
            .I(N__80685));
    InMux I__20242 (
            .O(N__80729),
            .I(N__80682));
    LocalMux I__20241 (
            .O(N__80726),
            .I(N__80679));
    Span4Mux_h I__20240 (
            .O(N__80723),
            .I(N__80674));
    LocalMux I__20239 (
            .O(N__80720),
            .I(N__80674));
    InMux I__20238 (
            .O(N__80719),
            .I(N__80668));
    InMux I__20237 (
            .O(N__80718),
            .I(N__80665));
    LocalMux I__20236 (
            .O(N__80715),
            .I(N__80662));
    LocalMux I__20235 (
            .O(N__80712),
            .I(N__80659));
    InMux I__20234 (
            .O(N__80711),
            .I(N__80656));
    InMux I__20233 (
            .O(N__80708),
            .I(N__80650));
    InMux I__20232 (
            .O(N__80707),
            .I(N__80650));
    LocalMux I__20231 (
            .O(N__80704),
            .I(N__80647));
    InMux I__20230 (
            .O(N__80703),
            .I(N__80644));
    LocalMux I__20229 (
            .O(N__80700),
            .I(N__80641));
    InMux I__20228 (
            .O(N__80697),
            .I(N__80638));
    InMux I__20227 (
            .O(N__80696),
            .I(N__80635));
    InMux I__20226 (
            .O(N__80693),
            .I(N__80632));
    LocalMux I__20225 (
            .O(N__80688),
            .I(N__80627));
    LocalMux I__20224 (
            .O(N__80685),
            .I(N__80627));
    LocalMux I__20223 (
            .O(N__80682),
            .I(N__80624));
    Span4Mux_v I__20222 (
            .O(N__80679),
            .I(N__80619));
    Span4Mux_v I__20221 (
            .O(N__80674),
            .I(N__80619));
    CascadeMux I__20220 (
            .O(N__80673),
            .I(N__80612));
    InMux I__20219 (
            .O(N__80672),
            .I(N__80609));
    CascadeMux I__20218 (
            .O(N__80671),
            .I(N__80606));
    LocalMux I__20217 (
            .O(N__80668),
            .I(N__80602));
    LocalMux I__20216 (
            .O(N__80665),
            .I(N__80595));
    Span4Mux_h I__20215 (
            .O(N__80662),
            .I(N__80595));
    Span4Mux_v I__20214 (
            .O(N__80659),
            .I(N__80595));
    LocalMux I__20213 (
            .O(N__80656),
            .I(N__80592));
    InMux I__20212 (
            .O(N__80655),
            .I(N__80589));
    LocalMux I__20211 (
            .O(N__80650),
            .I(N__80586));
    Span4Mux_h I__20210 (
            .O(N__80647),
            .I(N__80581));
    LocalMux I__20209 (
            .O(N__80644),
            .I(N__80581));
    Span4Mux_v I__20208 (
            .O(N__80641),
            .I(N__80576));
    LocalMux I__20207 (
            .O(N__80638),
            .I(N__80576));
    LocalMux I__20206 (
            .O(N__80635),
            .I(N__80568));
    LocalMux I__20205 (
            .O(N__80632),
            .I(N__80568));
    Span4Mux_v I__20204 (
            .O(N__80627),
            .I(N__80568));
    Span4Mux_v I__20203 (
            .O(N__80624),
            .I(N__80565));
    Span4Mux_h I__20202 (
            .O(N__80619),
            .I(N__80562));
    InMux I__20201 (
            .O(N__80618),
            .I(N__80557));
    InMux I__20200 (
            .O(N__80617),
            .I(N__80557));
    InMux I__20199 (
            .O(N__80616),
            .I(N__80554));
    InMux I__20198 (
            .O(N__80615),
            .I(N__80549));
    InMux I__20197 (
            .O(N__80612),
            .I(N__80549));
    LocalMux I__20196 (
            .O(N__80609),
            .I(N__80546));
    InMux I__20195 (
            .O(N__80606),
            .I(N__80543));
    InMux I__20194 (
            .O(N__80605),
            .I(N__80540));
    Span4Mux_v I__20193 (
            .O(N__80602),
            .I(N__80535));
    Span4Mux_v I__20192 (
            .O(N__80595),
            .I(N__80535));
    Span4Mux_v I__20191 (
            .O(N__80592),
            .I(N__80532));
    LocalMux I__20190 (
            .O(N__80589),
            .I(N__80527));
    Span4Mux_v I__20189 (
            .O(N__80586),
            .I(N__80527));
    Span4Mux_v I__20188 (
            .O(N__80581),
            .I(N__80524));
    Span4Mux_h I__20187 (
            .O(N__80576),
            .I(N__80521));
    InMux I__20186 (
            .O(N__80575),
            .I(N__80518));
    Span4Mux_v I__20185 (
            .O(N__80568),
            .I(N__80515));
    Span4Mux_v I__20184 (
            .O(N__80565),
            .I(N__80510));
    Span4Mux_h I__20183 (
            .O(N__80562),
            .I(N__80510));
    LocalMux I__20182 (
            .O(N__80557),
            .I(N__80505));
    LocalMux I__20181 (
            .O(N__80554),
            .I(N__80502));
    LocalMux I__20180 (
            .O(N__80549),
            .I(N__80497));
    Span4Mux_v I__20179 (
            .O(N__80546),
            .I(N__80497));
    LocalMux I__20178 (
            .O(N__80543),
            .I(N__80492));
    LocalMux I__20177 (
            .O(N__80540),
            .I(N__80492));
    Span4Mux_h I__20176 (
            .O(N__80535),
            .I(N__80487));
    Span4Mux_v I__20175 (
            .O(N__80532),
            .I(N__80487));
    Span4Mux_v I__20174 (
            .O(N__80527),
            .I(N__80484));
    Sp12to4 I__20173 (
            .O(N__80524),
            .I(N__80481));
    Sp12to4 I__20172 (
            .O(N__80521),
            .I(N__80478));
    LocalMux I__20171 (
            .O(N__80518),
            .I(N__80471));
    Sp12to4 I__20170 (
            .O(N__80515),
            .I(N__80471));
    Sp12to4 I__20169 (
            .O(N__80510),
            .I(N__80471));
    InMux I__20168 (
            .O(N__80509),
            .I(N__80466));
    InMux I__20167 (
            .O(N__80508),
            .I(N__80466));
    Span12Mux_h I__20166 (
            .O(N__80505),
            .I(N__80463));
    Span4Mux_h I__20165 (
            .O(N__80502),
            .I(N__80458));
    Span4Mux_h I__20164 (
            .O(N__80497),
            .I(N__80458));
    Span4Mux_v I__20163 (
            .O(N__80492),
            .I(N__80453));
    Span4Mux_v I__20162 (
            .O(N__80487),
            .I(N__80453));
    Sp12to4 I__20161 (
            .O(N__80484),
            .I(N__80444));
    Span12Mux_h I__20160 (
            .O(N__80481),
            .I(N__80444));
    Span12Mux_v I__20159 (
            .O(N__80478),
            .I(N__80444));
    Span12Mux_h I__20158 (
            .O(N__80471),
            .I(N__80444));
    LocalMux I__20157 (
            .O(N__80466),
            .I(rx_data_0));
    Odrv12 I__20156 (
            .O(N__80463),
            .I(rx_data_0));
    Odrv4 I__20155 (
            .O(N__80458),
            .I(rx_data_0));
    Odrv4 I__20154 (
            .O(N__80453),
            .I(rx_data_0));
    Odrv12 I__20153 (
            .O(N__80444),
            .I(rx_data_0));
    InMux I__20152 (
            .O(N__80433),
            .I(N__80407));
    InMux I__20151 (
            .O(N__80432),
            .I(N__80407));
    InMux I__20150 (
            .O(N__80431),
            .I(N__80404));
    InMux I__20149 (
            .O(N__80430),
            .I(N__80392));
    InMux I__20148 (
            .O(N__80429),
            .I(N__80389));
    InMux I__20147 (
            .O(N__80428),
            .I(N__80386));
    InMux I__20146 (
            .O(N__80427),
            .I(N__80382));
    InMux I__20145 (
            .O(N__80426),
            .I(N__80379));
    InMux I__20144 (
            .O(N__80425),
            .I(N__80376));
    InMux I__20143 (
            .O(N__80424),
            .I(N__80373));
    InMux I__20142 (
            .O(N__80423),
            .I(N__80368));
    InMux I__20141 (
            .O(N__80422),
            .I(N__80368));
    InMux I__20140 (
            .O(N__80421),
            .I(N__80365));
    InMux I__20139 (
            .O(N__80420),
            .I(N__80360));
    InMux I__20138 (
            .O(N__80419),
            .I(N__80360));
    InMux I__20137 (
            .O(N__80418),
            .I(N__80355));
    InMux I__20136 (
            .O(N__80417),
            .I(N__80355));
    InMux I__20135 (
            .O(N__80416),
            .I(N__80344));
    InMux I__20134 (
            .O(N__80415),
            .I(N__80344));
    InMux I__20133 (
            .O(N__80414),
            .I(N__80344));
    InMux I__20132 (
            .O(N__80413),
            .I(N__80344));
    InMux I__20131 (
            .O(N__80412),
            .I(N__80344));
    LocalMux I__20130 (
            .O(N__80407),
            .I(N__80341));
    LocalMux I__20129 (
            .O(N__80404),
            .I(N__80338));
    InMux I__20128 (
            .O(N__80403),
            .I(N__80329));
    InMux I__20127 (
            .O(N__80402),
            .I(N__80329));
    InMux I__20126 (
            .O(N__80401),
            .I(N__80329));
    InMux I__20125 (
            .O(N__80400),
            .I(N__80329));
    InMux I__20124 (
            .O(N__80399),
            .I(N__80325));
    InMux I__20123 (
            .O(N__80398),
            .I(N__80315));
    InMux I__20122 (
            .O(N__80397),
            .I(N__80312));
    InMux I__20121 (
            .O(N__80396),
            .I(N__80307));
    InMux I__20120 (
            .O(N__80395),
            .I(N__80307));
    LocalMux I__20119 (
            .O(N__80392),
            .I(N__80304));
    LocalMux I__20118 (
            .O(N__80389),
            .I(N__80299));
    LocalMux I__20117 (
            .O(N__80386),
            .I(N__80299));
    InMux I__20116 (
            .O(N__80385),
            .I(N__80296));
    LocalMux I__20115 (
            .O(N__80382),
            .I(N__80293));
    LocalMux I__20114 (
            .O(N__80379),
            .I(N__80288));
    LocalMux I__20113 (
            .O(N__80376),
            .I(N__80288));
    LocalMux I__20112 (
            .O(N__80373),
            .I(N__80283));
    LocalMux I__20111 (
            .O(N__80368),
            .I(N__80283));
    LocalMux I__20110 (
            .O(N__80365),
            .I(N__80276));
    LocalMux I__20109 (
            .O(N__80360),
            .I(N__80276));
    LocalMux I__20108 (
            .O(N__80355),
            .I(N__80276));
    LocalMux I__20107 (
            .O(N__80344),
            .I(N__80267));
    Span4Mux_v I__20106 (
            .O(N__80341),
            .I(N__80267));
    Span4Mux_v I__20105 (
            .O(N__80338),
            .I(N__80267));
    LocalMux I__20104 (
            .O(N__80329),
            .I(N__80267));
    InMux I__20103 (
            .O(N__80328),
            .I(N__80256));
    LocalMux I__20102 (
            .O(N__80325),
            .I(N__80253));
    InMux I__20101 (
            .O(N__80324),
            .I(N__80250));
    InMux I__20100 (
            .O(N__80323),
            .I(N__80241));
    InMux I__20099 (
            .O(N__80322),
            .I(N__80241));
    InMux I__20098 (
            .O(N__80321),
            .I(N__80241));
    InMux I__20097 (
            .O(N__80320),
            .I(N__80241));
    InMux I__20096 (
            .O(N__80319),
            .I(N__80236));
    InMux I__20095 (
            .O(N__80318),
            .I(N__80236));
    LocalMux I__20094 (
            .O(N__80315),
            .I(N__80233));
    LocalMux I__20093 (
            .O(N__80312),
            .I(N__80230));
    LocalMux I__20092 (
            .O(N__80307),
            .I(N__80227));
    Span4Mux_v I__20091 (
            .O(N__80304),
            .I(N__80224));
    Span4Mux_v I__20090 (
            .O(N__80299),
            .I(N__80221));
    LocalMux I__20089 (
            .O(N__80296),
            .I(N__80218));
    Span4Mux_h I__20088 (
            .O(N__80293),
            .I(N__80213));
    Span4Mux_v I__20087 (
            .O(N__80288),
            .I(N__80213));
    Span4Mux_v I__20086 (
            .O(N__80283),
            .I(N__80206));
    Span4Mux_v I__20085 (
            .O(N__80276),
            .I(N__80206));
    Span4Mux_h I__20084 (
            .O(N__80267),
            .I(N__80206));
    InMux I__20083 (
            .O(N__80266),
            .I(N__80203));
    InMux I__20082 (
            .O(N__80265),
            .I(N__80200));
    InMux I__20081 (
            .O(N__80264),
            .I(N__80197));
    InMux I__20080 (
            .O(N__80263),
            .I(N__80186));
    InMux I__20079 (
            .O(N__80262),
            .I(N__80186));
    InMux I__20078 (
            .O(N__80261),
            .I(N__80186));
    InMux I__20077 (
            .O(N__80260),
            .I(N__80186));
    InMux I__20076 (
            .O(N__80259),
            .I(N__80186));
    LocalMux I__20075 (
            .O(N__80256),
            .I(N__80183));
    Span4Mux_h I__20074 (
            .O(N__80253),
            .I(N__80180));
    LocalMux I__20073 (
            .O(N__80250),
            .I(N__80171));
    LocalMux I__20072 (
            .O(N__80241),
            .I(N__80171));
    LocalMux I__20071 (
            .O(N__80236),
            .I(N__80171));
    Span12Mux_v I__20070 (
            .O(N__80233),
            .I(N__80171));
    Span4Mux_v I__20069 (
            .O(N__80230),
            .I(N__80162));
    Span4Mux_v I__20068 (
            .O(N__80227),
            .I(N__80162));
    Span4Mux_h I__20067 (
            .O(N__80224),
            .I(N__80162));
    Span4Mux_h I__20066 (
            .O(N__80221),
            .I(N__80162));
    Span4Mux_h I__20065 (
            .O(N__80218),
            .I(N__80155));
    Span4Mux_v I__20064 (
            .O(N__80213),
            .I(N__80155));
    Span4Mux_h I__20063 (
            .O(N__80206),
            .I(N__80155));
    LocalMux I__20062 (
            .O(N__80203),
            .I(\c0.n22104 ));
    LocalMux I__20061 (
            .O(N__80200),
            .I(\c0.n22104 ));
    LocalMux I__20060 (
            .O(N__80197),
            .I(\c0.n22104 ));
    LocalMux I__20059 (
            .O(N__80186),
            .I(\c0.n22104 ));
    Odrv4 I__20058 (
            .O(N__80183),
            .I(\c0.n22104 ));
    Odrv4 I__20057 (
            .O(N__80180),
            .I(\c0.n22104 ));
    Odrv12 I__20056 (
            .O(N__80171),
            .I(\c0.n22104 ));
    Odrv4 I__20055 (
            .O(N__80162),
            .I(\c0.n22104 ));
    Odrv4 I__20054 (
            .O(N__80155),
            .I(\c0.n22104 ));
    InMux I__20053 (
            .O(N__80136),
            .I(N__80132));
    InMux I__20052 (
            .O(N__80135),
            .I(N__80128));
    LocalMux I__20051 (
            .O(N__80132),
            .I(N__80125));
    CascadeMux I__20050 (
            .O(N__80131),
            .I(N__80122));
    LocalMux I__20049 (
            .O(N__80128),
            .I(N__80119));
    Span4Mux_h I__20048 (
            .O(N__80125),
            .I(N__80116));
    InMux I__20047 (
            .O(N__80122),
            .I(N__80113));
    Span4Mux_h I__20046 (
            .O(N__80119),
            .I(N__80110));
    Span4Mux_h I__20045 (
            .O(N__80116),
            .I(N__80107));
    LocalMux I__20044 (
            .O(N__80113),
            .I(\c0.data_in_frame_23_0 ));
    Odrv4 I__20043 (
            .O(N__80110),
            .I(\c0.data_in_frame_23_0 ));
    Odrv4 I__20042 (
            .O(N__80107),
            .I(\c0.data_in_frame_23_0 ));
    CascadeMux I__20041 (
            .O(N__80100),
            .I(N__80090));
    CascadeMux I__20040 (
            .O(N__80099),
            .I(N__80087));
    CascadeMux I__20039 (
            .O(N__80098),
            .I(N__80084));
    CascadeMux I__20038 (
            .O(N__80097),
            .I(N__80081));
    InMux I__20037 (
            .O(N__80096),
            .I(N__80076));
    InMux I__20036 (
            .O(N__80095),
            .I(N__80073));
    InMux I__20035 (
            .O(N__80094),
            .I(N__80070));
    InMux I__20034 (
            .O(N__80093),
            .I(N__80067));
    InMux I__20033 (
            .O(N__80090),
            .I(N__80064));
    InMux I__20032 (
            .O(N__80087),
            .I(N__80061));
    InMux I__20031 (
            .O(N__80084),
            .I(N__80055));
    InMux I__20030 (
            .O(N__80081),
            .I(N__80055));
    CascadeMux I__20029 (
            .O(N__80080),
            .I(N__80052));
    InMux I__20028 (
            .O(N__80079),
            .I(N__80048));
    LocalMux I__20027 (
            .O(N__80076),
            .I(N__80045));
    LocalMux I__20026 (
            .O(N__80073),
            .I(N__80041));
    LocalMux I__20025 (
            .O(N__80070),
            .I(N__80036));
    LocalMux I__20024 (
            .O(N__80067),
            .I(N__80036));
    LocalMux I__20023 (
            .O(N__80064),
            .I(N__80033));
    LocalMux I__20022 (
            .O(N__80061),
            .I(N__80026));
    InMux I__20021 (
            .O(N__80060),
            .I(N__80023));
    LocalMux I__20020 (
            .O(N__80055),
            .I(N__80020));
    InMux I__20019 (
            .O(N__80052),
            .I(N__80017));
    InMux I__20018 (
            .O(N__80051),
            .I(N__80013));
    LocalMux I__20017 (
            .O(N__80048),
            .I(N__80010));
    Span4Mux_h I__20016 (
            .O(N__80045),
            .I(N__80004));
    InMux I__20015 (
            .O(N__80044),
            .I(N__80001));
    Span4Mux_h I__20014 (
            .O(N__80041),
            .I(N__79998));
    Span4Mux_v I__20013 (
            .O(N__80036),
            .I(N__79995));
    Span4Mux_h I__20012 (
            .O(N__80033),
            .I(N__79992));
    CascadeMux I__20011 (
            .O(N__80032),
            .I(N__79989));
    InMux I__20010 (
            .O(N__80031),
            .I(N__79980));
    InMux I__20009 (
            .O(N__80030),
            .I(N__79975));
    InMux I__20008 (
            .O(N__80029),
            .I(N__79975));
    Span4Mux_h I__20007 (
            .O(N__80026),
            .I(N__79972));
    LocalMux I__20006 (
            .O(N__80023),
            .I(N__79967));
    Span4Mux_v I__20005 (
            .O(N__80020),
            .I(N__79967));
    LocalMux I__20004 (
            .O(N__80017),
            .I(N__79964));
    InMux I__20003 (
            .O(N__80016),
            .I(N__79961));
    LocalMux I__20002 (
            .O(N__80013),
            .I(N__79958));
    Span4Mux_h I__20001 (
            .O(N__80010),
            .I(N__79955));
    CascadeMux I__20000 (
            .O(N__80009),
            .I(N__79949));
    InMux I__19999 (
            .O(N__80008),
            .I(N__79944));
    InMux I__19998 (
            .O(N__80007),
            .I(N__79941));
    Span4Mux_h I__19997 (
            .O(N__80004),
            .I(N__79938));
    LocalMux I__19996 (
            .O(N__80001),
            .I(N__79929));
    Span4Mux_h I__19995 (
            .O(N__79998),
            .I(N__79929));
    Span4Mux_h I__19994 (
            .O(N__79995),
            .I(N__79929));
    Span4Mux_v I__19993 (
            .O(N__79992),
            .I(N__79929));
    InMux I__19992 (
            .O(N__79989),
            .I(N__79922));
    InMux I__19991 (
            .O(N__79988),
            .I(N__79922));
    InMux I__19990 (
            .O(N__79987),
            .I(N__79922));
    InMux I__19989 (
            .O(N__79986),
            .I(N__79919));
    InMux I__19988 (
            .O(N__79985),
            .I(N__79914));
    InMux I__19987 (
            .O(N__79984),
            .I(N__79914));
    InMux I__19986 (
            .O(N__79983),
            .I(N__79911));
    LocalMux I__19985 (
            .O(N__79980),
            .I(N__79908));
    LocalMux I__19984 (
            .O(N__79975),
            .I(N__79901));
    Span4Mux_h I__19983 (
            .O(N__79972),
            .I(N__79901));
    Span4Mux_h I__19982 (
            .O(N__79967),
            .I(N__79901));
    Span4Mux_v I__19981 (
            .O(N__79964),
            .I(N__79892));
    LocalMux I__19980 (
            .O(N__79961),
            .I(N__79892));
    Span4Mux_h I__19979 (
            .O(N__79958),
            .I(N__79892));
    Span4Mux_v I__19978 (
            .O(N__79955),
            .I(N__79892));
    CascadeMux I__19977 (
            .O(N__79954),
            .I(N__79889));
    InMux I__19976 (
            .O(N__79953),
            .I(N__79886));
    InMux I__19975 (
            .O(N__79952),
            .I(N__79883));
    InMux I__19974 (
            .O(N__79949),
            .I(N__79878));
    InMux I__19973 (
            .O(N__79948),
            .I(N__79878));
    InMux I__19972 (
            .O(N__79947),
            .I(N__79875));
    LocalMux I__19971 (
            .O(N__79944),
            .I(N__79868));
    LocalMux I__19970 (
            .O(N__79941),
            .I(N__79868));
    Span4Mux_h I__19969 (
            .O(N__79938),
            .I(N__79868));
    Span4Mux_v I__19968 (
            .O(N__79929),
            .I(N__79865));
    LocalMux I__19967 (
            .O(N__79922),
            .I(N__79860));
    LocalMux I__19966 (
            .O(N__79919),
            .I(N__79860));
    LocalMux I__19965 (
            .O(N__79914),
            .I(N__79857));
    LocalMux I__19964 (
            .O(N__79911),
            .I(N__79848));
    Span12Mux_s10_v I__19963 (
            .O(N__79908),
            .I(N__79848));
    Sp12to4 I__19962 (
            .O(N__79901),
            .I(N__79848));
    Sp12to4 I__19961 (
            .O(N__79892),
            .I(N__79848));
    InMux I__19960 (
            .O(N__79889),
            .I(N__79845));
    LocalMux I__19959 (
            .O(N__79886),
            .I(N__79842));
    LocalMux I__19958 (
            .O(N__79883),
            .I(N__79833));
    LocalMux I__19957 (
            .O(N__79878),
            .I(N__79833));
    LocalMux I__19956 (
            .O(N__79875),
            .I(N__79833));
    Span4Mux_v I__19955 (
            .O(N__79868),
            .I(N__79833));
    Span4Mux_v I__19954 (
            .O(N__79865),
            .I(N__79830));
    Span4Mux_v I__19953 (
            .O(N__79860),
            .I(N__79827));
    Span12Mux_v I__19952 (
            .O(N__79857),
            .I(N__79824));
    Span12Mux_v I__19951 (
            .O(N__79848),
            .I(N__79821));
    LocalMux I__19950 (
            .O(N__79845),
            .I(N__79814));
    Span4Mux_h I__19949 (
            .O(N__79842),
            .I(N__79814));
    Span4Mux_v I__19948 (
            .O(N__79833),
            .I(N__79814));
    Span4Mux_v I__19947 (
            .O(N__79830),
            .I(N__79811));
    Odrv4 I__19946 (
            .O(N__79827),
            .I(\c0.n9_adj_4552 ));
    Odrv12 I__19945 (
            .O(N__79824),
            .I(\c0.n9_adj_4552 ));
    Odrv12 I__19944 (
            .O(N__79821),
            .I(\c0.n9_adj_4552 ));
    Odrv4 I__19943 (
            .O(N__79814),
            .I(\c0.n9_adj_4552 ));
    Odrv4 I__19942 (
            .O(N__79811),
            .I(\c0.n9_adj_4552 ));
    CascadeMux I__19941 (
            .O(N__79800),
            .I(N__79797));
    InMux I__19940 (
            .O(N__79797),
            .I(N__79793));
    CascadeMux I__19939 (
            .O(N__79796),
            .I(N__79788));
    LocalMux I__19938 (
            .O(N__79793),
            .I(N__79781));
    InMux I__19937 (
            .O(N__79792),
            .I(N__79778));
    InMux I__19936 (
            .O(N__79791),
            .I(N__79769));
    InMux I__19935 (
            .O(N__79788),
            .I(N__79769));
    InMux I__19934 (
            .O(N__79787),
            .I(N__79769));
    InMux I__19933 (
            .O(N__79786),
            .I(N__79766));
    InMux I__19932 (
            .O(N__79785),
            .I(N__79763));
    InMux I__19931 (
            .O(N__79784),
            .I(N__79760));
    Span4Mux_h I__19930 (
            .O(N__79781),
            .I(N__79751));
    LocalMux I__19929 (
            .O(N__79778),
            .I(N__79751));
    InMux I__19928 (
            .O(N__79777),
            .I(N__79746));
    InMux I__19927 (
            .O(N__79776),
            .I(N__79746));
    LocalMux I__19926 (
            .O(N__79769),
            .I(N__79743));
    LocalMux I__19925 (
            .O(N__79766),
            .I(N__79740));
    LocalMux I__19924 (
            .O(N__79763),
            .I(N__79737));
    LocalMux I__19923 (
            .O(N__79760),
            .I(N__79734));
    InMux I__19922 (
            .O(N__79759),
            .I(N__79729));
    InMux I__19921 (
            .O(N__79758),
            .I(N__79729));
    InMux I__19920 (
            .O(N__79757),
            .I(N__79724));
    CascadeMux I__19919 (
            .O(N__79756),
            .I(N__79721));
    Span4Mux_v I__19918 (
            .O(N__79751),
            .I(N__79718));
    LocalMux I__19917 (
            .O(N__79746),
            .I(N__79709));
    Span4Mux_v I__19916 (
            .O(N__79743),
            .I(N__79709));
    Span4Mux_h I__19915 (
            .O(N__79740),
            .I(N__79709));
    Span4Mux_v I__19914 (
            .O(N__79737),
            .I(N__79709));
    Span4Mux_h I__19913 (
            .O(N__79734),
            .I(N__79704));
    LocalMux I__19912 (
            .O(N__79729),
            .I(N__79704));
    CascadeMux I__19911 (
            .O(N__79728),
            .I(N__79699));
    InMux I__19910 (
            .O(N__79727),
            .I(N__79695));
    LocalMux I__19909 (
            .O(N__79724),
            .I(N__79692));
    InMux I__19908 (
            .O(N__79721),
            .I(N__79689));
    Span4Mux_h I__19907 (
            .O(N__79718),
            .I(N__79686));
    Span4Mux_h I__19906 (
            .O(N__79709),
            .I(N__79681));
    Span4Mux_v I__19905 (
            .O(N__79704),
            .I(N__79681));
    InMux I__19904 (
            .O(N__79703),
            .I(N__79678));
    InMux I__19903 (
            .O(N__79702),
            .I(N__79674));
    InMux I__19902 (
            .O(N__79699),
            .I(N__79671));
    InMux I__19901 (
            .O(N__79698),
            .I(N__79668));
    LocalMux I__19900 (
            .O(N__79695),
            .I(N__79665));
    Span4Mux_h I__19899 (
            .O(N__79692),
            .I(N__79662));
    LocalMux I__19898 (
            .O(N__79689),
            .I(N__79653));
    Span4Mux_h I__19897 (
            .O(N__79686),
            .I(N__79653));
    Span4Mux_h I__19896 (
            .O(N__79681),
            .I(N__79653));
    LocalMux I__19895 (
            .O(N__79678),
            .I(N__79653));
    CascadeMux I__19894 (
            .O(N__79677),
            .I(N__79650));
    LocalMux I__19893 (
            .O(N__79674),
            .I(N__79641));
    LocalMux I__19892 (
            .O(N__79671),
            .I(N__79641));
    LocalMux I__19891 (
            .O(N__79668),
            .I(N__79632));
    Span4Mux_h I__19890 (
            .O(N__79665),
            .I(N__79632));
    Span4Mux_v I__19889 (
            .O(N__79662),
            .I(N__79632));
    Span4Mux_v I__19888 (
            .O(N__79653),
            .I(N__79632));
    InMux I__19887 (
            .O(N__79650),
            .I(N__79629));
    CascadeMux I__19886 (
            .O(N__79649),
            .I(N__79623));
    InMux I__19885 (
            .O(N__79648),
            .I(N__79619));
    InMux I__19884 (
            .O(N__79647),
            .I(N__79616));
    InMux I__19883 (
            .O(N__79646),
            .I(N__79613));
    Span4Mux_v I__19882 (
            .O(N__79641),
            .I(N__79608));
    Span4Mux_v I__19881 (
            .O(N__79632),
            .I(N__79608));
    LocalMux I__19880 (
            .O(N__79629),
            .I(N__79605));
    InMux I__19879 (
            .O(N__79628),
            .I(N__79602));
    InMux I__19878 (
            .O(N__79627),
            .I(N__79599));
    InMux I__19877 (
            .O(N__79626),
            .I(N__79596));
    InMux I__19876 (
            .O(N__79623),
            .I(N__79593));
    InMux I__19875 (
            .O(N__79622),
            .I(N__79590));
    LocalMux I__19874 (
            .O(N__79619),
            .I(N__79582));
    LocalMux I__19873 (
            .O(N__79616),
            .I(N__79582));
    LocalMux I__19872 (
            .O(N__79613),
            .I(N__79579));
    Span4Mux_h I__19871 (
            .O(N__79608),
            .I(N__79576));
    Span4Mux_h I__19870 (
            .O(N__79605),
            .I(N__79571));
    LocalMux I__19869 (
            .O(N__79602),
            .I(N__79571));
    LocalMux I__19868 (
            .O(N__79599),
            .I(N__79568));
    LocalMux I__19867 (
            .O(N__79596),
            .I(N__79565));
    LocalMux I__19866 (
            .O(N__79593),
            .I(N__79560));
    LocalMux I__19865 (
            .O(N__79590),
            .I(N__79560));
    InMux I__19864 (
            .O(N__79589),
            .I(N__79557));
    InMux I__19863 (
            .O(N__79588),
            .I(N__79554));
    InMux I__19862 (
            .O(N__79587),
            .I(N__79551));
    Span12Mux_h I__19861 (
            .O(N__79582),
            .I(N__79548));
    Span4Mux_h I__19860 (
            .O(N__79579),
            .I(N__79543));
    Span4Mux_v I__19859 (
            .O(N__79576),
            .I(N__79543));
    Sp12to4 I__19858 (
            .O(N__79571),
            .I(N__79537));
    Span12Mux_v I__19857 (
            .O(N__79568),
            .I(N__79537));
    Span12Mux_h I__19856 (
            .O(N__79565),
            .I(N__79532));
    Sp12to4 I__19855 (
            .O(N__79560),
            .I(N__79532));
    LocalMux I__19854 (
            .O(N__79557),
            .I(N__79527));
    LocalMux I__19853 (
            .O(N__79554),
            .I(N__79527));
    LocalMux I__19852 (
            .O(N__79551),
            .I(N__79522));
    Span12Mux_v I__19851 (
            .O(N__79548),
            .I(N__79522));
    Span4Mux_v I__19850 (
            .O(N__79543),
            .I(N__79519));
    InMux I__19849 (
            .O(N__79542),
            .I(N__79516));
    Span12Mux_v I__19848 (
            .O(N__79537),
            .I(N__79513));
    Span12Mux_v I__19847 (
            .O(N__79532),
            .I(N__79510));
    Span12Mux_h I__19846 (
            .O(N__79527),
            .I(N__79505));
    Span12Mux_h I__19845 (
            .O(N__79522),
            .I(N__79505));
    Span4Mux_v I__19844 (
            .O(N__79519),
            .I(N__79502));
    LocalMux I__19843 (
            .O(N__79516),
            .I(rx_data_5));
    Odrv12 I__19842 (
            .O(N__79513),
            .I(rx_data_5));
    Odrv12 I__19841 (
            .O(N__79510),
            .I(rx_data_5));
    Odrv12 I__19840 (
            .O(N__79505),
            .I(rx_data_5));
    Odrv4 I__19839 (
            .O(N__79502),
            .I(rx_data_5));
    InMux I__19838 (
            .O(N__79491),
            .I(N__79485));
    InMux I__19837 (
            .O(N__79490),
            .I(N__79478));
    InMux I__19836 (
            .O(N__79489),
            .I(N__79473));
    InMux I__19835 (
            .O(N__79488),
            .I(N__79468));
    LocalMux I__19834 (
            .O(N__79485),
            .I(N__79465));
    InMux I__19833 (
            .O(N__79484),
            .I(N__79458));
    InMux I__19832 (
            .O(N__79483),
            .I(N__79458));
    InMux I__19831 (
            .O(N__79482),
            .I(N__79453));
    InMux I__19830 (
            .O(N__79481),
            .I(N__79450));
    LocalMux I__19829 (
            .O(N__79478),
            .I(N__79447));
    CascadeMux I__19828 (
            .O(N__79477),
            .I(N__79444));
    InMux I__19827 (
            .O(N__79476),
            .I(N__79436));
    LocalMux I__19826 (
            .O(N__79473),
            .I(N__79433));
    InMux I__19825 (
            .O(N__79472),
            .I(N__79428));
    InMux I__19824 (
            .O(N__79471),
            .I(N__79428));
    LocalMux I__19823 (
            .O(N__79468),
            .I(N__79425));
    Span4Mux_h I__19822 (
            .O(N__79465),
            .I(N__79422));
    InMux I__19821 (
            .O(N__79464),
            .I(N__79415));
    InMux I__19820 (
            .O(N__79463),
            .I(N__79415));
    LocalMux I__19819 (
            .O(N__79458),
            .I(N__79412));
    InMux I__19818 (
            .O(N__79457),
            .I(N__79407));
    InMux I__19817 (
            .O(N__79456),
            .I(N__79407));
    LocalMux I__19816 (
            .O(N__79453),
            .I(N__79404));
    LocalMux I__19815 (
            .O(N__79450),
            .I(N__79399));
    Span4Mux_v I__19814 (
            .O(N__79447),
            .I(N__79399));
    InMux I__19813 (
            .O(N__79444),
            .I(N__79393));
    InMux I__19812 (
            .O(N__79443),
            .I(N__79388));
    InMux I__19811 (
            .O(N__79442),
            .I(N__79388));
    InMux I__19810 (
            .O(N__79441),
            .I(N__79385));
    InMux I__19809 (
            .O(N__79440),
            .I(N__79380));
    InMux I__19808 (
            .O(N__79439),
            .I(N__79380));
    LocalMux I__19807 (
            .O(N__79436),
            .I(N__79373));
    Span4Mux_v I__19806 (
            .O(N__79433),
            .I(N__79373));
    LocalMux I__19805 (
            .O(N__79428),
            .I(N__79373));
    Span4Mux_v I__19804 (
            .O(N__79425),
            .I(N__79370));
    Span4Mux_v I__19803 (
            .O(N__79422),
            .I(N__79367));
    InMux I__19802 (
            .O(N__79421),
            .I(N__79351));
    InMux I__19801 (
            .O(N__79420),
            .I(N__79348));
    LocalMux I__19800 (
            .O(N__79415),
            .I(N__79345));
    Span12Mux_s7_v I__19799 (
            .O(N__79412),
            .I(N__79342));
    LocalMux I__19798 (
            .O(N__79407),
            .I(N__79337));
    Span4Mux_v I__19797 (
            .O(N__79404),
            .I(N__79337));
    Span4Mux_h I__19796 (
            .O(N__79399),
            .I(N__79334));
    InMux I__19795 (
            .O(N__79398),
            .I(N__79327));
    InMux I__19794 (
            .O(N__79397),
            .I(N__79327));
    InMux I__19793 (
            .O(N__79396),
            .I(N__79327));
    LocalMux I__19792 (
            .O(N__79393),
            .I(N__79324));
    LocalMux I__19791 (
            .O(N__79388),
            .I(N__79321));
    LocalMux I__19790 (
            .O(N__79385),
            .I(N__79316));
    LocalMux I__19789 (
            .O(N__79380),
            .I(N__79316));
    Span4Mux_v I__19788 (
            .O(N__79373),
            .I(N__79311));
    Span4Mux_h I__19787 (
            .O(N__79370),
            .I(N__79311));
    Span4Mux_v I__19786 (
            .O(N__79367),
            .I(N__79308));
    InMux I__19785 (
            .O(N__79366),
            .I(N__79305));
    InMux I__19784 (
            .O(N__79365),
            .I(N__79300));
    InMux I__19783 (
            .O(N__79364),
            .I(N__79300));
    InMux I__19782 (
            .O(N__79363),
            .I(N__79295));
    InMux I__19781 (
            .O(N__79362),
            .I(N__79295));
    InMux I__19780 (
            .O(N__79361),
            .I(N__79288));
    InMux I__19779 (
            .O(N__79360),
            .I(N__79288));
    InMux I__19778 (
            .O(N__79359),
            .I(N__79288));
    InMux I__19777 (
            .O(N__79358),
            .I(N__79277));
    InMux I__19776 (
            .O(N__79357),
            .I(N__79277));
    InMux I__19775 (
            .O(N__79356),
            .I(N__79277));
    InMux I__19774 (
            .O(N__79355),
            .I(N__79277));
    InMux I__19773 (
            .O(N__79354),
            .I(N__79277));
    LocalMux I__19772 (
            .O(N__79351),
            .I(N__79274));
    LocalMux I__19771 (
            .O(N__79348),
            .I(N__79269));
    Span4Mux_v I__19770 (
            .O(N__79345),
            .I(N__79269));
    Span12Mux_v I__19769 (
            .O(N__79342),
            .I(N__79266));
    Span4Mux_h I__19768 (
            .O(N__79337),
            .I(N__79261));
    Span4Mux_h I__19767 (
            .O(N__79334),
            .I(N__79261));
    LocalMux I__19766 (
            .O(N__79327),
            .I(N__79248));
    Span4Mux_v I__19765 (
            .O(N__79324),
            .I(N__79248));
    Span4Mux_h I__19764 (
            .O(N__79321),
            .I(N__79248));
    Span4Mux_v I__19763 (
            .O(N__79316),
            .I(N__79248));
    Span4Mux_h I__19762 (
            .O(N__79311),
            .I(N__79248));
    Span4Mux_h I__19761 (
            .O(N__79308),
            .I(N__79248));
    LocalMux I__19760 (
            .O(N__79305),
            .I(\c0.n22134 ));
    LocalMux I__19759 (
            .O(N__79300),
            .I(\c0.n22134 ));
    LocalMux I__19758 (
            .O(N__79295),
            .I(\c0.n22134 ));
    LocalMux I__19757 (
            .O(N__79288),
            .I(\c0.n22134 ));
    LocalMux I__19756 (
            .O(N__79277),
            .I(\c0.n22134 ));
    Odrv4 I__19755 (
            .O(N__79274),
            .I(\c0.n22134 ));
    Odrv4 I__19754 (
            .O(N__79269),
            .I(\c0.n22134 ));
    Odrv12 I__19753 (
            .O(N__79266),
            .I(\c0.n22134 ));
    Odrv4 I__19752 (
            .O(N__79261),
            .I(\c0.n22134 ));
    Odrv4 I__19751 (
            .O(N__79248),
            .I(\c0.n22134 ));
    CascadeMux I__19750 (
            .O(N__79227),
            .I(N__79223));
    InMux I__19749 (
            .O(N__79226),
            .I(N__79220));
    InMux I__19748 (
            .O(N__79223),
            .I(N__79217));
    LocalMux I__19747 (
            .O(N__79220),
            .I(N__79214));
    LocalMux I__19746 (
            .O(N__79217),
            .I(\c0.data_in_frame_28_5 ));
    Odrv4 I__19745 (
            .O(N__79214),
            .I(\c0.data_in_frame_28_5 ));
    InMux I__19744 (
            .O(N__79209),
            .I(N__79206));
    LocalMux I__19743 (
            .O(N__79206),
            .I(N__79200));
    InMux I__19742 (
            .O(N__79205),
            .I(N__79197));
    CascadeMux I__19741 (
            .O(N__79204),
            .I(N__79194));
    InMux I__19740 (
            .O(N__79203),
            .I(N__79186));
    Span4Mux_h I__19739 (
            .O(N__79200),
            .I(N__79177));
    LocalMux I__19738 (
            .O(N__79197),
            .I(N__79177));
    InMux I__19737 (
            .O(N__79194),
            .I(N__79174));
    CascadeMux I__19736 (
            .O(N__79193),
            .I(N__79169));
    InMux I__19735 (
            .O(N__79192),
            .I(N__79164));
    CascadeMux I__19734 (
            .O(N__79191),
            .I(N__79161));
    InMux I__19733 (
            .O(N__79190),
            .I(N__79158));
    InMux I__19732 (
            .O(N__79189),
            .I(N__79155));
    LocalMux I__19731 (
            .O(N__79186),
            .I(N__79152));
    InMux I__19730 (
            .O(N__79185),
            .I(N__79149));
    CascadeMux I__19729 (
            .O(N__79184),
            .I(N__79145));
    CascadeMux I__19728 (
            .O(N__79183),
            .I(N__79142));
    CascadeMux I__19727 (
            .O(N__79182),
            .I(N__79137));
    Span4Mux_v I__19726 (
            .O(N__79177),
            .I(N__79132));
    LocalMux I__19725 (
            .O(N__79174),
            .I(N__79132));
    InMux I__19724 (
            .O(N__79173),
            .I(N__79129));
    InMux I__19723 (
            .O(N__79172),
            .I(N__79126));
    InMux I__19722 (
            .O(N__79169),
            .I(N__79120));
    InMux I__19721 (
            .O(N__79168),
            .I(N__79120));
    InMux I__19720 (
            .O(N__79167),
            .I(N__79117));
    LocalMux I__19719 (
            .O(N__79164),
            .I(N__79114));
    InMux I__19718 (
            .O(N__79161),
            .I(N__79111));
    LocalMux I__19717 (
            .O(N__79158),
            .I(N__79101));
    LocalMux I__19716 (
            .O(N__79155),
            .I(N__79101));
    Span4Mux_h I__19715 (
            .O(N__79152),
            .I(N__79096));
    LocalMux I__19714 (
            .O(N__79149),
            .I(N__79096));
    InMux I__19713 (
            .O(N__79148),
            .I(N__79093));
    InMux I__19712 (
            .O(N__79145),
            .I(N__79088));
    InMux I__19711 (
            .O(N__79142),
            .I(N__79088));
    CascadeMux I__19710 (
            .O(N__79141),
            .I(N__79085));
    InMux I__19709 (
            .O(N__79140),
            .I(N__79078));
    InMux I__19708 (
            .O(N__79137),
            .I(N__79078));
    Span4Mux_h I__19707 (
            .O(N__79132),
            .I(N__79075));
    LocalMux I__19706 (
            .O(N__79129),
            .I(N__79072));
    LocalMux I__19705 (
            .O(N__79126),
            .I(N__79069));
    InMux I__19704 (
            .O(N__79125),
            .I(N__79066));
    LocalMux I__19703 (
            .O(N__79120),
            .I(N__79063));
    LocalMux I__19702 (
            .O(N__79117),
            .I(N__79060));
    Span4Mux_v I__19701 (
            .O(N__79114),
            .I(N__79055));
    LocalMux I__19700 (
            .O(N__79111),
            .I(N__79055));
    InMux I__19699 (
            .O(N__79110),
            .I(N__79052));
    InMux I__19698 (
            .O(N__79109),
            .I(N__79046));
    InMux I__19697 (
            .O(N__79108),
            .I(N__79046));
    InMux I__19696 (
            .O(N__79107),
            .I(N__79043));
    InMux I__19695 (
            .O(N__79106),
            .I(N__79040));
    Span4Mux_v I__19694 (
            .O(N__79101),
            .I(N__79037));
    Span4Mux_h I__19693 (
            .O(N__79096),
            .I(N__79034));
    LocalMux I__19692 (
            .O(N__79093),
            .I(N__79029));
    LocalMux I__19691 (
            .O(N__79088),
            .I(N__79029));
    InMux I__19690 (
            .O(N__79085),
            .I(N__79022));
    InMux I__19689 (
            .O(N__79084),
            .I(N__79022));
    InMux I__19688 (
            .O(N__79083),
            .I(N__79022));
    LocalMux I__19687 (
            .O(N__79078),
            .I(N__79019));
    Span4Mux_v I__19686 (
            .O(N__79075),
            .I(N__79016));
    Span4Mux_h I__19685 (
            .O(N__79072),
            .I(N__79009));
    Span4Mux_v I__19684 (
            .O(N__79069),
            .I(N__79009));
    LocalMux I__19683 (
            .O(N__79066),
            .I(N__79009));
    Span4Mux_v I__19682 (
            .O(N__79063),
            .I(N__79006));
    Span4Mux_v I__19681 (
            .O(N__79060),
            .I(N__79001));
    Span4Mux_h I__19680 (
            .O(N__79055),
            .I(N__79001));
    LocalMux I__19679 (
            .O(N__79052),
            .I(N__78998));
    CascadeMux I__19678 (
            .O(N__79051),
            .I(N__78995));
    LocalMux I__19677 (
            .O(N__79046),
            .I(N__78985));
    LocalMux I__19676 (
            .O(N__79043),
            .I(N__78985));
    LocalMux I__19675 (
            .O(N__79040),
            .I(N__78985));
    Sp12to4 I__19674 (
            .O(N__79037),
            .I(N__78985));
    Span4Mux_v I__19673 (
            .O(N__79034),
            .I(N__78980));
    Span4Mux_v I__19672 (
            .O(N__79029),
            .I(N__78980));
    LocalMux I__19671 (
            .O(N__79022),
            .I(N__78975));
    Span4Mux_h I__19670 (
            .O(N__79019),
            .I(N__78970));
    Span4Mux_v I__19669 (
            .O(N__79016),
            .I(N__78970));
    Span4Mux_v I__19668 (
            .O(N__79009),
            .I(N__78963));
    Span4Mux_v I__19667 (
            .O(N__79006),
            .I(N__78963));
    Span4Mux_v I__19666 (
            .O(N__79001),
            .I(N__78963));
    Span4Mux_h I__19665 (
            .O(N__78998),
            .I(N__78960));
    InMux I__19664 (
            .O(N__78995),
            .I(N__78955));
    InMux I__19663 (
            .O(N__78994),
            .I(N__78955));
    Span12Mux_h I__19662 (
            .O(N__78985),
            .I(N__78952));
    Sp12to4 I__19661 (
            .O(N__78980),
            .I(N__78949));
    InMux I__19660 (
            .O(N__78979),
            .I(N__78946));
    InMux I__19659 (
            .O(N__78978),
            .I(N__78943));
    Span4Mux_h I__19658 (
            .O(N__78975),
            .I(N__78938));
    Span4Mux_h I__19657 (
            .O(N__78970),
            .I(N__78938));
    Span4Mux_h I__19656 (
            .O(N__78963),
            .I(N__78933));
    Span4Mux_v I__19655 (
            .O(N__78960),
            .I(N__78933));
    LocalMux I__19654 (
            .O(N__78955),
            .I(N__78926));
    Span12Mux_v I__19653 (
            .O(N__78952),
            .I(N__78926));
    Span12Mux_v I__19652 (
            .O(N__78949),
            .I(N__78926));
    LocalMux I__19651 (
            .O(N__78946),
            .I(rx_data_2));
    LocalMux I__19650 (
            .O(N__78943),
            .I(rx_data_2));
    Odrv4 I__19649 (
            .O(N__78938),
            .I(rx_data_2));
    Odrv4 I__19648 (
            .O(N__78933),
            .I(rx_data_2));
    Odrv12 I__19647 (
            .O(N__78926),
            .I(rx_data_2));
    InMux I__19646 (
            .O(N__78915),
            .I(N__78912));
    LocalMux I__19645 (
            .O(N__78912),
            .I(N__78908));
    InMux I__19644 (
            .O(N__78911),
            .I(N__78905));
    Span4Mux_v I__19643 (
            .O(N__78908),
            .I(N__78901));
    LocalMux I__19642 (
            .O(N__78905),
            .I(N__78898));
    InMux I__19641 (
            .O(N__78904),
            .I(N__78892));
    Span4Mux_h I__19640 (
            .O(N__78901),
            .I(N__78887));
    Span4Mux_v I__19639 (
            .O(N__78898),
            .I(N__78884));
    InMux I__19638 (
            .O(N__78897),
            .I(N__78881));
    InMux I__19637 (
            .O(N__78896),
            .I(N__78876));
    InMux I__19636 (
            .O(N__78895),
            .I(N__78876));
    LocalMux I__19635 (
            .O(N__78892),
            .I(N__78873));
    InMux I__19634 (
            .O(N__78891),
            .I(N__78870));
    InMux I__19633 (
            .O(N__78890),
            .I(N__78867));
    Odrv4 I__19632 (
            .O(N__78887),
            .I(n22110));
    Odrv4 I__19631 (
            .O(N__78884),
            .I(n22110));
    LocalMux I__19630 (
            .O(N__78881),
            .I(n22110));
    LocalMux I__19629 (
            .O(N__78876),
            .I(n22110));
    Odrv12 I__19628 (
            .O(N__78873),
            .I(n22110));
    LocalMux I__19627 (
            .O(N__78870),
            .I(n22110));
    LocalMux I__19626 (
            .O(N__78867),
            .I(n22110));
    InMux I__19625 (
            .O(N__78852),
            .I(N__78849));
    LocalMux I__19624 (
            .O(N__78849),
            .I(N__78846));
    Span4Mux_h I__19623 (
            .O(N__78846),
            .I(N__78843));
    Span4Mux_v I__19622 (
            .O(N__78843),
            .I(N__78838));
    InMux I__19621 (
            .O(N__78842),
            .I(N__78833));
    InMux I__19620 (
            .O(N__78841),
            .I(N__78833));
    Span4Mux_v I__19619 (
            .O(N__78838),
            .I(N__78830));
    LocalMux I__19618 (
            .O(N__78833),
            .I(data_in_frame_22_2));
    Odrv4 I__19617 (
            .O(N__78830),
            .I(data_in_frame_22_2));
    ClkMux I__19616 (
            .O(N__78825),
            .I(N__78033));
    ClkMux I__19615 (
            .O(N__78824),
            .I(N__78033));
    ClkMux I__19614 (
            .O(N__78823),
            .I(N__78033));
    ClkMux I__19613 (
            .O(N__78822),
            .I(N__78033));
    ClkMux I__19612 (
            .O(N__78821),
            .I(N__78033));
    ClkMux I__19611 (
            .O(N__78820),
            .I(N__78033));
    ClkMux I__19610 (
            .O(N__78819),
            .I(N__78033));
    ClkMux I__19609 (
            .O(N__78818),
            .I(N__78033));
    ClkMux I__19608 (
            .O(N__78817),
            .I(N__78033));
    ClkMux I__19607 (
            .O(N__78816),
            .I(N__78033));
    ClkMux I__19606 (
            .O(N__78815),
            .I(N__78033));
    ClkMux I__19605 (
            .O(N__78814),
            .I(N__78033));
    ClkMux I__19604 (
            .O(N__78813),
            .I(N__78033));
    ClkMux I__19603 (
            .O(N__78812),
            .I(N__78033));
    ClkMux I__19602 (
            .O(N__78811),
            .I(N__78033));
    ClkMux I__19601 (
            .O(N__78810),
            .I(N__78033));
    ClkMux I__19600 (
            .O(N__78809),
            .I(N__78033));
    ClkMux I__19599 (
            .O(N__78808),
            .I(N__78033));
    ClkMux I__19598 (
            .O(N__78807),
            .I(N__78033));
    ClkMux I__19597 (
            .O(N__78806),
            .I(N__78033));
    ClkMux I__19596 (
            .O(N__78805),
            .I(N__78033));
    ClkMux I__19595 (
            .O(N__78804),
            .I(N__78033));
    ClkMux I__19594 (
            .O(N__78803),
            .I(N__78033));
    ClkMux I__19593 (
            .O(N__78802),
            .I(N__78033));
    ClkMux I__19592 (
            .O(N__78801),
            .I(N__78033));
    ClkMux I__19591 (
            .O(N__78800),
            .I(N__78033));
    ClkMux I__19590 (
            .O(N__78799),
            .I(N__78033));
    ClkMux I__19589 (
            .O(N__78798),
            .I(N__78033));
    ClkMux I__19588 (
            .O(N__78797),
            .I(N__78033));
    ClkMux I__19587 (
            .O(N__78796),
            .I(N__78033));
    ClkMux I__19586 (
            .O(N__78795),
            .I(N__78033));
    ClkMux I__19585 (
            .O(N__78794),
            .I(N__78033));
    ClkMux I__19584 (
            .O(N__78793),
            .I(N__78033));
    ClkMux I__19583 (
            .O(N__78792),
            .I(N__78033));
    ClkMux I__19582 (
            .O(N__78791),
            .I(N__78033));
    ClkMux I__19581 (
            .O(N__78790),
            .I(N__78033));
    ClkMux I__19580 (
            .O(N__78789),
            .I(N__78033));
    ClkMux I__19579 (
            .O(N__78788),
            .I(N__78033));
    ClkMux I__19578 (
            .O(N__78787),
            .I(N__78033));
    ClkMux I__19577 (
            .O(N__78786),
            .I(N__78033));
    ClkMux I__19576 (
            .O(N__78785),
            .I(N__78033));
    ClkMux I__19575 (
            .O(N__78784),
            .I(N__78033));
    ClkMux I__19574 (
            .O(N__78783),
            .I(N__78033));
    ClkMux I__19573 (
            .O(N__78782),
            .I(N__78033));
    ClkMux I__19572 (
            .O(N__78781),
            .I(N__78033));
    ClkMux I__19571 (
            .O(N__78780),
            .I(N__78033));
    ClkMux I__19570 (
            .O(N__78779),
            .I(N__78033));
    ClkMux I__19569 (
            .O(N__78778),
            .I(N__78033));
    ClkMux I__19568 (
            .O(N__78777),
            .I(N__78033));
    ClkMux I__19567 (
            .O(N__78776),
            .I(N__78033));
    ClkMux I__19566 (
            .O(N__78775),
            .I(N__78033));
    ClkMux I__19565 (
            .O(N__78774),
            .I(N__78033));
    ClkMux I__19564 (
            .O(N__78773),
            .I(N__78033));
    ClkMux I__19563 (
            .O(N__78772),
            .I(N__78033));
    ClkMux I__19562 (
            .O(N__78771),
            .I(N__78033));
    ClkMux I__19561 (
            .O(N__78770),
            .I(N__78033));
    ClkMux I__19560 (
            .O(N__78769),
            .I(N__78033));
    ClkMux I__19559 (
            .O(N__78768),
            .I(N__78033));
    ClkMux I__19558 (
            .O(N__78767),
            .I(N__78033));
    ClkMux I__19557 (
            .O(N__78766),
            .I(N__78033));
    ClkMux I__19556 (
            .O(N__78765),
            .I(N__78033));
    ClkMux I__19555 (
            .O(N__78764),
            .I(N__78033));
    ClkMux I__19554 (
            .O(N__78763),
            .I(N__78033));
    ClkMux I__19553 (
            .O(N__78762),
            .I(N__78033));
    ClkMux I__19552 (
            .O(N__78761),
            .I(N__78033));
    ClkMux I__19551 (
            .O(N__78760),
            .I(N__78033));
    ClkMux I__19550 (
            .O(N__78759),
            .I(N__78033));
    ClkMux I__19549 (
            .O(N__78758),
            .I(N__78033));
    ClkMux I__19548 (
            .O(N__78757),
            .I(N__78033));
    ClkMux I__19547 (
            .O(N__78756),
            .I(N__78033));
    ClkMux I__19546 (
            .O(N__78755),
            .I(N__78033));
    ClkMux I__19545 (
            .O(N__78754),
            .I(N__78033));
    ClkMux I__19544 (
            .O(N__78753),
            .I(N__78033));
    ClkMux I__19543 (
            .O(N__78752),
            .I(N__78033));
    ClkMux I__19542 (
            .O(N__78751),
            .I(N__78033));
    ClkMux I__19541 (
            .O(N__78750),
            .I(N__78033));
    ClkMux I__19540 (
            .O(N__78749),
            .I(N__78033));
    ClkMux I__19539 (
            .O(N__78748),
            .I(N__78033));
    ClkMux I__19538 (
            .O(N__78747),
            .I(N__78033));
    ClkMux I__19537 (
            .O(N__78746),
            .I(N__78033));
    ClkMux I__19536 (
            .O(N__78745),
            .I(N__78033));
    ClkMux I__19535 (
            .O(N__78744),
            .I(N__78033));
    ClkMux I__19534 (
            .O(N__78743),
            .I(N__78033));
    ClkMux I__19533 (
            .O(N__78742),
            .I(N__78033));
    ClkMux I__19532 (
            .O(N__78741),
            .I(N__78033));
    ClkMux I__19531 (
            .O(N__78740),
            .I(N__78033));
    ClkMux I__19530 (
            .O(N__78739),
            .I(N__78033));
    ClkMux I__19529 (
            .O(N__78738),
            .I(N__78033));
    ClkMux I__19528 (
            .O(N__78737),
            .I(N__78033));
    ClkMux I__19527 (
            .O(N__78736),
            .I(N__78033));
    ClkMux I__19526 (
            .O(N__78735),
            .I(N__78033));
    ClkMux I__19525 (
            .O(N__78734),
            .I(N__78033));
    ClkMux I__19524 (
            .O(N__78733),
            .I(N__78033));
    ClkMux I__19523 (
            .O(N__78732),
            .I(N__78033));
    ClkMux I__19522 (
            .O(N__78731),
            .I(N__78033));
    ClkMux I__19521 (
            .O(N__78730),
            .I(N__78033));
    ClkMux I__19520 (
            .O(N__78729),
            .I(N__78033));
    ClkMux I__19519 (
            .O(N__78728),
            .I(N__78033));
    ClkMux I__19518 (
            .O(N__78727),
            .I(N__78033));
    ClkMux I__19517 (
            .O(N__78726),
            .I(N__78033));
    ClkMux I__19516 (
            .O(N__78725),
            .I(N__78033));
    ClkMux I__19515 (
            .O(N__78724),
            .I(N__78033));
    ClkMux I__19514 (
            .O(N__78723),
            .I(N__78033));
    ClkMux I__19513 (
            .O(N__78722),
            .I(N__78033));
    ClkMux I__19512 (
            .O(N__78721),
            .I(N__78033));
    ClkMux I__19511 (
            .O(N__78720),
            .I(N__78033));
    ClkMux I__19510 (
            .O(N__78719),
            .I(N__78033));
    ClkMux I__19509 (
            .O(N__78718),
            .I(N__78033));
    ClkMux I__19508 (
            .O(N__78717),
            .I(N__78033));
    ClkMux I__19507 (
            .O(N__78716),
            .I(N__78033));
    ClkMux I__19506 (
            .O(N__78715),
            .I(N__78033));
    ClkMux I__19505 (
            .O(N__78714),
            .I(N__78033));
    ClkMux I__19504 (
            .O(N__78713),
            .I(N__78033));
    ClkMux I__19503 (
            .O(N__78712),
            .I(N__78033));
    ClkMux I__19502 (
            .O(N__78711),
            .I(N__78033));
    ClkMux I__19501 (
            .O(N__78710),
            .I(N__78033));
    ClkMux I__19500 (
            .O(N__78709),
            .I(N__78033));
    ClkMux I__19499 (
            .O(N__78708),
            .I(N__78033));
    ClkMux I__19498 (
            .O(N__78707),
            .I(N__78033));
    ClkMux I__19497 (
            .O(N__78706),
            .I(N__78033));
    ClkMux I__19496 (
            .O(N__78705),
            .I(N__78033));
    ClkMux I__19495 (
            .O(N__78704),
            .I(N__78033));
    ClkMux I__19494 (
            .O(N__78703),
            .I(N__78033));
    ClkMux I__19493 (
            .O(N__78702),
            .I(N__78033));
    ClkMux I__19492 (
            .O(N__78701),
            .I(N__78033));
    ClkMux I__19491 (
            .O(N__78700),
            .I(N__78033));
    ClkMux I__19490 (
            .O(N__78699),
            .I(N__78033));
    ClkMux I__19489 (
            .O(N__78698),
            .I(N__78033));
    ClkMux I__19488 (
            .O(N__78697),
            .I(N__78033));
    ClkMux I__19487 (
            .O(N__78696),
            .I(N__78033));
    ClkMux I__19486 (
            .O(N__78695),
            .I(N__78033));
    ClkMux I__19485 (
            .O(N__78694),
            .I(N__78033));
    ClkMux I__19484 (
            .O(N__78693),
            .I(N__78033));
    ClkMux I__19483 (
            .O(N__78692),
            .I(N__78033));
    ClkMux I__19482 (
            .O(N__78691),
            .I(N__78033));
    ClkMux I__19481 (
            .O(N__78690),
            .I(N__78033));
    ClkMux I__19480 (
            .O(N__78689),
            .I(N__78033));
    ClkMux I__19479 (
            .O(N__78688),
            .I(N__78033));
    ClkMux I__19478 (
            .O(N__78687),
            .I(N__78033));
    ClkMux I__19477 (
            .O(N__78686),
            .I(N__78033));
    ClkMux I__19476 (
            .O(N__78685),
            .I(N__78033));
    ClkMux I__19475 (
            .O(N__78684),
            .I(N__78033));
    ClkMux I__19474 (
            .O(N__78683),
            .I(N__78033));
    ClkMux I__19473 (
            .O(N__78682),
            .I(N__78033));
    ClkMux I__19472 (
            .O(N__78681),
            .I(N__78033));
    ClkMux I__19471 (
            .O(N__78680),
            .I(N__78033));
    ClkMux I__19470 (
            .O(N__78679),
            .I(N__78033));
    ClkMux I__19469 (
            .O(N__78678),
            .I(N__78033));
    ClkMux I__19468 (
            .O(N__78677),
            .I(N__78033));
    ClkMux I__19467 (
            .O(N__78676),
            .I(N__78033));
    ClkMux I__19466 (
            .O(N__78675),
            .I(N__78033));
    ClkMux I__19465 (
            .O(N__78674),
            .I(N__78033));
    ClkMux I__19464 (
            .O(N__78673),
            .I(N__78033));
    ClkMux I__19463 (
            .O(N__78672),
            .I(N__78033));
    ClkMux I__19462 (
            .O(N__78671),
            .I(N__78033));
    ClkMux I__19461 (
            .O(N__78670),
            .I(N__78033));
    ClkMux I__19460 (
            .O(N__78669),
            .I(N__78033));
    ClkMux I__19459 (
            .O(N__78668),
            .I(N__78033));
    ClkMux I__19458 (
            .O(N__78667),
            .I(N__78033));
    ClkMux I__19457 (
            .O(N__78666),
            .I(N__78033));
    ClkMux I__19456 (
            .O(N__78665),
            .I(N__78033));
    ClkMux I__19455 (
            .O(N__78664),
            .I(N__78033));
    ClkMux I__19454 (
            .O(N__78663),
            .I(N__78033));
    ClkMux I__19453 (
            .O(N__78662),
            .I(N__78033));
    ClkMux I__19452 (
            .O(N__78661),
            .I(N__78033));
    ClkMux I__19451 (
            .O(N__78660),
            .I(N__78033));
    ClkMux I__19450 (
            .O(N__78659),
            .I(N__78033));
    ClkMux I__19449 (
            .O(N__78658),
            .I(N__78033));
    ClkMux I__19448 (
            .O(N__78657),
            .I(N__78033));
    ClkMux I__19447 (
            .O(N__78656),
            .I(N__78033));
    ClkMux I__19446 (
            .O(N__78655),
            .I(N__78033));
    ClkMux I__19445 (
            .O(N__78654),
            .I(N__78033));
    ClkMux I__19444 (
            .O(N__78653),
            .I(N__78033));
    ClkMux I__19443 (
            .O(N__78652),
            .I(N__78033));
    ClkMux I__19442 (
            .O(N__78651),
            .I(N__78033));
    ClkMux I__19441 (
            .O(N__78650),
            .I(N__78033));
    ClkMux I__19440 (
            .O(N__78649),
            .I(N__78033));
    ClkMux I__19439 (
            .O(N__78648),
            .I(N__78033));
    ClkMux I__19438 (
            .O(N__78647),
            .I(N__78033));
    ClkMux I__19437 (
            .O(N__78646),
            .I(N__78033));
    ClkMux I__19436 (
            .O(N__78645),
            .I(N__78033));
    ClkMux I__19435 (
            .O(N__78644),
            .I(N__78033));
    ClkMux I__19434 (
            .O(N__78643),
            .I(N__78033));
    ClkMux I__19433 (
            .O(N__78642),
            .I(N__78033));
    ClkMux I__19432 (
            .O(N__78641),
            .I(N__78033));
    ClkMux I__19431 (
            .O(N__78640),
            .I(N__78033));
    ClkMux I__19430 (
            .O(N__78639),
            .I(N__78033));
    ClkMux I__19429 (
            .O(N__78638),
            .I(N__78033));
    ClkMux I__19428 (
            .O(N__78637),
            .I(N__78033));
    ClkMux I__19427 (
            .O(N__78636),
            .I(N__78033));
    ClkMux I__19426 (
            .O(N__78635),
            .I(N__78033));
    ClkMux I__19425 (
            .O(N__78634),
            .I(N__78033));
    ClkMux I__19424 (
            .O(N__78633),
            .I(N__78033));
    ClkMux I__19423 (
            .O(N__78632),
            .I(N__78033));
    ClkMux I__19422 (
            .O(N__78631),
            .I(N__78033));
    ClkMux I__19421 (
            .O(N__78630),
            .I(N__78033));
    ClkMux I__19420 (
            .O(N__78629),
            .I(N__78033));
    ClkMux I__19419 (
            .O(N__78628),
            .I(N__78033));
    ClkMux I__19418 (
            .O(N__78627),
            .I(N__78033));
    ClkMux I__19417 (
            .O(N__78626),
            .I(N__78033));
    ClkMux I__19416 (
            .O(N__78625),
            .I(N__78033));
    ClkMux I__19415 (
            .O(N__78624),
            .I(N__78033));
    ClkMux I__19414 (
            .O(N__78623),
            .I(N__78033));
    ClkMux I__19413 (
            .O(N__78622),
            .I(N__78033));
    ClkMux I__19412 (
            .O(N__78621),
            .I(N__78033));
    ClkMux I__19411 (
            .O(N__78620),
            .I(N__78033));
    ClkMux I__19410 (
            .O(N__78619),
            .I(N__78033));
    ClkMux I__19409 (
            .O(N__78618),
            .I(N__78033));
    ClkMux I__19408 (
            .O(N__78617),
            .I(N__78033));
    ClkMux I__19407 (
            .O(N__78616),
            .I(N__78033));
    ClkMux I__19406 (
            .O(N__78615),
            .I(N__78033));
    ClkMux I__19405 (
            .O(N__78614),
            .I(N__78033));
    ClkMux I__19404 (
            .O(N__78613),
            .I(N__78033));
    ClkMux I__19403 (
            .O(N__78612),
            .I(N__78033));
    ClkMux I__19402 (
            .O(N__78611),
            .I(N__78033));
    ClkMux I__19401 (
            .O(N__78610),
            .I(N__78033));
    ClkMux I__19400 (
            .O(N__78609),
            .I(N__78033));
    ClkMux I__19399 (
            .O(N__78608),
            .I(N__78033));
    ClkMux I__19398 (
            .O(N__78607),
            .I(N__78033));
    ClkMux I__19397 (
            .O(N__78606),
            .I(N__78033));
    ClkMux I__19396 (
            .O(N__78605),
            .I(N__78033));
    ClkMux I__19395 (
            .O(N__78604),
            .I(N__78033));
    ClkMux I__19394 (
            .O(N__78603),
            .I(N__78033));
    ClkMux I__19393 (
            .O(N__78602),
            .I(N__78033));
    ClkMux I__19392 (
            .O(N__78601),
            .I(N__78033));
    ClkMux I__19391 (
            .O(N__78600),
            .I(N__78033));
    ClkMux I__19390 (
            .O(N__78599),
            .I(N__78033));
    ClkMux I__19389 (
            .O(N__78598),
            .I(N__78033));
    ClkMux I__19388 (
            .O(N__78597),
            .I(N__78033));
    ClkMux I__19387 (
            .O(N__78596),
            .I(N__78033));
    ClkMux I__19386 (
            .O(N__78595),
            .I(N__78033));
    ClkMux I__19385 (
            .O(N__78594),
            .I(N__78033));
    ClkMux I__19384 (
            .O(N__78593),
            .I(N__78033));
    ClkMux I__19383 (
            .O(N__78592),
            .I(N__78033));
    ClkMux I__19382 (
            .O(N__78591),
            .I(N__78033));
    ClkMux I__19381 (
            .O(N__78590),
            .I(N__78033));
    ClkMux I__19380 (
            .O(N__78589),
            .I(N__78033));
    ClkMux I__19379 (
            .O(N__78588),
            .I(N__78033));
    ClkMux I__19378 (
            .O(N__78587),
            .I(N__78033));
    ClkMux I__19377 (
            .O(N__78586),
            .I(N__78033));
    ClkMux I__19376 (
            .O(N__78585),
            .I(N__78033));
    ClkMux I__19375 (
            .O(N__78584),
            .I(N__78033));
    ClkMux I__19374 (
            .O(N__78583),
            .I(N__78033));
    ClkMux I__19373 (
            .O(N__78582),
            .I(N__78033));
    ClkMux I__19372 (
            .O(N__78581),
            .I(N__78033));
    ClkMux I__19371 (
            .O(N__78580),
            .I(N__78033));
    ClkMux I__19370 (
            .O(N__78579),
            .I(N__78033));
    ClkMux I__19369 (
            .O(N__78578),
            .I(N__78033));
    ClkMux I__19368 (
            .O(N__78577),
            .I(N__78033));
    ClkMux I__19367 (
            .O(N__78576),
            .I(N__78033));
    ClkMux I__19366 (
            .O(N__78575),
            .I(N__78033));
    ClkMux I__19365 (
            .O(N__78574),
            .I(N__78033));
    ClkMux I__19364 (
            .O(N__78573),
            .I(N__78033));
    ClkMux I__19363 (
            .O(N__78572),
            .I(N__78033));
    ClkMux I__19362 (
            .O(N__78571),
            .I(N__78033));
    ClkMux I__19361 (
            .O(N__78570),
            .I(N__78033));
    ClkMux I__19360 (
            .O(N__78569),
            .I(N__78033));
    ClkMux I__19359 (
            .O(N__78568),
            .I(N__78033));
    ClkMux I__19358 (
            .O(N__78567),
            .I(N__78033));
    ClkMux I__19357 (
            .O(N__78566),
            .I(N__78033));
    ClkMux I__19356 (
            .O(N__78565),
            .I(N__78033));
    ClkMux I__19355 (
            .O(N__78564),
            .I(N__78033));
    ClkMux I__19354 (
            .O(N__78563),
            .I(N__78033));
    ClkMux I__19353 (
            .O(N__78562),
            .I(N__78033));
    GlobalMux I__19352 (
            .O(N__78033),
            .I(N__78030));
    gio2CtrlBuf I__19351 (
            .O(N__78030),
            .I(CLK_c));
    InMux I__19350 (
            .O(N__78027),
            .I(N__78021));
    InMux I__19349 (
            .O(N__78026),
            .I(N__78014));
    InMux I__19348 (
            .O(N__78025),
            .I(N__78009));
    InMux I__19347 (
            .O(N__78024),
            .I(N__78009));
    LocalMux I__19346 (
            .O(N__78021),
            .I(N__78006));
    InMux I__19345 (
            .O(N__78020),
            .I(N__78003));
    InMux I__19344 (
            .O(N__78019),
            .I(N__77998));
    InMux I__19343 (
            .O(N__78018),
            .I(N__77998));
    CascadeMux I__19342 (
            .O(N__78017),
            .I(N__77995));
    LocalMux I__19341 (
            .O(N__78014),
            .I(N__77992));
    LocalMux I__19340 (
            .O(N__78009),
            .I(N__77987));
    Span4Mux_v I__19339 (
            .O(N__78006),
            .I(N__77987));
    LocalMux I__19338 (
            .O(N__78003),
            .I(N__77982));
    LocalMux I__19337 (
            .O(N__77998),
            .I(N__77982));
    InMux I__19336 (
            .O(N__77995),
            .I(N__77979));
    Span4Mux_v I__19335 (
            .O(N__77992),
            .I(N__77976));
    Span4Mux_h I__19334 (
            .O(N__77987),
            .I(N__77971));
    Span4Mux_v I__19333 (
            .O(N__77982),
            .I(N__77971));
    LocalMux I__19332 (
            .O(N__77979),
            .I(N__77966));
    Span4Mux_h I__19331 (
            .O(N__77976),
            .I(N__77966));
    Span4Mux_h I__19330 (
            .O(N__77971),
            .I(N__77963));
    Odrv4 I__19329 (
            .O(N__77966),
            .I(\c0.data_in_frame_24_0 ));
    Odrv4 I__19328 (
            .O(N__77963),
            .I(\c0.data_in_frame_24_0 ));
    InMux I__19327 (
            .O(N__77958),
            .I(N__77951));
    InMux I__19326 (
            .O(N__77957),
            .I(N__77948));
    InMux I__19325 (
            .O(N__77956),
            .I(N__77945));
    InMux I__19324 (
            .O(N__77955),
            .I(N__77942));
    InMux I__19323 (
            .O(N__77954),
            .I(N__77939));
    LocalMux I__19322 (
            .O(N__77951),
            .I(N__77933));
    LocalMux I__19321 (
            .O(N__77948),
            .I(N__77933));
    LocalMux I__19320 (
            .O(N__77945),
            .I(N__77928));
    LocalMux I__19319 (
            .O(N__77942),
            .I(N__77928));
    LocalMux I__19318 (
            .O(N__77939),
            .I(N__77925));
    InMux I__19317 (
            .O(N__77938),
            .I(N__77922));
    Span4Mux_v I__19316 (
            .O(N__77933),
            .I(N__77919));
    Span4Mux_h I__19315 (
            .O(N__77928),
            .I(N__77914));
    Span4Mux_v I__19314 (
            .O(N__77925),
            .I(N__77914));
    LocalMux I__19313 (
            .O(N__77922),
            .I(N__77911));
    Span4Mux_v I__19312 (
            .O(N__77919),
            .I(N__77906));
    Span4Mux_v I__19311 (
            .O(N__77914),
            .I(N__77906));
    Span12Mux_h I__19310 (
            .O(N__77911),
            .I(N__77903));
    Odrv4 I__19309 (
            .O(N__77906),
            .I(\c0.n29_adj_4362 ));
    Odrv12 I__19308 (
            .O(N__77903),
            .I(\c0.n29_adj_4362 ));
    InMux I__19307 (
            .O(N__77898),
            .I(N__77895));
    LocalMux I__19306 (
            .O(N__77895),
            .I(N__77892));
    Span4Mux_v I__19305 (
            .O(N__77892),
            .I(N__77889));
    Span4Mux_h I__19304 (
            .O(N__77889),
            .I(N__77886));
    Odrv4 I__19303 (
            .O(N__77886),
            .I(\c0.n24_adj_4531 ));
    InMux I__19302 (
            .O(N__77883),
            .I(N__77880));
    LocalMux I__19301 (
            .O(N__77880),
            .I(N__77876));
    InMux I__19300 (
            .O(N__77879),
            .I(N__77873));
    Span4Mux_h I__19299 (
            .O(N__77876),
            .I(N__77869));
    LocalMux I__19298 (
            .O(N__77873),
            .I(N__77866));
    InMux I__19297 (
            .O(N__77872),
            .I(N__77863));
    Span4Mux_h I__19296 (
            .O(N__77869),
            .I(N__77858));
    Span4Mux_v I__19295 (
            .O(N__77866),
            .I(N__77858));
    LocalMux I__19294 (
            .O(N__77863),
            .I(N__77853));
    Span4Mux_v I__19293 (
            .O(N__77858),
            .I(N__77850));
    InMux I__19292 (
            .O(N__77857),
            .I(N__77847));
    InMux I__19291 (
            .O(N__77856),
            .I(N__77841));
    Span12Mux_v I__19290 (
            .O(N__77853),
            .I(N__77838));
    Span4Mux_h I__19289 (
            .O(N__77850),
            .I(N__77833));
    LocalMux I__19288 (
            .O(N__77847),
            .I(N__77833));
    InMux I__19287 (
            .O(N__77846),
            .I(N__77826));
    InMux I__19286 (
            .O(N__77845),
            .I(N__77826));
    InMux I__19285 (
            .O(N__77844),
            .I(N__77826));
    LocalMux I__19284 (
            .O(N__77841),
            .I(data_in_frame_6_3));
    Odrv12 I__19283 (
            .O(N__77838),
            .I(data_in_frame_6_3));
    Odrv4 I__19282 (
            .O(N__77833),
            .I(data_in_frame_6_3));
    LocalMux I__19281 (
            .O(N__77826),
            .I(data_in_frame_6_3));
    InMux I__19280 (
            .O(N__77817),
            .I(N__77813));
    InMux I__19279 (
            .O(N__77816),
            .I(N__77807));
    LocalMux I__19278 (
            .O(N__77813),
            .I(N__77804));
    InMux I__19277 (
            .O(N__77812),
            .I(N__77799));
    InMux I__19276 (
            .O(N__77811),
            .I(N__77799));
    InMux I__19275 (
            .O(N__77810),
            .I(N__77796));
    LocalMux I__19274 (
            .O(N__77807),
            .I(N__77793));
    Span4Mux_v I__19273 (
            .O(N__77804),
            .I(N__77789));
    LocalMux I__19272 (
            .O(N__77799),
            .I(N__77784));
    LocalMux I__19271 (
            .O(N__77796),
            .I(N__77784));
    Span4Mux_v I__19270 (
            .O(N__77793),
            .I(N__77781));
    InMux I__19269 (
            .O(N__77792),
            .I(N__77778));
    Span4Mux_h I__19268 (
            .O(N__77789),
            .I(N__77771));
    Span4Mux_v I__19267 (
            .O(N__77784),
            .I(N__77771));
    Span4Mux_v I__19266 (
            .O(N__77781),
            .I(N__77766));
    LocalMux I__19265 (
            .O(N__77778),
            .I(N__77766));
    InMux I__19264 (
            .O(N__77777),
            .I(N__77761));
    InMux I__19263 (
            .O(N__77776),
            .I(N__77761));
    Odrv4 I__19262 (
            .O(N__77771),
            .I(\c0.n23267 ));
    Odrv4 I__19261 (
            .O(N__77766),
            .I(\c0.n23267 ));
    LocalMux I__19260 (
            .O(N__77761),
            .I(\c0.n23267 ));
    CascadeMux I__19259 (
            .O(N__77754),
            .I(\c0.n18_cascade_ ));
    InMux I__19258 (
            .O(N__77751),
            .I(N__77748));
    LocalMux I__19257 (
            .O(N__77748),
            .I(N__77745));
    Span4Mux_h I__19256 (
            .O(N__77745),
            .I(N__77742));
    Odrv4 I__19255 (
            .O(N__77742),
            .I(\c0.n16_adj_4666 ));
    InMux I__19254 (
            .O(N__77739),
            .I(N__77736));
    LocalMux I__19253 (
            .O(N__77736),
            .I(\c0.n28_adj_4667 ));
    CascadeMux I__19252 (
            .O(N__77733),
            .I(\c0.n24_adj_4653_cascade_ ));
    InMux I__19251 (
            .O(N__77730),
            .I(N__77727));
    LocalMux I__19250 (
            .O(N__77727),
            .I(N__77723));
    InMux I__19249 (
            .O(N__77726),
            .I(N__77720));
    Span4Mux_v I__19248 (
            .O(N__77723),
            .I(N__77715));
    LocalMux I__19247 (
            .O(N__77720),
            .I(N__77715));
    Span4Mux_h I__19246 (
            .O(N__77715),
            .I(N__77712));
    Odrv4 I__19245 (
            .O(N__77712),
            .I(\c0.n22369 ));
    InMux I__19244 (
            .O(N__77709),
            .I(N__77706));
    LocalMux I__19243 (
            .O(N__77706),
            .I(N__77702));
    CascadeMux I__19242 (
            .O(N__77705),
            .I(N__77699));
    Span4Mux_h I__19241 (
            .O(N__77702),
            .I(N__77696));
    InMux I__19240 (
            .O(N__77699),
            .I(N__77693));
    Odrv4 I__19239 (
            .O(N__77696),
            .I(\c0.n6_adj_4587 ));
    LocalMux I__19238 (
            .O(N__77693),
            .I(\c0.n6_adj_4587 ));
    InMux I__19237 (
            .O(N__77688),
            .I(N__77684));
    InMux I__19236 (
            .O(N__77687),
            .I(N__77681));
    LocalMux I__19235 (
            .O(N__77684),
            .I(N__77678));
    LocalMux I__19234 (
            .O(N__77681),
            .I(N__77675));
    Span4Mux_h I__19233 (
            .O(N__77678),
            .I(N__77668));
    Span4Mux_h I__19232 (
            .O(N__77675),
            .I(N__77668));
    InMux I__19231 (
            .O(N__77674),
            .I(N__77663));
    InMux I__19230 (
            .O(N__77673),
            .I(N__77663));
    Span4Mux_h I__19229 (
            .O(N__77668),
            .I(N__77658));
    LocalMux I__19228 (
            .O(N__77663),
            .I(N__77658));
    Odrv4 I__19227 (
            .O(N__77658),
            .I(\c0.n22586 ));
    CascadeMux I__19226 (
            .O(N__77655),
            .I(N__77651));
    InMux I__19225 (
            .O(N__77654),
            .I(N__77646));
    InMux I__19224 (
            .O(N__77651),
            .I(N__77643));
    InMux I__19223 (
            .O(N__77650),
            .I(N__77640));
    CascadeMux I__19222 (
            .O(N__77649),
            .I(N__77635));
    LocalMux I__19221 (
            .O(N__77646),
            .I(N__77632));
    LocalMux I__19220 (
            .O(N__77643),
            .I(N__77629));
    LocalMux I__19219 (
            .O(N__77640),
            .I(N__77626));
    InMux I__19218 (
            .O(N__77639),
            .I(N__77623));
    InMux I__19217 (
            .O(N__77638),
            .I(N__77620));
    InMux I__19216 (
            .O(N__77635),
            .I(N__77617));
    Span4Mux_v I__19215 (
            .O(N__77632),
            .I(N__77614));
    Span4Mux_v I__19214 (
            .O(N__77629),
            .I(N__77611));
    Span4Mux_v I__19213 (
            .O(N__77626),
            .I(N__77608));
    LocalMux I__19212 (
            .O(N__77623),
            .I(N__77605));
    LocalMux I__19211 (
            .O(N__77620),
            .I(N__77602));
    LocalMux I__19210 (
            .O(N__77617),
            .I(N__77593));
    Span4Mux_h I__19209 (
            .O(N__77614),
            .I(N__77593));
    Span4Mux_v I__19208 (
            .O(N__77611),
            .I(N__77593));
    Span4Mux_v I__19207 (
            .O(N__77608),
            .I(N__77593));
    Span4Mux_v I__19206 (
            .O(N__77605),
            .I(N__77590));
    Odrv12 I__19205 (
            .O(N__77602),
            .I(\c0.data_in_frame_19_6 ));
    Odrv4 I__19204 (
            .O(N__77593),
            .I(\c0.data_in_frame_19_6 ));
    Odrv4 I__19203 (
            .O(N__77590),
            .I(\c0.data_in_frame_19_6 ));
    InMux I__19202 (
            .O(N__77583),
            .I(N__77580));
    LocalMux I__19201 (
            .O(N__77580),
            .I(N__77575));
    InMux I__19200 (
            .O(N__77579),
            .I(N__77570));
    InMux I__19199 (
            .O(N__77578),
            .I(N__77566));
    Span4Mux_v I__19198 (
            .O(N__77575),
            .I(N__77563));
    InMux I__19197 (
            .O(N__77574),
            .I(N__77560));
    InMux I__19196 (
            .O(N__77573),
            .I(N__77557));
    LocalMux I__19195 (
            .O(N__77570),
            .I(N__77554));
    CascadeMux I__19194 (
            .O(N__77569),
            .I(N__77551));
    LocalMux I__19193 (
            .O(N__77566),
            .I(N__77546));
    Span4Mux_h I__19192 (
            .O(N__77563),
            .I(N__77546));
    LocalMux I__19191 (
            .O(N__77560),
            .I(N__77543));
    LocalMux I__19190 (
            .O(N__77557),
            .I(N__77538));
    Span4Mux_h I__19189 (
            .O(N__77554),
            .I(N__77538));
    InMux I__19188 (
            .O(N__77551),
            .I(N__77535));
    Span4Mux_v I__19187 (
            .O(N__77546),
            .I(N__77532));
    Span4Mux_h I__19186 (
            .O(N__77543),
            .I(N__77529));
    Span4Mux_v I__19185 (
            .O(N__77538),
            .I(N__77526));
    LocalMux I__19184 (
            .O(N__77535),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__19183 (
            .O(N__77532),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__19182 (
            .O(N__77529),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__19181 (
            .O(N__77526),
            .I(\c0.data_in_frame_19_7 ));
    InMux I__19180 (
            .O(N__77517),
            .I(N__77514));
    LocalMux I__19179 (
            .O(N__77514),
            .I(N__77511));
    Odrv12 I__19178 (
            .O(N__77511),
            .I(\c0.n23433 ));
    InMux I__19177 (
            .O(N__77508),
            .I(N__77505));
    LocalMux I__19176 (
            .O(N__77505),
            .I(\c0.n15_adj_4625 ));
    InMux I__19175 (
            .O(N__77502),
            .I(N__77498));
    InMux I__19174 (
            .O(N__77501),
            .I(N__77495));
    LocalMux I__19173 (
            .O(N__77498),
            .I(\c0.n17_adj_4626 ));
    LocalMux I__19172 (
            .O(N__77495),
            .I(\c0.n17_adj_4626 ));
    InMux I__19171 (
            .O(N__77490),
            .I(N__77486));
    InMux I__19170 (
            .O(N__77489),
            .I(N__77483));
    LocalMux I__19169 (
            .O(N__77486),
            .I(N__77480));
    LocalMux I__19168 (
            .O(N__77483),
            .I(N__77477));
    Span4Mux_v I__19167 (
            .O(N__77480),
            .I(N__77474));
    Span4Mux_h I__19166 (
            .O(N__77477),
            .I(N__77471));
    Odrv4 I__19165 (
            .O(N__77474),
            .I(\c0.n16_adj_4627 ));
    Odrv4 I__19164 (
            .O(N__77471),
            .I(\c0.n16_adj_4627 ));
    CascadeMux I__19163 (
            .O(N__77466),
            .I(\c0.n15_adj_4625_cascade_ ));
    InMux I__19162 (
            .O(N__77463),
            .I(N__77460));
    LocalMux I__19161 (
            .O(N__77460),
            .I(\c0.n18 ));
    InMux I__19160 (
            .O(N__77457),
            .I(N__77454));
    LocalMux I__19159 (
            .O(N__77454),
            .I(N__77450));
    InMux I__19158 (
            .O(N__77453),
            .I(N__77447));
    Span4Mux_v I__19157 (
            .O(N__77450),
            .I(N__77441));
    LocalMux I__19156 (
            .O(N__77447),
            .I(N__77441));
    InMux I__19155 (
            .O(N__77446),
            .I(N__77437));
    Span4Mux_v I__19154 (
            .O(N__77441),
            .I(N__77434));
    InMux I__19153 (
            .O(N__77440),
            .I(N__77431));
    LocalMux I__19152 (
            .O(N__77437),
            .I(N__77428));
    Odrv4 I__19151 (
            .O(N__77434),
            .I(\c0.n22605 ));
    LocalMux I__19150 (
            .O(N__77431),
            .I(\c0.n22605 ));
    Odrv12 I__19149 (
            .O(N__77428),
            .I(\c0.n22605 ));
    InMux I__19148 (
            .O(N__77421),
            .I(N__77418));
    LocalMux I__19147 (
            .O(N__77418),
            .I(N__77414));
    InMux I__19146 (
            .O(N__77417),
            .I(N__77411));
    Span4Mux_v I__19145 (
            .O(N__77414),
            .I(N__77406));
    LocalMux I__19144 (
            .O(N__77411),
            .I(N__77406));
    Span4Mux_h I__19143 (
            .O(N__77406),
            .I(N__77402));
    InMux I__19142 (
            .O(N__77405),
            .I(N__77399));
    Odrv4 I__19141 (
            .O(N__77402),
            .I(\c0.n13767 ));
    LocalMux I__19140 (
            .O(N__77399),
            .I(\c0.n13767 ));
    CascadeMux I__19139 (
            .O(N__77394),
            .I(N__77388));
    InMux I__19138 (
            .O(N__77393),
            .I(N__77383));
    InMux I__19137 (
            .O(N__77392),
            .I(N__77383));
    InMux I__19136 (
            .O(N__77391),
            .I(N__77380));
    InMux I__19135 (
            .O(N__77388),
            .I(N__77377));
    LocalMux I__19134 (
            .O(N__77383),
            .I(N__77373));
    LocalMux I__19133 (
            .O(N__77380),
            .I(N__77368));
    LocalMux I__19132 (
            .O(N__77377),
            .I(N__77368));
    InMux I__19131 (
            .O(N__77376),
            .I(N__77365));
    Span4Mux_h I__19130 (
            .O(N__77373),
            .I(N__77362));
    Odrv4 I__19129 (
            .O(N__77368),
            .I(\c0.n13468 ));
    LocalMux I__19128 (
            .O(N__77365),
            .I(\c0.n13468 ));
    Odrv4 I__19127 (
            .O(N__77362),
            .I(\c0.n13468 ));
    CascadeMux I__19126 (
            .O(N__77355),
            .I(\c0.n20239_cascade_ ));
    InMux I__19125 (
            .O(N__77352),
            .I(N__77348));
    InMux I__19124 (
            .O(N__77351),
            .I(N__77345));
    LocalMux I__19123 (
            .O(N__77348),
            .I(N__77342));
    LocalMux I__19122 (
            .O(N__77345),
            .I(N__77336));
    Span4Mux_v I__19121 (
            .O(N__77342),
            .I(N__77336));
    InMux I__19120 (
            .O(N__77341),
            .I(N__77333));
    Span4Mux_h I__19119 (
            .O(N__77336),
            .I(N__77329));
    LocalMux I__19118 (
            .O(N__77333),
            .I(N__77326));
    CascadeMux I__19117 (
            .O(N__77332),
            .I(N__77323));
    Sp12to4 I__19116 (
            .O(N__77329),
            .I(N__77318));
    Sp12to4 I__19115 (
            .O(N__77326),
            .I(N__77318));
    InMux I__19114 (
            .O(N__77323),
            .I(N__77315));
    Span12Mux_s10_v I__19113 (
            .O(N__77318),
            .I(N__77312));
    LocalMux I__19112 (
            .O(N__77315),
            .I(\c0.data_in_frame_26_4 ));
    Odrv12 I__19111 (
            .O(N__77312),
            .I(\c0.data_in_frame_26_4 ));
    InMux I__19110 (
            .O(N__77307),
            .I(N__77304));
    LocalMux I__19109 (
            .O(N__77304),
            .I(N__77301));
    Odrv12 I__19108 (
            .O(N__77301),
            .I(\c0.n10_adj_4457 ));
    InMux I__19107 (
            .O(N__77298),
            .I(N__77295));
    LocalMux I__19106 (
            .O(N__77295),
            .I(\c0.n6_adj_4668 ));
    CascadeMux I__19105 (
            .O(N__77292),
            .I(N__77288));
    InMux I__19104 (
            .O(N__77291),
            .I(N__77284));
    InMux I__19103 (
            .O(N__77288),
            .I(N__77281));
    InMux I__19102 (
            .O(N__77287),
            .I(N__77277));
    LocalMux I__19101 (
            .O(N__77284),
            .I(N__77274));
    LocalMux I__19100 (
            .O(N__77281),
            .I(N__77270));
    InMux I__19099 (
            .O(N__77280),
            .I(N__77267));
    LocalMux I__19098 (
            .O(N__77277),
            .I(N__77261));
    Span4Mux_h I__19097 (
            .O(N__77274),
            .I(N__77261));
    InMux I__19096 (
            .O(N__77273),
            .I(N__77258));
    Span4Mux_v I__19095 (
            .O(N__77270),
            .I(N__77255));
    LocalMux I__19094 (
            .O(N__77267),
            .I(N__77252));
    InMux I__19093 (
            .O(N__77266),
            .I(N__77249));
    Span4Mux_h I__19092 (
            .O(N__77261),
            .I(N__77246));
    LocalMux I__19091 (
            .O(N__77258),
            .I(N__77243));
    Span4Mux_h I__19090 (
            .O(N__77255),
            .I(N__77238));
    Span4Mux_h I__19089 (
            .O(N__77252),
            .I(N__77238));
    LocalMux I__19088 (
            .O(N__77249),
            .I(\c0.data_in_frame_23_2 ));
    Odrv4 I__19087 (
            .O(N__77246),
            .I(\c0.data_in_frame_23_2 ));
    Odrv12 I__19086 (
            .O(N__77243),
            .I(\c0.data_in_frame_23_2 ));
    Odrv4 I__19085 (
            .O(N__77238),
            .I(\c0.data_in_frame_23_2 ));
    InMux I__19084 (
            .O(N__77229),
            .I(N__77226));
    LocalMux I__19083 (
            .O(N__77226),
            .I(N__77223));
    Span4Mux_h I__19082 (
            .O(N__77223),
            .I(N__77220));
    Odrv4 I__19081 (
            .O(N__77220),
            .I(\c0.n13314 ));
    InMux I__19080 (
            .O(N__77217),
            .I(N__77213));
    InMux I__19079 (
            .O(N__77216),
            .I(N__77210));
    LocalMux I__19078 (
            .O(N__77213),
            .I(N__77204));
    LocalMux I__19077 (
            .O(N__77210),
            .I(N__77204));
    CascadeMux I__19076 (
            .O(N__77209),
            .I(N__77201));
    Span4Mux_v I__19075 (
            .O(N__77204),
            .I(N__77198));
    InMux I__19074 (
            .O(N__77201),
            .I(N__77195));
    Odrv4 I__19073 (
            .O(N__77198),
            .I(\c0.n6227 ));
    LocalMux I__19072 (
            .O(N__77195),
            .I(\c0.n6227 ));
    InMux I__19071 (
            .O(N__77190),
            .I(N__77184));
    CascadeMux I__19070 (
            .O(N__77189),
            .I(N__77181));
    InMux I__19069 (
            .O(N__77188),
            .I(N__77177));
    InMux I__19068 (
            .O(N__77187),
            .I(N__77174));
    LocalMux I__19067 (
            .O(N__77184),
            .I(N__77171));
    InMux I__19066 (
            .O(N__77181),
            .I(N__77168));
    InMux I__19065 (
            .O(N__77180),
            .I(N__77165));
    LocalMux I__19064 (
            .O(N__77177),
            .I(N__77162));
    LocalMux I__19063 (
            .O(N__77174),
            .I(data_in_frame_21_7));
    Odrv4 I__19062 (
            .O(N__77171),
            .I(data_in_frame_21_7));
    LocalMux I__19061 (
            .O(N__77168),
            .I(data_in_frame_21_7));
    LocalMux I__19060 (
            .O(N__77165),
            .I(data_in_frame_21_7));
    Odrv4 I__19059 (
            .O(N__77162),
            .I(data_in_frame_21_7));
    InMux I__19058 (
            .O(N__77151),
            .I(N__77147));
    InMux I__19057 (
            .O(N__77150),
            .I(N__77144));
    LocalMux I__19056 (
            .O(N__77147),
            .I(N__77141));
    LocalMux I__19055 (
            .O(N__77144),
            .I(N__77138));
    Odrv4 I__19054 (
            .O(N__77141),
            .I(\c0.n20350 ));
    Odrv4 I__19053 (
            .O(N__77138),
            .I(\c0.n20350 ));
    CascadeMux I__19052 (
            .O(N__77133),
            .I(N__77125));
    CascadeMux I__19051 (
            .O(N__77132),
            .I(N__77118));
    InMux I__19050 (
            .O(N__77131),
            .I(N__77115));
    InMux I__19049 (
            .O(N__77130),
            .I(N__77112));
    InMux I__19048 (
            .O(N__77129),
            .I(N__77107));
    InMux I__19047 (
            .O(N__77128),
            .I(N__77103));
    InMux I__19046 (
            .O(N__77125),
            .I(N__77093));
    InMux I__19045 (
            .O(N__77124),
            .I(N__77093));
    InMux I__19044 (
            .O(N__77123),
            .I(N__77087));
    InMux I__19043 (
            .O(N__77122),
            .I(N__77084));
    CascadeMux I__19042 (
            .O(N__77121),
            .I(N__77081));
    InMux I__19041 (
            .O(N__77118),
            .I(N__77078));
    LocalMux I__19040 (
            .O(N__77115),
            .I(N__77075));
    LocalMux I__19039 (
            .O(N__77112),
            .I(N__77072));
    InMux I__19038 (
            .O(N__77111),
            .I(N__77069));
    InMux I__19037 (
            .O(N__77110),
            .I(N__77066));
    LocalMux I__19036 (
            .O(N__77107),
            .I(N__77062));
    InMux I__19035 (
            .O(N__77106),
            .I(N__77059));
    LocalMux I__19034 (
            .O(N__77103),
            .I(N__77055));
    InMux I__19033 (
            .O(N__77102),
            .I(N__77052));
    InMux I__19032 (
            .O(N__77101),
            .I(N__77049));
    InMux I__19031 (
            .O(N__77100),
            .I(N__77046));
    CascadeMux I__19030 (
            .O(N__77099),
            .I(N__77041));
    CascadeMux I__19029 (
            .O(N__77098),
            .I(N__77038));
    LocalMux I__19028 (
            .O(N__77093),
            .I(N__77035));
    InMux I__19027 (
            .O(N__77092),
            .I(N__77028));
    InMux I__19026 (
            .O(N__77091),
            .I(N__77028));
    InMux I__19025 (
            .O(N__77090),
            .I(N__77028));
    LocalMux I__19024 (
            .O(N__77087),
            .I(N__77023));
    LocalMux I__19023 (
            .O(N__77084),
            .I(N__77023));
    InMux I__19022 (
            .O(N__77081),
            .I(N__77020));
    LocalMux I__19021 (
            .O(N__77078),
            .I(N__77017));
    Span4Mux_h I__19020 (
            .O(N__77075),
            .I(N__77012));
    Span4Mux_h I__19019 (
            .O(N__77072),
            .I(N__77012));
    LocalMux I__19018 (
            .O(N__77069),
            .I(N__77009));
    LocalMux I__19017 (
            .O(N__77066),
            .I(N__77006));
    InMux I__19016 (
            .O(N__77065),
            .I(N__77003));
    Span4Mux_v I__19015 (
            .O(N__77062),
            .I(N__76998));
    LocalMux I__19014 (
            .O(N__77059),
            .I(N__76998));
    InMux I__19013 (
            .O(N__77058),
            .I(N__76994));
    Span4Mux_v I__19012 (
            .O(N__77055),
            .I(N__76985));
    LocalMux I__19011 (
            .O(N__77052),
            .I(N__76985));
    LocalMux I__19010 (
            .O(N__77049),
            .I(N__76985));
    LocalMux I__19009 (
            .O(N__77046),
            .I(N__76985));
    InMux I__19008 (
            .O(N__77045),
            .I(N__76982));
    InMux I__19007 (
            .O(N__77044),
            .I(N__76979));
    InMux I__19006 (
            .O(N__77041),
            .I(N__76974));
    InMux I__19005 (
            .O(N__77038),
            .I(N__76974));
    Span4Mux_v I__19004 (
            .O(N__77035),
            .I(N__76963));
    LocalMux I__19003 (
            .O(N__77028),
            .I(N__76963));
    Span4Mux_h I__19002 (
            .O(N__77023),
            .I(N__76963));
    LocalMux I__19001 (
            .O(N__77020),
            .I(N__76963));
    Span4Mux_v I__19000 (
            .O(N__77017),
            .I(N__76963));
    Span4Mux_h I__18999 (
            .O(N__77012),
            .I(N__76958));
    Span4Mux_v I__18998 (
            .O(N__77009),
            .I(N__76958));
    Span4Mux_v I__18997 (
            .O(N__77006),
            .I(N__76955));
    LocalMux I__18996 (
            .O(N__77003),
            .I(N__76949));
    Span4Mux_h I__18995 (
            .O(N__76998),
            .I(N__76949));
    InMux I__18994 (
            .O(N__76997),
            .I(N__76946));
    LocalMux I__18993 (
            .O(N__76994),
            .I(N__76941));
    Span4Mux_h I__18992 (
            .O(N__76985),
            .I(N__76936));
    LocalMux I__18991 (
            .O(N__76982),
            .I(N__76936));
    LocalMux I__18990 (
            .O(N__76979),
            .I(N__76933));
    LocalMux I__18989 (
            .O(N__76974),
            .I(N__76926));
    Span4Mux_h I__18988 (
            .O(N__76963),
            .I(N__76926));
    Span4Mux_v I__18987 (
            .O(N__76958),
            .I(N__76926));
    Span4Mux_v I__18986 (
            .O(N__76955),
            .I(N__76923));
    InMux I__18985 (
            .O(N__76954),
            .I(N__76920));
    Span4Mux_v I__18984 (
            .O(N__76949),
            .I(N__76917));
    LocalMux I__18983 (
            .O(N__76946),
            .I(N__76913));
    InMux I__18982 (
            .O(N__76945),
            .I(N__76909));
    InMux I__18981 (
            .O(N__76944),
            .I(N__76906));
    Span4Mux_v I__18980 (
            .O(N__76941),
            .I(N__76903));
    Span4Mux_h I__18979 (
            .O(N__76936),
            .I(N__76900));
    Span4Mux_h I__18978 (
            .O(N__76933),
            .I(N__76895));
    Span4Mux_v I__18977 (
            .O(N__76926),
            .I(N__76895));
    Span4Mux_v I__18976 (
            .O(N__76923),
            .I(N__76892));
    LocalMux I__18975 (
            .O(N__76920),
            .I(N__76887));
    Span4Mux_v I__18974 (
            .O(N__76917),
            .I(N__76887));
    CascadeMux I__18973 (
            .O(N__76916),
            .I(N__76884));
    Span4Mux_v I__18972 (
            .O(N__76913),
            .I(N__76880));
    InMux I__18971 (
            .O(N__76912),
            .I(N__76877));
    LocalMux I__18970 (
            .O(N__76909),
            .I(N__76874));
    LocalMux I__18969 (
            .O(N__76906),
            .I(N__76865));
    Span4Mux_h I__18968 (
            .O(N__76903),
            .I(N__76865));
    Span4Mux_v I__18967 (
            .O(N__76900),
            .I(N__76865));
    Span4Mux_v I__18966 (
            .O(N__76895),
            .I(N__76865));
    Span4Mux_h I__18965 (
            .O(N__76892),
            .I(N__76860));
    Span4Mux_v I__18964 (
            .O(N__76887),
            .I(N__76860));
    InMux I__18963 (
            .O(N__76884),
            .I(N__76855));
    InMux I__18962 (
            .O(N__76883),
            .I(N__76855));
    Span4Mux_v I__18961 (
            .O(N__76880),
            .I(N__76852));
    LocalMux I__18960 (
            .O(N__76877),
            .I(N__76845));
    Span4Mux_v I__18959 (
            .O(N__76874),
            .I(N__76845));
    Span4Mux_h I__18958 (
            .O(N__76865),
            .I(N__76845));
    Span4Mux_h I__18957 (
            .O(N__76860),
            .I(N__76842));
    LocalMux I__18956 (
            .O(N__76855),
            .I(rx_data_3));
    Odrv4 I__18955 (
            .O(N__76852),
            .I(rx_data_3));
    Odrv4 I__18954 (
            .O(N__76845),
            .I(rx_data_3));
    Odrv4 I__18953 (
            .O(N__76842),
            .I(rx_data_3));
    InMux I__18952 (
            .O(N__76833),
            .I(N__76829));
    InMux I__18951 (
            .O(N__76832),
            .I(N__76825));
    LocalMux I__18950 (
            .O(N__76829),
            .I(N__76822));
    InMux I__18949 (
            .O(N__76828),
            .I(N__76819));
    LocalMux I__18948 (
            .O(N__76825),
            .I(N__76816));
    Span4Mux_v I__18947 (
            .O(N__76822),
            .I(N__76810));
    LocalMux I__18946 (
            .O(N__76819),
            .I(N__76810));
    Span4Mux_h I__18945 (
            .O(N__76816),
            .I(N__76807));
    CascadeMux I__18944 (
            .O(N__76815),
            .I(N__76804));
    Span4Mux_h I__18943 (
            .O(N__76810),
            .I(N__76801));
    Span4Mux_h I__18942 (
            .O(N__76807),
            .I(N__76798));
    InMux I__18941 (
            .O(N__76804),
            .I(N__76794));
    Span4Mux_h I__18940 (
            .O(N__76801),
            .I(N__76791));
    Span4Mux_v I__18939 (
            .O(N__76798),
            .I(N__76788));
    InMux I__18938 (
            .O(N__76797),
            .I(N__76785));
    LocalMux I__18937 (
            .O(N__76794),
            .I(\c0.data_in_frame_23_3 ));
    Odrv4 I__18936 (
            .O(N__76791),
            .I(\c0.data_in_frame_23_3 ));
    Odrv4 I__18935 (
            .O(N__76788),
            .I(\c0.data_in_frame_23_3 ));
    LocalMux I__18934 (
            .O(N__76785),
            .I(\c0.data_in_frame_23_3 ));
    InMux I__18933 (
            .O(N__76776),
            .I(N__76773));
    LocalMux I__18932 (
            .O(N__76773),
            .I(N__76770));
    Odrv4 I__18931 (
            .O(N__76770),
            .I(\c0.n25484 ));
    InMux I__18930 (
            .O(N__76767),
            .I(N__76764));
    LocalMux I__18929 (
            .O(N__76764),
            .I(N__76761));
    Odrv4 I__18928 (
            .O(N__76761),
            .I(\c0.n62 ));
    CascadeMux I__18927 (
            .O(N__76758),
            .I(N__76755));
    InMux I__18926 (
            .O(N__76755),
            .I(N__76752));
    LocalMux I__18925 (
            .O(N__76752),
            .I(\c0.n21_adj_4481 ));
    InMux I__18924 (
            .O(N__76749),
            .I(N__76746));
    LocalMux I__18923 (
            .O(N__76746),
            .I(N__76743));
    Span4Mux_v I__18922 (
            .O(N__76743),
            .I(N__76738));
    InMux I__18921 (
            .O(N__76742),
            .I(N__76735));
    InMux I__18920 (
            .O(N__76741),
            .I(N__76732));
    Span4Mux_h I__18919 (
            .O(N__76738),
            .I(N__76727));
    LocalMux I__18918 (
            .O(N__76735),
            .I(N__76727));
    LocalMux I__18917 (
            .O(N__76732),
            .I(N__76723));
    Span4Mux_h I__18916 (
            .O(N__76727),
            .I(N__76720));
    InMux I__18915 (
            .O(N__76726),
            .I(N__76717));
    Odrv12 I__18914 (
            .O(N__76723),
            .I(\c0.n6_adj_4462 ));
    Odrv4 I__18913 (
            .O(N__76720),
            .I(\c0.n6_adj_4462 ));
    LocalMux I__18912 (
            .O(N__76717),
            .I(\c0.n6_adj_4462 ));
    InMux I__18911 (
            .O(N__76710),
            .I(N__76707));
    LocalMux I__18910 (
            .O(N__76707),
            .I(N__76704));
    Span4Mux_h I__18909 (
            .O(N__76704),
            .I(N__76701));
    Span4Mux_h I__18908 (
            .O(N__76701),
            .I(N__76698));
    Odrv4 I__18907 (
            .O(N__76698),
            .I(\c0.n30_adj_4482 ));
    InMux I__18906 (
            .O(N__76695),
            .I(N__76688));
    InMux I__18905 (
            .O(N__76694),
            .I(N__76688));
    InMux I__18904 (
            .O(N__76693),
            .I(N__76684));
    LocalMux I__18903 (
            .O(N__76688),
            .I(N__76679));
    InMux I__18902 (
            .O(N__76687),
            .I(N__76676));
    LocalMux I__18901 (
            .O(N__76684),
            .I(N__76671));
    InMux I__18900 (
            .O(N__76683),
            .I(N__76668));
    InMux I__18899 (
            .O(N__76682),
            .I(N__76665));
    Span4Mux_v I__18898 (
            .O(N__76679),
            .I(N__76660));
    LocalMux I__18897 (
            .O(N__76676),
            .I(N__76660));
    InMux I__18896 (
            .O(N__76675),
            .I(N__76657));
    InMux I__18895 (
            .O(N__76674),
            .I(N__76649));
    Span4Mux_v I__18894 (
            .O(N__76671),
            .I(N__76644));
    LocalMux I__18893 (
            .O(N__76668),
            .I(N__76644));
    LocalMux I__18892 (
            .O(N__76665),
            .I(N__76641));
    Span4Mux_v I__18891 (
            .O(N__76660),
            .I(N__76636));
    LocalMux I__18890 (
            .O(N__76657),
            .I(N__76636));
    InMux I__18889 (
            .O(N__76656),
            .I(N__76631));
    InMux I__18888 (
            .O(N__76655),
            .I(N__76631));
    InMux I__18887 (
            .O(N__76654),
            .I(N__76626));
    InMux I__18886 (
            .O(N__76653),
            .I(N__76617));
    InMux I__18885 (
            .O(N__76652),
            .I(N__76617));
    LocalMux I__18884 (
            .O(N__76649),
            .I(N__76614));
    Span4Mux_v I__18883 (
            .O(N__76644),
            .I(N__76607));
    Span4Mux_v I__18882 (
            .O(N__76641),
            .I(N__76600));
    Span4Mux_v I__18881 (
            .O(N__76636),
            .I(N__76600));
    LocalMux I__18880 (
            .O(N__76631),
            .I(N__76600));
    CascadeMux I__18879 (
            .O(N__76630),
            .I(N__76596));
    InMux I__18878 (
            .O(N__76629),
            .I(N__76592));
    LocalMux I__18877 (
            .O(N__76626),
            .I(N__76589));
    InMux I__18876 (
            .O(N__76625),
            .I(N__76586));
    InMux I__18875 (
            .O(N__76624),
            .I(N__76583));
    InMux I__18874 (
            .O(N__76623),
            .I(N__76579));
    InMux I__18873 (
            .O(N__76622),
            .I(N__76576));
    LocalMux I__18872 (
            .O(N__76617),
            .I(N__76573));
    Span4Mux_h I__18871 (
            .O(N__76614),
            .I(N__76570));
    InMux I__18870 (
            .O(N__76613),
            .I(N__76567));
    InMux I__18869 (
            .O(N__76612),
            .I(N__76564));
    InMux I__18868 (
            .O(N__76611),
            .I(N__76559));
    InMux I__18867 (
            .O(N__76610),
            .I(N__76559));
    Span4Mux_h I__18866 (
            .O(N__76607),
            .I(N__76554));
    Span4Mux_h I__18865 (
            .O(N__76600),
            .I(N__76554));
    CascadeMux I__18864 (
            .O(N__76599),
            .I(N__76551));
    InMux I__18863 (
            .O(N__76596),
            .I(N__76545));
    InMux I__18862 (
            .O(N__76595),
            .I(N__76542));
    LocalMux I__18861 (
            .O(N__76592),
            .I(N__76539));
    Span4Mux_v I__18860 (
            .O(N__76589),
            .I(N__76536));
    LocalMux I__18859 (
            .O(N__76586),
            .I(N__76531));
    LocalMux I__18858 (
            .O(N__76583),
            .I(N__76531));
    InMux I__18857 (
            .O(N__76582),
            .I(N__76526));
    LocalMux I__18856 (
            .O(N__76579),
            .I(N__76520));
    LocalMux I__18855 (
            .O(N__76576),
            .I(N__76520));
    Span4Mux_v I__18854 (
            .O(N__76573),
            .I(N__76513));
    Span4Mux_h I__18853 (
            .O(N__76570),
            .I(N__76513));
    LocalMux I__18852 (
            .O(N__76567),
            .I(N__76513));
    LocalMux I__18851 (
            .O(N__76564),
            .I(N__76510));
    LocalMux I__18850 (
            .O(N__76559),
            .I(N__76505));
    Span4Mux_v I__18849 (
            .O(N__76554),
            .I(N__76505));
    InMux I__18848 (
            .O(N__76551),
            .I(N__76502));
    InMux I__18847 (
            .O(N__76550),
            .I(N__76499));
    InMux I__18846 (
            .O(N__76549),
            .I(N__76496));
    InMux I__18845 (
            .O(N__76548),
            .I(N__76493));
    LocalMux I__18844 (
            .O(N__76545),
            .I(N__76484));
    LocalMux I__18843 (
            .O(N__76542),
            .I(N__76484));
    Span4Mux_h I__18842 (
            .O(N__76539),
            .I(N__76484));
    Span4Mux_v I__18841 (
            .O(N__76536),
            .I(N__76484));
    Span4Mux_v I__18840 (
            .O(N__76531),
            .I(N__76481));
    InMux I__18839 (
            .O(N__76530),
            .I(N__76478));
    InMux I__18838 (
            .O(N__76529),
            .I(N__76475));
    LocalMux I__18837 (
            .O(N__76526),
            .I(N__76472));
    InMux I__18836 (
            .O(N__76525),
            .I(N__76469));
    Span4Mux_v I__18835 (
            .O(N__76520),
            .I(N__76464));
    Span4Mux_v I__18834 (
            .O(N__76513),
            .I(N__76464));
    Span4Mux_h I__18833 (
            .O(N__76510),
            .I(N__76459));
    Span4Mux_v I__18832 (
            .O(N__76505),
            .I(N__76459));
    LocalMux I__18831 (
            .O(N__76502),
            .I(N__76456));
    LocalMux I__18830 (
            .O(N__76499),
            .I(N__76449));
    LocalMux I__18829 (
            .O(N__76496),
            .I(N__76449));
    LocalMux I__18828 (
            .O(N__76493),
            .I(N__76449));
    Span4Mux_h I__18827 (
            .O(N__76484),
            .I(N__76446));
    Sp12to4 I__18826 (
            .O(N__76481),
            .I(N__76443));
    LocalMux I__18825 (
            .O(N__76478),
            .I(N__76434));
    LocalMux I__18824 (
            .O(N__76475),
            .I(N__76434));
    Span12Mux_v I__18823 (
            .O(N__76472),
            .I(N__76434));
    LocalMux I__18822 (
            .O(N__76469),
            .I(N__76434));
    Span4Mux_h I__18821 (
            .O(N__76464),
            .I(N__76429));
    Span4Mux_v I__18820 (
            .O(N__76459),
            .I(N__76429));
    Span4Mux_v I__18819 (
            .O(N__76456),
            .I(N__76426));
    Span4Mux_v I__18818 (
            .O(N__76449),
            .I(N__76423));
    Span4Mux_h I__18817 (
            .O(N__76446),
            .I(N__76420));
    Span12Mux_h I__18816 (
            .O(N__76443),
            .I(N__76417));
    Span12Mux_v I__18815 (
            .O(N__76434),
            .I(N__76414));
    Span4Mux_v I__18814 (
            .O(N__76429),
            .I(N__76411));
    Odrv4 I__18813 (
            .O(N__76426),
            .I(\c0.n9_adj_4273 ));
    Odrv4 I__18812 (
            .O(N__76423),
            .I(\c0.n9_adj_4273 ));
    Odrv4 I__18811 (
            .O(N__76420),
            .I(\c0.n9_adj_4273 ));
    Odrv12 I__18810 (
            .O(N__76417),
            .I(\c0.n9_adj_4273 ));
    Odrv12 I__18809 (
            .O(N__76414),
            .I(\c0.n9_adj_4273 ));
    Odrv4 I__18808 (
            .O(N__76411),
            .I(\c0.n9_adj_4273 ));
    CascadeMux I__18807 (
            .O(N__76398),
            .I(N__76395));
    InMux I__18806 (
            .O(N__76395),
            .I(N__76390));
    InMux I__18805 (
            .O(N__76394),
            .I(N__76386));
    InMux I__18804 (
            .O(N__76393),
            .I(N__76379));
    LocalMux I__18803 (
            .O(N__76390),
            .I(N__76375));
    InMux I__18802 (
            .O(N__76389),
            .I(N__76372));
    LocalMux I__18801 (
            .O(N__76386),
            .I(N__76369));
    InMux I__18800 (
            .O(N__76385),
            .I(N__76366));
    InMux I__18799 (
            .O(N__76384),
            .I(N__76362));
    CascadeMux I__18798 (
            .O(N__76383),
            .I(N__76359));
    CascadeMux I__18797 (
            .O(N__76382),
            .I(N__76356));
    LocalMux I__18796 (
            .O(N__76379),
            .I(N__76351));
    InMux I__18795 (
            .O(N__76378),
            .I(N__76348));
    Span4Mux_h I__18794 (
            .O(N__76375),
            .I(N__76343));
    LocalMux I__18793 (
            .O(N__76372),
            .I(N__76343));
    Span4Mux_v I__18792 (
            .O(N__76369),
            .I(N__76338));
    LocalMux I__18791 (
            .O(N__76366),
            .I(N__76338));
    CascadeMux I__18790 (
            .O(N__76365),
            .I(N__76335));
    LocalMux I__18789 (
            .O(N__76362),
            .I(N__76332));
    InMux I__18788 (
            .O(N__76359),
            .I(N__76329));
    InMux I__18787 (
            .O(N__76356),
            .I(N__76326));
    InMux I__18786 (
            .O(N__76355),
            .I(N__76321));
    InMux I__18785 (
            .O(N__76354),
            .I(N__76318));
    Span4Mux_v I__18784 (
            .O(N__76351),
            .I(N__76310));
    LocalMux I__18783 (
            .O(N__76348),
            .I(N__76310));
    Span4Mux_v I__18782 (
            .O(N__76343),
            .I(N__76305));
    Span4Mux_h I__18781 (
            .O(N__76338),
            .I(N__76305));
    InMux I__18780 (
            .O(N__76335),
            .I(N__76302));
    Span4Mux_h I__18779 (
            .O(N__76332),
            .I(N__76295));
    LocalMux I__18778 (
            .O(N__76329),
            .I(N__76295));
    LocalMux I__18777 (
            .O(N__76326),
            .I(N__76295));
    CascadeMux I__18776 (
            .O(N__76325),
            .I(N__76290));
    InMux I__18775 (
            .O(N__76324),
            .I(N__76286));
    LocalMux I__18774 (
            .O(N__76321),
            .I(N__76282));
    LocalMux I__18773 (
            .O(N__76318),
            .I(N__76279));
    InMux I__18772 (
            .O(N__76317),
            .I(N__76276));
    InMux I__18771 (
            .O(N__76316),
            .I(N__76271));
    InMux I__18770 (
            .O(N__76315),
            .I(N__76268));
    Span4Mux_v I__18769 (
            .O(N__76310),
            .I(N__76265));
    Span4Mux_h I__18768 (
            .O(N__76305),
            .I(N__76260));
    LocalMux I__18767 (
            .O(N__76302),
            .I(N__76260));
    Span4Mux_v I__18766 (
            .O(N__76295),
            .I(N__76257));
    CascadeMux I__18765 (
            .O(N__76294),
            .I(N__76254));
    InMux I__18764 (
            .O(N__76293),
            .I(N__76251));
    InMux I__18763 (
            .O(N__76290),
            .I(N__76248));
    InMux I__18762 (
            .O(N__76289),
            .I(N__76245));
    LocalMux I__18761 (
            .O(N__76286),
            .I(N__76242));
    InMux I__18760 (
            .O(N__76285),
            .I(N__76239));
    Span4Mux_v I__18759 (
            .O(N__76282),
            .I(N__76232));
    Span4Mux_h I__18758 (
            .O(N__76279),
            .I(N__76232));
    LocalMux I__18757 (
            .O(N__76276),
            .I(N__76232));
    CascadeMux I__18756 (
            .O(N__76275),
            .I(N__76229));
    InMux I__18755 (
            .O(N__76274),
            .I(N__76224));
    LocalMux I__18754 (
            .O(N__76271),
            .I(N__76221));
    LocalMux I__18753 (
            .O(N__76268),
            .I(N__76218));
    Span4Mux_h I__18752 (
            .O(N__76265),
            .I(N__76215));
    Span4Mux_v I__18751 (
            .O(N__76260),
            .I(N__76212));
    Span4Mux_h I__18750 (
            .O(N__76257),
            .I(N__76209));
    InMux I__18749 (
            .O(N__76254),
            .I(N__76206));
    LocalMux I__18748 (
            .O(N__76251),
            .I(N__76199));
    LocalMux I__18747 (
            .O(N__76248),
            .I(N__76199));
    LocalMux I__18746 (
            .O(N__76245),
            .I(N__76199));
    Span4Mux_v I__18745 (
            .O(N__76242),
            .I(N__76194));
    LocalMux I__18744 (
            .O(N__76239),
            .I(N__76194));
    Span4Mux_v I__18743 (
            .O(N__76232),
            .I(N__76191));
    InMux I__18742 (
            .O(N__76229),
            .I(N__76188));
    InMux I__18741 (
            .O(N__76228),
            .I(N__76183));
    InMux I__18740 (
            .O(N__76227),
            .I(N__76183));
    LocalMux I__18739 (
            .O(N__76224),
            .I(N__76180));
    Span4Mux_v I__18738 (
            .O(N__76221),
            .I(N__76175));
    Span4Mux_h I__18737 (
            .O(N__76218),
            .I(N__76175));
    Sp12to4 I__18736 (
            .O(N__76215),
            .I(N__76172));
    Sp12to4 I__18735 (
            .O(N__76212),
            .I(N__76167));
    Sp12to4 I__18734 (
            .O(N__76209),
            .I(N__76167));
    LocalMux I__18733 (
            .O(N__76206),
            .I(N__76164));
    Span4Mux_v I__18732 (
            .O(N__76199),
            .I(N__76161));
    Span4Mux_h I__18731 (
            .O(N__76194),
            .I(N__76158));
    Span4Mux_h I__18730 (
            .O(N__76191),
            .I(N__76155));
    LocalMux I__18729 (
            .O(N__76188),
            .I(N__76135));
    LocalMux I__18728 (
            .O(N__76183),
            .I(N__76135));
    Span12Mux_h I__18727 (
            .O(N__76180),
            .I(N__76135));
    Sp12to4 I__18726 (
            .O(N__76175),
            .I(N__76135));
    Span12Mux_h I__18725 (
            .O(N__76172),
            .I(N__76135));
    Span12Mux_h I__18724 (
            .O(N__76167),
            .I(N__76135));
    Span4Mux_v I__18723 (
            .O(N__76164),
            .I(N__76130));
    Span4Mux_v I__18722 (
            .O(N__76161),
            .I(N__76130));
    Span4Mux_v I__18721 (
            .O(N__76158),
            .I(N__76125));
    Span4Mux_v I__18720 (
            .O(N__76155),
            .I(N__76125));
    InMux I__18719 (
            .O(N__76154),
            .I(N__76122));
    InMux I__18718 (
            .O(N__76153),
            .I(N__76117));
    InMux I__18717 (
            .O(N__76152),
            .I(N__76117));
    InMux I__18716 (
            .O(N__76151),
            .I(N__76112));
    InMux I__18715 (
            .O(N__76150),
            .I(N__76112));
    InMux I__18714 (
            .O(N__76149),
            .I(N__76107));
    InMux I__18713 (
            .O(N__76148),
            .I(N__76107));
    Span12Mux_v I__18712 (
            .O(N__76135),
            .I(N__76104));
    Span4Mux_h I__18711 (
            .O(N__76130),
            .I(N__76099));
    Span4Mux_v I__18710 (
            .O(N__76125),
            .I(N__76099));
    LocalMux I__18709 (
            .O(N__76122),
            .I(rx_data_7));
    LocalMux I__18708 (
            .O(N__76117),
            .I(rx_data_7));
    LocalMux I__18707 (
            .O(N__76112),
            .I(rx_data_7));
    LocalMux I__18706 (
            .O(N__76107),
            .I(rx_data_7));
    Odrv12 I__18705 (
            .O(N__76104),
            .I(rx_data_7));
    Odrv4 I__18704 (
            .O(N__76099),
            .I(rx_data_7));
    InMux I__18703 (
            .O(N__76086),
            .I(N__76083));
    LocalMux I__18702 (
            .O(N__76083),
            .I(N__76079));
    InMux I__18701 (
            .O(N__76082),
            .I(N__76076));
    Span4Mux_h I__18700 (
            .O(N__76079),
            .I(N__76071));
    LocalMux I__18699 (
            .O(N__76076),
            .I(N__76071));
    Span4Mux_h I__18698 (
            .O(N__76071),
            .I(N__76067));
    CascadeMux I__18697 (
            .O(N__76070),
            .I(N__76064));
    Sp12to4 I__18696 (
            .O(N__76067),
            .I(N__76061));
    InMux I__18695 (
            .O(N__76064),
            .I(N__76058));
    Odrv12 I__18694 (
            .O(N__76061),
            .I(\c0.n23598 ));
    LocalMux I__18693 (
            .O(N__76058),
            .I(\c0.n23598 ));
    InMux I__18692 (
            .O(N__76053),
            .I(N__76049));
    InMux I__18691 (
            .O(N__76052),
            .I(N__76044));
    LocalMux I__18690 (
            .O(N__76049),
            .I(N__76041));
    CascadeMux I__18689 (
            .O(N__76048),
            .I(N__76038));
    CascadeMux I__18688 (
            .O(N__76047),
            .I(N__76033));
    LocalMux I__18687 (
            .O(N__76044),
            .I(N__76030));
    Span4Mux_v I__18686 (
            .O(N__76041),
            .I(N__76027));
    InMux I__18685 (
            .O(N__76038),
            .I(N__76022));
    InMux I__18684 (
            .O(N__76037),
            .I(N__76022));
    InMux I__18683 (
            .O(N__76036),
            .I(N__76019));
    InMux I__18682 (
            .O(N__76033),
            .I(N__76016));
    Span4Mux_h I__18681 (
            .O(N__76030),
            .I(N__76013));
    Span4Mux_h I__18680 (
            .O(N__76027),
            .I(N__76008));
    LocalMux I__18679 (
            .O(N__76022),
            .I(N__76008));
    LocalMux I__18678 (
            .O(N__76019),
            .I(N__76005));
    LocalMux I__18677 (
            .O(N__76016),
            .I(\c0.data_in_frame_8_4 ));
    Odrv4 I__18676 (
            .O(N__76013),
            .I(\c0.data_in_frame_8_4 ));
    Odrv4 I__18675 (
            .O(N__76008),
            .I(\c0.data_in_frame_8_4 ));
    Odrv12 I__18674 (
            .O(N__76005),
            .I(\c0.data_in_frame_8_4 ));
    CascadeMux I__18673 (
            .O(N__75996),
            .I(N__75993));
    InMux I__18672 (
            .O(N__75993),
            .I(N__75990));
    LocalMux I__18671 (
            .O(N__75990),
            .I(N__75986));
    CascadeMux I__18670 (
            .O(N__75989),
            .I(N__75983));
    Span12Mux_s10_h I__18669 (
            .O(N__75986),
            .I(N__75980));
    InMux I__18668 (
            .O(N__75983),
            .I(N__75977));
    Span12Mux_v I__18667 (
            .O(N__75980),
            .I(N__75974));
    LocalMux I__18666 (
            .O(N__75977),
            .I(\c0.data_in_frame_26_6 ));
    Odrv12 I__18665 (
            .O(N__75974),
            .I(\c0.data_in_frame_26_6 ));
    InMux I__18664 (
            .O(N__75969),
            .I(N__75966));
    LocalMux I__18663 (
            .O(N__75966),
            .I(N__75963));
    Span12Mux_h I__18662 (
            .O(N__75963),
            .I(N__75959));
    InMux I__18661 (
            .O(N__75962),
            .I(N__75956));
    Odrv12 I__18660 (
            .O(N__75959),
            .I(\c0.n22769 ));
    LocalMux I__18659 (
            .O(N__75956),
            .I(\c0.n22769 ));
    InMux I__18658 (
            .O(N__75951),
            .I(N__75948));
    LocalMux I__18657 (
            .O(N__75948),
            .I(N__75943));
    InMux I__18656 (
            .O(N__75947),
            .I(N__75940));
    InMux I__18655 (
            .O(N__75946),
            .I(N__75935));
    Span4Mux_h I__18654 (
            .O(N__75943),
            .I(N__75932));
    LocalMux I__18653 (
            .O(N__75940),
            .I(N__75929));
    InMux I__18652 (
            .O(N__75939),
            .I(N__75926));
    CascadeMux I__18651 (
            .O(N__75938),
            .I(N__75923));
    LocalMux I__18650 (
            .O(N__75935),
            .I(N__75920));
    Span4Mux_v I__18649 (
            .O(N__75932),
            .I(N__75913));
    Span4Mux_h I__18648 (
            .O(N__75929),
            .I(N__75913));
    LocalMux I__18647 (
            .O(N__75926),
            .I(N__75913));
    InMux I__18646 (
            .O(N__75923),
            .I(N__75910));
    Span4Mux_h I__18645 (
            .O(N__75920),
            .I(N__75906));
    Span4Mux_v I__18644 (
            .O(N__75913),
            .I(N__75903));
    LocalMux I__18643 (
            .O(N__75910),
            .I(N__75900));
    InMux I__18642 (
            .O(N__75909),
            .I(N__75897));
    Span4Mux_h I__18641 (
            .O(N__75906),
            .I(N__75894));
    Span4Mux_h I__18640 (
            .O(N__75903),
            .I(N__75891));
    Span12Mux_v I__18639 (
            .O(N__75900),
            .I(N__75888));
    LocalMux I__18638 (
            .O(N__75897),
            .I(N__75883));
    Span4Mux_v I__18637 (
            .O(N__75894),
            .I(N__75883));
    Span4Mux_h I__18636 (
            .O(N__75891),
            .I(N__75880));
    Odrv12 I__18635 (
            .O(N__75888),
            .I(data_in_frame_21_5));
    Odrv4 I__18634 (
            .O(N__75883),
            .I(data_in_frame_21_5));
    Odrv4 I__18633 (
            .O(N__75880),
            .I(data_in_frame_21_5));
    InMux I__18632 (
            .O(N__75873),
            .I(N__75870));
    LocalMux I__18631 (
            .O(N__75870),
            .I(N__75867));
    Span4Mux_v I__18630 (
            .O(N__75867),
            .I(N__75864));
    Span4Mux_h I__18629 (
            .O(N__75864),
            .I(N__75861));
    Odrv4 I__18628 (
            .O(N__75861),
            .I(\c0.n22698 ));
    CascadeMux I__18627 (
            .O(N__75858),
            .I(N__75854));
    CascadeMux I__18626 (
            .O(N__75857),
            .I(N__75851));
    InMux I__18625 (
            .O(N__75854),
            .I(N__75848));
    InMux I__18624 (
            .O(N__75851),
            .I(N__75844));
    LocalMux I__18623 (
            .O(N__75848),
            .I(N__75841));
    InMux I__18622 (
            .O(N__75847),
            .I(N__75838));
    LocalMux I__18621 (
            .O(N__75844),
            .I(N__75831));
    Span4Mux_v I__18620 (
            .O(N__75841),
            .I(N__75831));
    LocalMux I__18619 (
            .O(N__75838),
            .I(N__75831));
    Span4Mux_h I__18618 (
            .O(N__75831),
            .I(N__75827));
    CascadeMux I__18617 (
            .O(N__75830),
            .I(N__75824));
    Span4Mux_h I__18616 (
            .O(N__75827),
            .I(N__75820));
    InMux I__18615 (
            .O(N__75824),
            .I(N__75815));
    InMux I__18614 (
            .O(N__75823),
            .I(N__75815));
    Odrv4 I__18613 (
            .O(N__75820),
            .I(\c0.data_in_frame_23_6 ));
    LocalMux I__18612 (
            .O(N__75815),
            .I(\c0.data_in_frame_23_6 ));
    InMux I__18611 (
            .O(N__75810),
            .I(N__75807));
    LocalMux I__18610 (
            .O(N__75807),
            .I(N__75804));
    Span4Mux_h I__18609 (
            .O(N__75804),
            .I(N__75801));
    Span4Mux_h I__18608 (
            .O(N__75801),
            .I(N__75798));
    Odrv4 I__18607 (
            .O(N__75798),
            .I(\c0.n4_adj_4464 ));
    InMux I__18606 (
            .O(N__75795),
            .I(N__75792));
    LocalMux I__18605 (
            .O(N__75792),
            .I(N__75789));
    Odrv12 I__18604 (
            .O(N__75789),
            .I(\c0.n14_adj_4465 ));
    InMux I__18603 (
            .O(N__75786),
            .I(N__75779));
    InMux I__18602 (
            .O(N__75785),
            .I(N__75779));
    InMux I__18601 (
            .O(N__75784),
            .I(N__75775));
    LocalMux I__18600 (
            .O(N__75779),
            .I(N__75772));
    InMux I__18599 (
            .O(N__75778),
            .I(N__75769));
    LocalMux I__18598 (
            .O(N__75775),
            .I(N__75766));
    Span4Mux_h I__18597 (
            .O(N__75772),
            .I(N__75762));
    LocalMux I__18596 (
            .O(N__75769),
            .I(N__75757));
    Span4Mux_h I__18595 (
            .O(N__75766),
            .I(N__75757));
    CascadeMux I__18594 (
            .O(N__75765),
            .I(N__75754));
    Sp12to4 I__18593 (
            .O(N__75762),
            .I(N__75751));
    Span4Mux_v I__18592 (
            .O(N__75757),
            .I(N__75748));
    InMux I__18591 (
            .O(N__75754),
            .I(N__75745));
    Span12Mux_v I__18590 (
            .O(N__75751),
            .I(N__75742));
    Span4Mux_v I__18589 (
            .O(N__75748),
            .I(N__75739));
    LocalMux I__18588 (
            .O(N__75745),
            .I(\c0.data_in_frame_20_3 ));
    Odrv12 I__18587 (
            .O(N__75742),
            .I(\c0.data_in_frame_20_3 ));
    Odrv4 I__18586 (
            .O(N__75739),
            .I(\c0.data_in_frame_20_3 ));
    InMux I__18585 (
            .O(N__75732),
            .I(N__75726));
    InMux I__18584 (
            .O(N__75731),
            .I(N__75719));
    InMux I__18583 (
            .O(N__75730),
            .I(N__75719));
    InMux I__18582 (
            .O(N__75729),
            .I(N__75719));
    LocalMux I__18581 (
            .O(N__75726),
            .I(N__75716));
    LocalMux I__18580 (
            .O(N__75719),
            .I(N__75713));
    Odrv12 I__18579 (
            .O(N__75716),
            .I(\c0.n21412 ));
    Odrv4 I__18578 (
            .O(N__75713),
            .I(\c0.n21412 ));
    InMux I__18577 (
            .O(N__75708),
            .I(N__75705));
    LocalMux I__18576 (
            .O(N__75705),
            .I(\c0.n4_adj_4369 ));
    CascadeMux I__18575 (
            .O(N__75702),
            .I(N__75697));
    CascadeMux I__18574 (
            .O(N__75701),
            .I(N__75694));
    CascadeMux I__18573 (
            .O(N__75700),
            .I(N__75691));
    InMux I__18572 (
            .O(N__75697),
            .I(N__75688));
    InMux I__18571 (
            .O(N__75694),
            .I(N__75685));
    InMux I__18570 (
            .O(N__75691),
            .I(N__75682));
    LocalMux I__18569 (
            .O(N__75688),
            .I(N__75679));
    LocalMux I__18568 (
            .O(N__75685),
            .I(N__75675));
    LocalMux I__18567 (
            .O(N__75682),
            .I(N__75672));
    Span4Mux_h I__18566 (
            .O(N__75679),
            .I(N__75669));
    CascadeMux I__18565 (
            .O(N__75678),
            .I(N__75666));
    Span4Mux_h I__18564 (
            .O(N__75675),
            .I(N__75663));
    Span4Mux_h I__18563 (
            .O(N__75672),
            .I(N__75660));
    Span4Mux_h I__18562 (
            .O(N__75669),
            .I(N__75657));
    InMux I__18561 (
            .O(N__75666),
            .I(N__75654));
    Span4Mux_h I__18560 (
            .O(N__75663),
            .I(N__75649));
    Span4Mux_h I__18559 (
            .O(N__75660),
            .I(N__75649));
    Span4Mux_v I__18558 (
            .O(N__75657),
            .I(N__75646));
    LocalMux I__18557 (
            .O(N__75654),
            .I(N__75641));
    Span4Mux_v I__18556 (
            .O(N__75649),
            .I(N__75641));
    Odrv4 I__18555 (
            .O(N__75646),
            .I(\c0.data_in_frame_27_0 ));
    Odrv4 I__18554 (
            .O(N__75641),
            .I(\c0.data_in_frame_27_0 ));
    CascadeMux I__18553 (
            .O(N__75636),
            .I(N__75633));
    InMux I__18552 (
            .O(N__75633),
            .I(N__75630));
    LocalMux I__18551 (
            .O(N__75630),
            .I(N__75627));
    Span4Mux_h I__18550 (
            .O(N__75627),
            .I(N__75624));
    Odrv4 I__18549 (
            .O(N__75624),
            .I(\c0.n73 ));
    InMux I__18548 (
            .O(N__75621),
            .I(N__75615));
    InMux I__18547 (
            .O(N__75620),
            .I(N__75615));
    LocalMux I__18546 (
            .O(N__75615),
            .I(N__75608));
    InMux I__18545 (
            .O(N__75614),
            .I(N__75605));
    InMux I__18544 (
            .O(N__75613),
            .I(N__75600));
    InMux I__18543 (
            .O(N__75612),
            .I(N__75600));
    InMux I__18542 (
            .O(N__75611),
            .I(N__75597));
    Span4Mux_v I__18541 (
            .O(N__75608),
            .I(N__75590));
    LocalMux I__18540 (
            .O(N__75605),
            .I(N__75590));
    LocalMux I__18539 (
            .O(N__75600),
            .I(N__75590));
    LocalMux I__18538 (
            .O(N__75597),
            .I(N__75587));
    Span4Mux_h I__18537 (
            .O(N__75590),
            .I(N__75584));
    Span4Mux_v I__18536 (
            .O(N__75587),
            .I(N__75579));
    Span4Mux_h I__18535 (
            .O(N__75584),
            .I(N__75579));
    Odrv4 I__18534 (
            .O(N__75579),
            .I(\c0.n20409 ));
    CascadeMux I__18533 (
            .O(N__75576),
            .I(N__75573));
    InMux I__18532 (
            .O(N__75573),
            .I(N__75570));
    LocalMux I__18531 (
            .O(N__75570),
            .I(N__75567));
    Span4Mux_h I__18530 (
            .O(N__75567),
            .I(N__75563));
    InMux I__18529 (
            .O(N__75566),
            .I(N__75559));
    Sp12to4 I__18528 (
            .O(N__75563),
            .I(N__75555));
    CascadeMux I__18527 (
            .O(N__75562),
            .I(N__75550));
    LocalMux I__18526 (
            .O(N__75559),
            .I(N__75545));
    InMux I__18525 (
            .O(N__75558),
            .I(N__75542));
    Span12Mux_v I__18524 (
            .O(N__75555),
            .I(N__75539));
    InMux I__18523 (
            .O(N__75554),
            .I(N__75536));
    InMux I__18522 (
            .O(N__75553),
            .I(N__75533));
    InMux I__18521 (
            .O(N__75550),
            .I(N__75528));
    InMux I__18520 (
            .O(N__75549),
            .I(N__75528));
    InMux I__18519 (
            .O(N__75548),
            .I(N__75525));
    Span4Mux_v I__18518 (
            .O(N__75545),
            .I(N__75522));
    LocalMux I__18517 (
            .O(N__75542),
            .I(data_in_frame_22_4));
    Odrv12 I__18516 (
            .O(N__75539),
            .I(data_in_frame_22_4));
    LocalMux I__18515 (
            .O(N__75536),
            .I(data_in_frame_22_4));
    LocalMux I__18514 (
            .O(N__75533),
            .I(data_in_frame_22_4));
    LocalMux I__18513 (
            .O(N__75528),
            .I(data_in_frame_22_4));
    LocalMux I__18512 (
            .O(N__75525),
            .I(data_in_frame_22_4));
    Odrv4 I__18511 (
            .O(N__75522),
            .I(data_in_frame_22_4));
    InMux I__18510 (
            .O(N__75507),
            .I(N__75501));
    InMux I__18509 (
            .O(N__75506),
            .I(N__75501));
    LocalMux I__18508 (
            .O(N__75501),
            .I(N__75495));
    InMux I__18507 (
            .O(N__75500),
            .I(N__75489));
    InMux I__18506 (
            .O(N__75499),
            .I(N__75484));
    InMux I__18505 (
            .O(N__75498),
            .I(N__75484));
    Span4Mux_h I__18504 (
            .O(N__75495),
            .I(N__75481));
    InMux I__18503 (
            .O(N__75494),
            .I(N__75476));
    InMux I__18502 (
            .O(N__75493),
            .I(N__75476));
    InMux I__18501 (
            .O(N__75492),
            .I(N__75473));
    LocalMux I__18500 (
            .O(N__75489),
            .I(N__75470));
    LocalMux I__18499 (
            .O(N__75484),
            .I(N__75467));
    Span4Mux_v I__18498 (
            .O(N__75481),
            .I(N__75464));
    LocalMux I__18497 (
            .O(N__75476),
            .I(N__75461));
    LocalMux I__18496 (
            .O(N__75473),
            .I(N__75458));
    Span4Mux_h I__18495 (
            .O(N__75470),
            .I(N__75455));
    Span4Mux_v I__18494 (
            .O(N__75467),
            .I(N__75452));
    Span4Mux_v I__18493 (
            .O(N__75464),
            .I(N__75449));
    Span4Mux_h I__18492 (
            .O(N__75461),
            .I(N__75442));
    Span4Mux_h I__18491 (
            .O(N__75458),
            .I(N__75442));
    Span4Mux_v I__18490 (
            .O(N__75455),
            .I(N__75442));
    Span4Mux_v I__18489 (
            .O(N__75452),
            .I(N__75439));
    Span4Mux_h I__18488 (
            .O(N__75449),
            .I(N__75436));
    Span4Mux_v I__18487 (
            .O(N__75442),
            .I(N__75433));
    Odrv4 I__18486 (
            .O(N__75439),
            .I(\c0.n12_adj_4672 ));
    Odrv4 I__18485 (
            .O(N__75436),
            .I(\c0.n12_adj_4672 ));
    Odrv4 I__18484 (
            .O(N__75433),
            .I(\c0.n12_adj_4672 ));
    CascadeMux I__18483 (
            .O(N__75426),
            .I(N__75423));
    InMux I__18482 (
            .O(N__75423),
            .I(N__75417));
    InMux I__18481 (
            .O(N__75422),
            .I(N__75408));
    InMux I__18480 (
            .O(N__75421),
            .I(N__75408));
    InMux I__18479 (
            .O(N__75420),
            .I(N__75408));
    LocalMux I__18478 (
            .O(N__75417),
            .I(N__75403));
    InMux I__18477 (
            .O(N__75416),
            .I(N__75400));
    InMux I__18476 (
            .O(N__75415),
            .I(N__75394));
    LocalMux I__18475 (
            .O(N__75408),
            .I(N__75390));
    InMux I__18474 (
            .O(N__75407),
            .I(N__75385));
    InMux I__18473 (
            .O(N__75406),
            .I(N__75385));
    Span4Mux_h I__18472 (
            .O(N__75403),
            .I(N__75380));
    LocalMux I__18471 (
            .O(N__75400),
            .I(N__75380));
    InMux I__18470 (
            .O(N__75399),
            .I(N__75375));
    InMux I__18469 (
            .O(N__75398),
            .I(N__75375));
    InMux I__18468 (
            .O(N__75397),
            .I(N__75370));
    LocalMux I__18467 (
            .O(N__75394),
            .I(N__75367));
    InMux I__18466 (
            .O(N__75393),
            .I(N__75364));
    Span4Mux_h I__18465 (
            .O(N__75390),
            .I(N__75359));
    LocalMux I__18464 (
            .O(N__75385),
            .I(N__75359));
    Span4Mux_h I__18463 (
            .O(N__75380),
            .I(N__75356));
    LocalMux I__18462 (
            .O(N__75375),
            .I(N__75353));
    InMux I__18461 (
            .O(N__75374),
            .I(N__75350));
    InMux I__18460 (
            .O(N__75373),
            .I(N__75347));
    LocalMux I__18459 (
            .O(N__75370),
            .I(N__75344));
    Span4Mux_h I__18458 (
            .O(N__75367),
            .I(N__75341));
    LocalMux I__18457 (
            .O(N__75364),
            .I(N__75338));
    Span4Mux_v I__18456 (
            .O(N__75359),
            .I(N__75334));
    Sp12to4 I__18455 (
            .O(N__75356),
            .I(N__75331));
    Span4Mux_v I__18454 (
            .O(N__75353),
            .I(N__75328));
    LocalMux I__18453 (
            .O(N__75350),
            .I(N__75321));
    LocalMux I__18452 (
            .O(N__75347),
            .I(N__75321));
    Span4Mux_v I__18451 (
            .O(N__75344),
            .I(N__75318));
    Span4Mux_h I__18450 (
            .O(N__75341),
            .I(N__75313));
    Span4Mux_v I__18449 (
            .O(N__75338),
            .I(N__75313));
    InMux I__18448 (
            .O(N__75337),
            .I(N__75310));
    Sp12to4 I__18447 (
            .O(N__75334),
            .I(N__75307));
    Span12Mux_v I__18446 (
            .O(N__75331),
            .I(N__75302));
    Sp12to4 I__18445 (
            .O(N__75328),
            .I(N__75302));
    InMux I__18444 (
            .O(N__75327),
            .I(N__75298));
    InMux I__18443 (
            .O(N__75326),
            .I(N__75295));
    Span4Mux_h I__18442 (
            .O(N__75321),
            .I(N__75290));
    Span4Mux_v I__18441 (
            .O(N__75318),
            .I(N__75290));
    Span4Mux_v I__18440 (
            .O(N__75313),
            .I(N__75287));
    LocalMux I__18439 (
            .O(N__75310),
            .I(N__75280));
    Span12Mux_h I__18438 (
            .O(N__75307),
            .I(N__75280));
    Span12Mux_h I__18437 (
            .O(N__75302),
            .I(N__75280));
    InMux I__18436 (
            .O(N__75301),
            .I(N__75277));
    LocalMux I__18435 (
            .O(N__75298),
            .I(N__75274));
    LocalMux I__18434 (
            .O(N__75295),
            .I(\c0.n22099 ));
    Odrv4 I__18433 (
            .O(N__75290),
            .I(\c0.n22099 ));
    Odrv4 I__18432 (
            .O(N__75287),
            .I(\c0.n22099 ));
    Odrv12 I__18431 (
            .O(N__75280),
            .I(\c0.n22099 ));
    LocalMux I__18430 (
            .O(N__75277),
            .I(\c0.n22099 ));
    Odrv12 I__18429 (
            .O(N__75274),
            .I(\c0.n22099 ));
    InMux I__18428 (
            .O(N__75261),
            .I(N__75258));
    LocalMux I__18427 (
            .O(N__75258),
            .I(N__75245));
    InMux I__18426 (
            .O(N__75257),
            .I(N__75239));
    InMux I__18425 (
            .O(N__75256),
            .I(N__75236));
    InMux I__18424 (
            .O(N__75255),
            .I(N__75233));
    CascadeMux I__18423 (
            .O(N__75254),
            .I(N__75230));
    InMux I__18422 (
            .O(N__75253),
            .I(N__75225));
    InMux I__18421 (
            .O(N__75252),
            .I(N__75219));
    InMux I__18420 (
            .O(N__75251),
            .I(N__75219));
    InMux I__18419 (
            .O(N__75250),
            .I(N__75216));
    InMux I__18418 (
            .O(N__75249),
            .I(N__75211));
    InMux I__18417 (
            .O(N__75248),
            .I(N__75211));
    Span4Mux_v I__18416 (
            .O(N__75245),
            .I(N__75208));
    InMux I__18415 (
            .O(N__75244),
            .I(N__75205));
    InMux I__18414 (
            .O(N__75243),
            .I(N__75202));
    InMux I__18413 (
            .O(N__75242),
            .I(N__75199));
    LocalMux I__18412 (
            .O(N__75239),
            .I(N__75196));
    LocalMux I__18411 (
            .O(N__75236),
            .I(N__75190));
    LocalMux I__18410 (
            .O(N__75233),
            .I(N__75190));
    InMux I__18409 (
            .O(N__75230),
            .I(N__75187));
    CascadeMux I__18408 (
            .O(N__75229),
            .I(N__75182));
    CascadeMux I__18407 (
            .O(N__75228),
            .I(N__75179));
    LocalMux I__18406 (
            .O(N__75225),
            .I(N__75174));
    InMux I__18405 (
            .O(N__75224),
            .I(N__75171));
    LocalMux I__18404 (
            .O(N__75219),
            .I(N__75166));
    LocalMux I__18403 (
            .O(N__75216),
            .I(N__75166));
    LocalMux I__18402 (
            .O(N__75211),
            .I(N__75163));
    Span4Mux_h I__18401 (
            .O(N__75208),
            .I(N__75160));
    LocalMux I__18400 (
            .O(N__75205),
            .I(N__75153));
    LocalMux I__18399 (
            .O(N__75202),
            .I(N__75153));
    LocalMux I__18398 (
            .O(N__75199),
            .I(N__75153));
    Span4Mux_h I__18397 (
            .O(N__75196),
            .I(N__75150));
    InMux I__18396 (
            .O(N__75195),
            .I(N__75147));
    Span4Mux_v I__18395 (
            .O(N__75190),
            .I(N__75142));
    LocalMux I__18394 (
            .O(N__75187),
            .I(N__75142));
    InMux I__18393 (
            .O(N__75186),
            .I(N__75139));
    InMux I__18392 (
            .O(N__75185),
            .I(N__75134));
    InMux I__18391 (
            .O(N__75182),
            .I(N__75131));
    InMux I__18390 (
            .O(N__75179),
            .I(N__75128));
    InMux I__18389 (
            .O(N__75178),
            .I(N__75125));
    InMux I__18388 (
            .O(N__75177),
            .I(N__75122));
    Span4Mux_v I__18387 (
            .O(N__75174),
            .I(N__75117));
    LocalMux I__18386 (
            .O(N__75171),
            .I(N__75117));
    Span4Mux_h I__18385 (
            .O(N__75166),
            .I(N__75114));
    Span4Mux_v I__18384 (
            .O(N__75163),
            .I(N__75103));
    Span4Mux_h I__18383 (
            .O(N__75160),
            .I(N__75103));
    Span4Mux_v I__18382 (
            .O(N__75153),
            .I(N__75103));
    Span4Mux_h I__18381 (
            .O(N__75150),
            .I(N__75098));
    LocalMux I__18380 (
            .O(N__75147),
            .I(N__75098));
    Span4Mux_v I__18379 (
            .O(N__75142),
            .I(N__75093));
    LocalMux I__18378 (
            .O(N__75139),
            .I(N__75093));
    InMux I__18377 (
            .O(N__75138),
            .I(N__75088));
    InMux I__18376 (
            .O(N__75137),
            .I(N__75088));
    LocalMux I__18375 (
            .O(N__75134),
            .I(N__75085));
    LocalMux I__18374 (
            .O(N__75131),
            .I(N__75080));
    LocalMux I__18373 (
            .O(N__75128),
            .I(N__75080));
    LocalMux I__18372 (
            .O(N__75125),
            .I(N__75077));
    LocalMux I__18371 (
            .O(N__75122),
            .I(N__75074));
    Span4Mux_v I__18370 (
            .O(N__75117),
            .I(N__75071));
    Span4Mux_v I__18369 (
            .O(N__75114),
            .I(N__75068));
    InMux I__18368 (
            .O(N__75113),
            .I(N__75065));
    InMux I__18367 (
            .O(N__75112),
            .I(N__75062));
    InMux I__18366 (
            .O(N__75111),
            .I(N__75057));
    InMux I__18365 (
            .O(N__75110),
            .I(N__75057));
    Sp12to4 I__18364 (
            .O(N__75103),
            .I(N__75054));
    Span4Mux_h I__18363 (
            .O(N__75098),
            .I(N__75051));
    Span4Mux_h I__18362 (
            .O(N__75093),
            .I(N__75048));
    LocalMux I__18361 (
            .O(N__75088),
            .I(N__75041));
    Span4Mux_h I__18360 (
            .O(N__75085),
            .I(N__75041));
    Span4Mux_v I__18359 (
            .O(N__75080),
            .I(N__75034));
    Span4Mux_v I__18358 (
            .O(N__75077),
            .I(N__75034));
    Span4Mux_v I__18357 (
            .O(N__75074),
            .I(N__75034));
    Span4Mux_h I__18356 (
            .O(N__75071),
            .I(N__75029));
    Span4Mux_v I__18355 (
            .O(N__75068),
            .I(N__75029));
    LocalMux I__18354 (
            .O(N__75065),
            .I(N__75022));
    LocalMux I__18353 (
            .O(N__75062),
            .I(N__75022));
    LocalMux I__18352 (
            .O(N__75057),
            .I(N__75019));
    Span12Mux_h I__18351 (
            .O(N__75054),
            .I(N__75012));
    Sp12to4 I__18350 (
            .O(N__75051),
            .I(N__75012));
    Sp12to4 I__18349 (
            .O(N__75048),
            .I(N__75012));
    InMux I__18348 (
            .O(N__75047),
            .I(N__75007));
    InMux I__18347 (
            .O(N__75046),
            .I(N__75007));
    Span4Mux_v I__18346 (
            .O(N__75041),
            .I(N__75002));
    Span4Mux_h I__18345 (
            .O(N__75034),
            .I(N__75002));
    Sp12to4 I__18344 (
            .O(N__75029),
            .I(N__74999));
    InMux I__18343 (
            .O(N__75028),
            .I(N__74996));
    InMux I__18342 (
            .O(N__75027),
            .I(N__74993));
    Span4Mux_v I__18341 (
            .O(N__75022),
            .I(N__74990));
    Span4Mux_h I__18340 (
            .O(N__75019),
            .I(N__74987));
    Span12Mux_v I__18339 (
            .O(N__75012),
            .I(N__74984));
    LocalMux I__18338 (
            .O(N__75007),
            .I(N__74977));
    Sp12to4 I__18337 (
            .O(N__75002),
            .I(N__74977));
    Span12Mux_s6_h I__18336 (
            .O(N__74999),
            .I(N__74977));
    LocalMux I__18335 (
            .O(N__74996),
            .I(rx_data_1));
    LocalMux I__18334 (
            .O(N__74993),
            .I(rx_data_1));
    Odrv4 I__18333 (
            .O(N__74990),
            .I(rx_data_1));
    Odrv4 I__18332 (
            .O(N__74987),
            .I(rx_data_1));
    Odrv12 I__18331 (
            .O(N__74984),
            .I(rx_data_1));
    Odrv12 I__18330 (
            .O(N__74977),
            .I(rx_data_1));
    CascadeMux I__18329 (
            .O(N__74964),
            .I(N__74958));
    CascadeMux I__18328 (
            .O(N__74963),
            .I(N__74955));
    InMux I__18327 (
            .O(N__74962),
            .I(N__74952));
    InMux I__18326 (
            .O(N__74961),
            .I(N__74949));
    InMux I__18325 (
            .O(N__74958),
            .I(N__74946));
    InMux I__18324 (
            .O(N__74955),
            .I(N__74943));
    LocalMux I__18323 (
            .O(N__74952),
            .I(N__74940));
    LocalMux I__18322 (
            .O(N__74949),
            .I(N__74937));
    LocalMux I__18321 (
            .O(N__74946),
            .I(N__74934));
    LocalMux I__18320 (
            .O(N__74943),
            .I(N__74930));
    Span4Mux_h I__18319 (
            .O(N__74940),
            .I(N__74927));
    Span4Mux_v I__18318 (
            .O(N__74937),
            .I(N__74922));
    Span4Mux_v I__18317 (
            .O(N__74934),
            .I(N__74922));
    InMux I__18316 (
            .O(N__74933),
            .I(N__74919));
    Span4Mux_h I__18315 (
            .O(N__74930),
            .I(N__74914));
    Span4Mux_v I__18314 (
            .O(N__74927),
            .I(N__74914));
    Span4Mux_h I__18313 (
            .O(N__74922),
            .I(N__74911));
    LocalMux I__18312 (
            .O(N__74919),
            .I(\c0.data_in_frame_13_1 ));
    Odrv4 I__18311 (
            .O(N__74914),
            .I(\c0.data_in_frame_13_1 ));
    Odrv4 I__18310 (
            .O(N__74911),
            .I(\c0.data_in_frame_13_1 ));
    InMux I__18309 (
            .O(N__74904),
            .I(N__74900));
    InMux I__18308 (
            .O(N__74903),
            .I(N__74897));
    LocalMux I__18307 (
            .O(N__74900),
            .I(N__74894));
    LocalMux I__18306 (
            .O(N__74897),
            .I(N__74890));
    Span4Mux_v I__18305 (
            .O(N__74894),
            .I(N__74887));
    InMux I__18304 (
            .O(N__74893),
            .I(N__74884));
    Span4Mux_h I__18303 (
            .O(N__74890),
            .I(N__74881));
    Odrv4 I__18302 (
            .O(N__74887),
            .I(\c0.n13490 ));
    LocalMux I__18301 (
            .O(N__74884),
            .I(\c0.n13490 ));
    Odrv4 I__18300 (
            .O(N__74881),
            .I(\c0.n13490 ));
    InMux I__18299 (
            .O(N__74874),
            .I(N__74871));
    LocalMux I__18298 (
            .O(N__74871),
            .I(N__74867));
    CascadeMux I__18297 (
            .O(N__74870),
            .I(N__74863));
    Span4Mux_h I__18296 (
            .O(N__74867),
            .I(N__74860));
    CascadeMux I__18295 (
            .O(N__74866),
            .I(N__74857));
    InMux I__18294 (
            .O(N__74863),
            .I(N__74854));
    Span4Mux_h I__18293 (
            .O(N__74860),
            .I(N__74851));
    InMux I__18292 (
            .O(N__74857),
            .I(N__74848));
    LocalMux I__18291 (
            .O(N__74854),
            .I(\c0.data_in_frame_24_5 ));
    Odrv4 I__18290 (
            .O(N__74851),
            .I(\c0.data_in_frame_24_5 ));
    LocalMux I__18289 (
            .O(N__74848),
            .I(\c0.data_in_frame_24_5 ));
    InMux I__18288 (
            .O(N__74841),
            .I(N__74838));
    LocalMux I__18287 (
            .O(N__74838),
            .I(N__74834));
    InMux I__18286 (
            .O(N__74837),
            .I(N__74831));
    Span4Mux_h I__18285 (
            .O(N__74834),
            .I(N__74828));
    LocalMux I__18284 (
            .O(N__74831),
            .I(N__74825));
    Span4Mux_h I__18283 (
            .O(N__74828),
            .I(N__74822));
    Odrv4 I__18282 (
            .O(N__74825),
            .I(\c0.n22505 ));
    Odrv4 I__18281 (
            .O(N__74822),
            .I(\c0.n22505 ));
    InMux I__18280 (
            .O(N__74817),
            .I(N__74812));
    InMux I__18279 (
            .O(N__74816),
            .I(N__74808));
    InMux I__18278 (
            .O(N__74815),
            .I(N__74805));
    LocalMux I__18277 (
            .O(N__74812),
            .I(N__74802));
    InMux I__18276 (
            .O(N__74811),
            .I(N__74799));
    LocalMux I__18275 (
            .O(N__74808),
            .I(N__74794));
    LocalMux I__18274 (
            .O(N__74805),
            .I(N__74794));
    Span4Mux_v I__18273 (
            .O(N__74802),
            .I(N__74789));
    LocalMux I__18272 (
            .O(N__74799),
            .I(N__74789));
    Span4Mux_v I__18271 (
            .O(N__74794),
            .I(N__74786));
    Span4Mux_h I__18270 (
            .O(N__74789),
            .I(N__74783));
    Odrv4 I__18269 (
            .O(N__74786),
            .I(\c0.n6718 ));
    Odrv4 I__18268 (
            .O(N__74783),
            .I(\c0.n6718 ));
    InMux I__18267 (
            .O(N__74778),
            .I(N__74775));
    LocalMux I__18266 (
            .O(N__74775),
            .I(N__74769));
    CascadeMux I__18265 (
            .O(N__74774),
            .I(N__74765));
    InMux I__18264 (
            .O(N__74773),
            .I(N__74760));
    InMux I__18263 (
            .O(N__74772),
            .I(N__74760));
    Span4Mux_h I__18262 (
            .O(N__74769),
            .I(N__74757));
    InMux I__18261 (
            .O(N__74768),
            .I(N__74752));
    InMux I__18260 (
            .O(N__74765),
            .I(N__74752));
    LocalMux I__18259 (
            .O(N__74760),
            .I(\c0.n13963 ));
    Odrv4 I__18258 (
            .O(N__74757),
            .I(\c0.n13963 ));
    LocalMux I__18257 (
            .O(N__74752),
            .I(\c0.n13963 ));
    InMux I__18256 (
            .O(N__74745),
            .I(N__74742));
    LocalMux I__18255 (
            .O(N__74742),
            .I(N__74739));
    Span4Mux_v I__18254 (
            .O(N__74739),
            .I(N__74736));
    Odrv4 I__18253 (
            .O(N__74736),
            .I(\c0.n21295 ));
    InMux I__18252 (
            .O(N__74733),
            .I(N__74730));
    LocalMux I__18251 (
            .O(N__74730),
            .I(N__74727));
    Span4Mux_h I__18250 (
            .O(N__74727),
            .I(N__74724));
    Span4Mux_h I__18249 (
            .O(N__74724),
            .I(N__74721));
    Odrv4 I__18248 (
            .O(N__74721),
            .I(\c0.n20239 ));
    CascadeMux I__18247 (
            .O(N__74718),
            .I(N__74715));
    InMux I__18246 (
            .O(N__74715),
            .I(N__74709));
    InMux I__18245 (
            .O(N__74714),
            .I(N__74704));
    InMux I__18244 (
            .O(N__74713),
            .I(N__74704));
    CascadeMux I__18243 (
            .O(N__74712),
            .I(N__74701));
    LocalMux I__18242 (
            .O(N__74709),
            .I(N__74698));
    LocalMux I__18241 (
            .O(N__74704),
            .I(N__74695));
    InMux I__18240 (
            .O(N__74701),
            .I(N__74692));
    Span12Mux_h I__18239 (
            .O(N__74698),
            .I(N__74689));
    Span4Mux_h I__18238 (
            .O(N__74695),
            .I(N__74686));
    LocalMux I__18237 (
            .O(N__74692),
            .I(\c0.data_in_frame_17_1 ));
    Odrv12 I__18236 (
            .O(N__74689),
            .I(\c0.data_in_frame_17_1 ));
    Odrv4 I__18235 (
            .O(N__74686),
            .I(\c0.data_in_frame_17_1 ));
    InMux I__18234 (
            .O(N__74679),
            .I(N__74675));
    InMux I__18233 (
            .O(N__74678),
            .I(N__74670));
    LocalMux I__18232 (
            .O(N__74675),
            .I(N__74667));
    CascadeMux I__18231 (
            .O(N__74674),
            .I(N__74663));
    InMux I__18230 (
            .O(N__74673),
            .I(N__74660));
    LocalMux I__18229 (
            .O(N__74670),
            .I(N__74655));
    Span4Mux_v I__18228 (
            .O(N__74667),
            .I(N__74652));
    InMux I__18227 (
            .O(N__74666),
            .I(N__74647));
    InMux I__18226 (
            .O(N__74663),
            .I(N__74647));
    LocalMux I__18225 (
            .O(N__74660),
            .I(N__74644));
    InMux I__18224 (
            .O(N__74659),
            .I(N__74637));
    InMux I__18223 (
            .O(N__74658),
            .I(N__74637));
    Span4Mux_h I__18222 (
            .O(N__74655),
            .I(N__74633));
    Sp12to4 I__18221 (
            .O(N__74652),
            .I(N__74626));
    LocalMux I__18220 (
            .O(N__74647),
            .I(N__74626));
    Span4Mux_h I__18219 (
            .O(N__74644),
            .I(N__74622));
    InMux I__18218 (
            .O(N__74643),
            .I(N__74619));
    InMux I__18217 (
            .O(N__74642),
            .I(N__74616));
    LocalMux I__18216 (
            .O(N__74637),
            .I(N__74613));
    InMux I__18215 (
            .O(N__74636),
            .I(N__74610));
    Sp12to4 I__18214 (
            .O(N__74633),
            .I(N__74607));
    InMux I__18213 (
            .O(N__74632),
            .I(N__74604));
    InMux I__18212 (
            .O(N__74631),
            .I(N__74601));
    Span12Mux_h I__18211 (
            .O(N__74626),
            .I(N__74598));
    InMux I__18210 (
            .O(N__74625),
            .I(N__74595));
    Span4Mux_v I__18209 (
            .O(N__74622),
            .I(N__74592));
    LocalMux I__18208 (
            .O(N__74619),
            .I(N__74589));
    LocalMux I__18207 (
            .O(N__74616),
            .I(N__74586));
    Span4Mux_v I__18206 (
            .O(N__74613),
            .I(N__74581));
    LocalMux I__18205 (
            .O(N__74610),
            .I(N__74581));
    Span12Mux_v I__18204 (
            .O(N__74607),
            .I(N__74578));
    LocalMux I__18203 (
            .O(N__74604),
            .I(N__74573));
    LocalMux I__18202 (
            .O(N__74601),
            .I(N__74573));
    Span12Mux_v I__18201 (
            .O(N__74598),
            .I(N__74570));
    LocalMux I__18200 (
            .O(N__74595),
            .I(N__74563));
    Span4Mux_v I__18199 (
            .O(N__74592),
            .I(N__74563));
    Span4Mux_h I__18198 (
            .O(N__74589),
            .I(N__74563));
    Span4Mux_v I__18197 (
            .O(N__74586),
            .I(N__74559));
    Span4Mux_v I__18196 (
            .O(N__74581),
            .I(N__74556));
    Span12Mux_v I__18195 (
            .O(N__74578),
            .I(N__74553));
    Span12Mux_h I__18194 (
            .O(N__74573),
            .I(N__74548));
    Span12Mux_h I__18193 (
            .O(N__74570),
            .I(N__74548));
    Span4Mux_v I__18192 (
            .O(N__74563),
            .I(N__74545));
    InMux I__18191 (
            .O(N__74562),
            .I(N__74542));
    Odrv4 I__18190 (
            .O(N__74559),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__18189 (
            .O(N__74556),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv12 I__18188 (
            .O(N__74553),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv12 I__18187 (
            .O(N__74548),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__18186 (
            .O(N__74545),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__18185 (
            .O(N__74542),
            .I(\c0.FRAME_MATCHER_i_2 ));
    InMux I__18184 (
            .O(N__74529),
            .I(N__74526));
    LocalMux I__18183 (
            .O(N__74526),
            .I(N__74521));
    InMux I__18182 (
            .O(N__74525),
            .I(N__74517));
    InMux I__18181 (
            .O(N__74524),
            .I(N__74514));
    Span4Mux_v I__18180 (
            .O(N__74521),
            .I(N__74511));
    InMux I__18179 (
            .O(N__74520),
            .I(N__74508));
    LocalMux I__18178 (
            .O(N__74517),
            .I(N__74504));
    LocalMux I__18177 (
            .O(N__74514),
            .I(N__74501));
    Span4Mux_h I__18176 (
            .O(N__74511),
            .I(N__74493));
    LocalMux I__18175 (
            .O(N__74508),
            .I(N__74493));
    InMux I__18174 (
            .O(N__74507),
            .I(N__74490));
    Span4Mux_v I__18173 (
            .O(N__74504),
            .I(N__74487));
    Span4Mux_v I__18172 (
            .O(N__74501),
            .I(N__74484));
    InMux I__18171 (
            .O(N__74500),
            .I(N__74481));
    InMux I__18170 (
            .O(N__74499),
            .I(N__74477));
    InMux I__18169 (
            .O(N__74498),
            .I(N__74474));
    Span4Mux_v I__18168 (
            .O(N__74493),
            .I(N__74471));
    LocalMux I__18167 (
            .O(N__74490),
            .I(N__74466));
    Span4Mux_h I__18166 (
            .O(N__74487),
            .I(N__74459));
    Span4Mux_v I__18165 (
            .O(N__74484),
            .I(N__74459));
    LocalMux I__18164 (
            .O(N__74481),
            .I(N__74459));
    InMux I__18163 (
            .O(N__74480),
            .I(N__74456));
    LocalMux I__18162 (
            .O(N__74477),
            .I(N__74453));
    LocalMux I__18161 (
            .O(N__74474),
            .I(N__74448));
    Span4Mux_v I__18160 (
            .O(N__74471),
            .I(N__74448));
    InMux I__18159 (
            .O(N__74470),
            .I(N__74442));
    InMux I__18158 (
            .O(N__74469),
            .I(N__74442));
    Span4Mux_v I__18157 (
            .O(N__74466),
            .I(N__74436));
    Span4Mux_v I__18156 (
            .O(N__74459),
            .I(N__74436));
    LocalMux I__18155 (
            .O(N__74456),
            .I(N__74429));
    Span4Mux_h I__18154 (
            .O(N__74453),
            .I(N__74429));
    Span4Mux_v I__18153 (
            .O(N__74448),
            .I(N__74429));
    InMux I__18152 (
            .O(N__74447),
            .I(N__74426));
    LocalMux I__18151 (
            .O(N__74442),
            .I(N__74423));
    InMux I__18150 (
            .O(N__74441),
            .I(N__74420));
    Span4Mux_h I__18149 (
            .O(N__74436),
            .I(N__74417));
    Span4Mux_v I__18148 (
            .O(N__74429),
            .I(N__74414));
    LocalMux I__18147 (
            .O(N__74426),
            .I(N__74407));
    Span12Mux_v I__18146 (
            .O(N__74423),
            .I(N__74407));
    LocalMux I__18145 (
            .O(N__74420),
            .I(N__74407));
    Span4Mux_v I__18144 (
            .O(N__74417),
            .I(N__74403));
    Sp12to4 I__18143 (
            .O(N__74414),
            .I(N__74398));
    Span12Mux_v I__18142 (
            .O(N__74407),
            .I(N__74398));
    InMux I__18141 (
            .O(N__74406),
            .I(N__74395));
    Odrv4 I__18140 (
            .O(N__74403),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv12 I__18139 (
            .O(N__74398),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__18138 (
            .O(N__74395),
            .I(\c0.FRAME_MATCHER_i_1 ));
    CascadeMux I__18137 (
            .O(N__74388),
            .I(N__74383));
    CascadeMux I__18136 (
            .O(N__74387),
            .I(N__74378));
    CascadeMux I__18135 (
            .O(N__74386),
            .I(N__74375));
    InMux I__18134 (
            .O(N__74383),
            .I(N__74372));
    InMux I__18133 (
            .O(N__74382),
            .I(N__74369));
    CascadeMux I__18132 (
            .O(N__74381),
            .I(N__74366));
    InMux I__18131 (
            .O(N__74378),
            .I(N__74362));
    InMux I__18130 (
            .O(N__74375),
            .I(N__74359));
    LocalMux I__18129 (
            .O(N__74372),
            .I(N__74355));
    LocalMux I__18128 (
            .O(N__74369),
            .I(N__74352));
    InMux I__18127 (
            .O(N__74366),
            .I(N__74349));
    InMux I__18126 (
            .O(N__74365),
            .I(N__74345));
    LocalMux I__18125 (
            .O(N__74362),
            .I(N__74341));
    LocalMux I__18124 (
            .O(N__74359),
            .I(N__74338));
    InMux I__18123 (
            .O(N__74358),
            .I(N__74335));
    Span4Mux_h I__18122 (
            .O(N__74355),
            .I(N__74332));
    Span4Mux_v I__18121 (
            .O(N__74352),
            .I(N__74329));
    LocalMux I__18120 (
            .O(N__74349),
            .I(N__74326));
    InMux I__18119 (
            .O(N__74348),
            .I(N__74323));
    LocalMux I__18118 (
            .O(N__74345),
            .I(N__74320));
    InMux I__18117 (
            .O(N__74344),
            .I(N__74317));
    Span4Mux_v I__18116 (
            .O(N__74341),
            .I(N__74312));
    Span4Mux_h I__18115 (
            .O(N__74338),
            .I(N__74312));
    LocalMux I__18114 (
            .O(N__74335),
            .I(N__74309));
    Span4Mux_h I__18113 (
            .O(N__74332),
            .I(N__74306));
    Span4Mux_v I__18112 (
            .O(N__74329),
            .I(N__74303));
    Span4Mux_v I__18111 (
            .O(N__74326),
            .I(N__74297));
    LocalMux I__18110 (
            .O(N__74323),
            .I(N__74297));
    Span4Mux_v I__18109 (
            .O(N__74320),
            .I(N__74292));
    LocalMux I__18108 (
            .O(N__74317),
            .I(N__74292));
    Span4Mux_v I__18107 (
            .O(N__74312),
            .I(N__74289));
    Span4Mux_h I__18106 (
            .O(N__74309),
            .I(N__74285));
    Span4Mux_v I__18105 (
            .O(N__74306),
            .I(N__74280));
    Span4Mux_h I__18104 (
            .O(N__74303),
            .I(N__74280));
    InMux I__18103 (
            .O(N__74302),
            .I(N__74276));
    Span4Mux_v I__18102 (
            .O(N__74297),
            .I(N__74273));
    Span4Mux_v I__18101 (
            .O(N__74292),
            .I(N__74270));
    Span4Mux_v I__18100 (
            .O(N__74289),
            .I(N__74267));
    InMux I__18099 (
            .O(N__74288),
            .I(N__74264));
    Span4Mux_h I__18098 (
            .O(N__74285),
            .I(N__74259));
    Span4Mux_v I__18097 (
            .O(N__74280),
            .I(N__74259));
    InMux I__18096 (
            .O(N__74279),
            .I(N__74256));
    LocalMux I__18095 (
            .O(N__74276),
            .I(N__74247));
    Span4Mux_h I__18094 (
            .O(N__74273),
            .I(N__74247));
    Span4Mux_h I__18093 (
            .O(N__74270),
            .I(N__74247));
    Span4Mux_v I__18092 (
            .O(N__74267),
            .I(N__74247));
    LocalMux I__18091 (
            .O(N__74264),
            .I(N__74242));
    Span4Mux_v I__18090 (
            .O(N__74259),
            .I(N__74242));
    LocalMux I__18089 (
            .O(N__74256),
            .I(N__74239));
    Span4Mux_v I__18088 (
            .O(N__74247),
            .I(N__74235));
    Sp12to4 I__18087 (
            .O(N__74242),
            .I(N__74230));
    Span12Mux_h I__18086 (
            .O(N__74239),
            .I(N__74230));
    InMux I__18085 (
            .O(N__74238),
            .I(N__74227));
    Odrv4 I__18084 (
            .O(N__74235),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv12 I__18083 (
            .O(N__74230),
            .I(\c0.FRAME_MATCHER_i_0 ));
    LocalMux I__18082 (
            .O(N__74227),
            .I(\c0.FRAME_MATCHER_i_0 ));
    InMux I__18081 (
            .O(N__74220),
            .I(N__74217));
    LocalMux I__18080 (
            .O(N__74217),
            .I(N__74213));
    InMux I__18079 (
            .O(N__74216),
            .I(N__74210));
    Span4Mux_h I__18078 (
            .O(N__74213),
            .I(N__74197));
    LocalMux I__18077 (
            .O(N__74210),
            .I(N__74197));
    InMux I__18076 (
            .O(N__74209),
            .I(N__74194));
    InMux I__18075 (
            .O(N__74208),
            .I(N__74189));
    InMux I__18074 (
            .O(N__74207),
            .I(N__74189));
    InMux I__18073 (
            .O(N__74206),
            .I(N__74184));
    InMux I__18072 (
            .O(N__74205),
            .I(N__74181));
    InMux I__18071 (
            .O(N__74204),
            .I(N__74171));
    InMux I__18070 (
            .O(N__74203),
            .I(N__74171));
    InMux I__18069 (
            .O(N__74202),
            .I(N__74171));
    Span4Mux_v I__18068 (
            .O(N__74197),
            .I(N__74166));
    LocalMux I__18067 (
            .O(N__74194),
            .I(N__74166));
    LocalMux I__18066 (
            .O(N__74189),
            .I(N__74163));
    InMux I__18065 (
            .O(N__74188),
            .I(N__74158));
    InMux I__18064 (
            .O(N__74187),
            .I(N__74158));
    LocalMux I__18063 (
            .O(N__74184),
            .I(N__74151));
    LocalMux I__18062 (
            .O(N__74181),
            .I(N__74151));
    InMux I__18061 (
            .O(N__74180),
            .I(N__74147));
    InMux I__18060 (
            .O(N__74179),
            .I(N__74142));
    InMux I__18059 (
            .O(N__74178),
            .I(N__74139));
    LocalMux I__18058 (
            .O(N__74171),
            .I(N__74136));
    Span4Mux_h I__18057 (
            .O(N__74166),
            .I(N__74132));
    Span4Mux_v I__18056 (
            .O(N__74163),
            .I(N__74127));
    LocalMux I__18055 (
            .O(N__74158),
            .I(N__74127));
    InMux I__18054 (
            .O(N__74157),
            .I(N__74124));
    InMux I__18053 (
            .O(N__74156),
            .I(N__74121));
    Span4Mux_h I__18052 (
            .O(N__74151),
            .I(N__74118));
    InMux I__18051 (
            .O(N__74150),
            .I(N__74112));
    LocalMux I__18050 (
            .O(N__74147),
            .I(N__74108));
    InMux I__18049 (
            .O(N__74146),
            .I(N__74105));
    InMux I__18048 (
            .O(N__74145),
            .I(N__74101));
    LocalMux I__18047 (
            .O(N__74142),
            .I(N__74098));
    LocalMux I__18046 (
            .O(N__74139),
            .I(N__74095));
    Span4Mux_v I__18045 (
            .O(N__74136),
            .I(N__74092));
    InMux I__18044 (
            .O(N__74135),
            .I(N__74089));
    Span4Mux_h I__18043 (
            .O(N__74132),
            .I(N__74086));
    Span4Mux_h I__18042 (
            .O(N__74127),
            .I(N__74081));
    LocalMux I__18041 (
            .O(N__74124),
            .I(N__74081));
    LocalMux I__18040 (
            .O(N__74121),
            .I(N__74076));
    Span4Mux_h I__18039 (
            .O(N__74118),
            .I(N__74076));
    InMux I__18038 (
            .O(N__74117),
            .I(N__74073));
    InMux I__18037 (
            .O(N__74116),
            .I(N__74070));
    InMux I__18036 (
            .O(N__74115),
            .I(N__74063));
    LocalMux I__18035 (
            .O(N__74112),
            .I(N__74060));
    InMux I__18034 (
            .O(N__74111),
            .I(N__74057));
    Span4Mux_v I__18033 (
            .O(N__74108),
            .I(N__74052));
    LocalMux I__18032 (
            .O(N__74105),
            .I(N__74052));
    InMux I__18031 (
            .O(N__74104),
            .I(N__74048));
    LocalMux I__18030 (
            .O(N__74101),
            .I(N__74045));
    Span4Mux_v I__18029 (
            .O(N__74098),
            .I(N__74040));
    Span4Mux_v I__18028 (
            .O(N__74095),
            .I(N__74040));
    Sp12to4 I__18027 (
            .O(N__74092),
            .I(N__74035));
    LocalMux I__18026 (
            .O(N__74089),
            .I(N__74035));
    Span4Mux_v I__18025 (
            .O(N__74086),
            .I(N__74030));
    Span4Mux_v I__18024 (
            .O(N__74081),
            .I(N__74030));
    Span4Mux_v I__18023 (
            .O(N__74076),
            .I(N__74025));
    LocalMux I__18022 (
            .O(N__74073),
            .I(N__74025));
    LocalMux I__18021 (
            .O(N__74070),
            .I(N__74022));
    InMux I__18020 (
            .O(N__74069),
            .I(N__74018));
    InMux I__18019 (
            .O(N__74068),
            .I(N__74015));
    InMux I__18018 (
            .O(N__74067),
            .I(N__74010));
    InMux I__18017 (
            .O(N__74066),
            .I(N__74010));
    LocalMux I__18016 (
            .O(N__74063),
            .I(N__74003));
    Span4Mux_h I__18015 (
            .O(N__74060),
            .I(N__74003));
    LocalMux I__18014 (
            .O(N__74057),
            .I(N__74003));
    Span4Mux_h I__18013 (
            .O(N__74052),
            .I(N__74000));
    InMux I__18012 (
            .O(N__74051),
            .I(N__73997));
    LocalMux I__18011 (
            .O(N__74048),
            .I(N__73990));
    Span4Mux_v I__18010 (
            .O(N__74045),
            .I(N__73990));
    Span4Mux_h I__18009 (
            .O(N__74040),
            .I(N__73990));
    Span12Mux_h I__18008 (
            .O(N__74035),
            .I(N__73981));
    Sp12to4 I__18007 (
            .O(N__74030),
            .I(N__73981));
    Sp12to4 I__18006 (
            .O(N__74025),
            .I(N__73981));
    Sp12to4 I__18005 (
            .O(N__74022),
            .I(N__73981));
    InMux I__18004 (
            .O(N__74021),
            .I(N__73978));
    LocalMux I__18003 (
            .O(N__74018),
            .I(N__73975));
    LocalMux I__18002 (
            .O(N__74015),
            .I(N__73972));
    LocalMux I__18001 (
            .O(N__74010),
            .I(N__73967));
    Span4Mux_h I__18000 (
            .O(N__74003),
            .I(N__73967));
    Span4Mux_v I__17999 (
            .O(N__74000),
            .I(N__73964));
    LocalMux I__17998 (
            .O(N__73997),
            .I(N__73957));
    Sp12to4 I__17997 (
            .O(N__73990),
            .I(N__73957));
    Span12Mux_v I__17996 (
            .O(N__73981),
            .I(N__73957));
    LocalMux I__17995 (
            .O(N__73978),
            .I(\c0.n9_adj_4601 ));
    Odrv4 I__17994 (
            .O(N__73975),
            .I(\c0.n9_adj_4601 ));
    Odrv4 I__17993 (
            .O(N__73972),
            .I(\c0.n9_adj_4601 ));
    Odrv4 I__17992 (
            .O(N__73967),
            .I(\c0.n9_adj_4601 ));
    Odrv4 I__17991 (
            .O(N__73964),
            .I(\c0.n9_adj_4601 ));
    Odrv12 I__17990 (
            .O(N__73957),
            .I(\c0.n9_adj_4601 ));
    InMux I__17989 (
            .O(N__73944),
            .I(N__73940));
    InMux I__17988 (
            .O(N__73943),
            .I(N__73936));
    LocalMux I__17987 (
            .O(N__73940),
            .I(N__73933));
    CascadeMux I__17986 (
            .O(N__73939),
            .I(N__73930));
    LocalMux I__17985 (
            .O(N__73936),
            .I(N__73927));
    Span4Mux_v I__17984 (
            .O(N__73933),
            .I(N__73924));
    InMux I__17983 (
            .O(N__73930),
            .I(N__73921));
    Span4Mux_h I__17982 (
            .O(N__73927),
            .I(N__73918));
    Span4Mux_h I__17981 (
            .O(N__73924),
            .I(N__73915));
    LocalMux I__17980 (
            .O(N__73921),
            .I(\c0.data_in_frame_25_1 ));
    Odrv4 I__17979 (
            .O(N__73918),
            .I(\c0.data_in_frame_25_1 ));
    Odrv4 I__17978 (
            .O(N__73915),
            .I(\c0.data_in_frame_25_1 ));
    CascadeMux I__17977 (
            .O(N__73908),
            .I(N__73905));
    InMux I__17976 (
            .O(N__73905),
            .I(N__73902));
    LocalMux I__17975 (
            .O(N__73902),
            .I(N__73896));
    CascadeMux I__17974 (
            .O(N__73901),
            .I(N__73893));
    InMux I__17973 (
            .O(N__73900),
            .I(N__73890));
    InMux I__17972 (
            .O(N__73899),
            .I(N__73887));
    Span4Mux_h I__17971 (
            .O(N__73896),
            .I(N__73884));
    InMux I__17970 (
            .O(N__73893),
            .I(N__73881));
    LocalMux I__17969 (
            .O(N__73890),
            .I(N__73876));
    LocalMux I__17968 (
            .O(N__73887),
            .I(N__73876));
    Span4Mux_v I__17967 (
            .O(N__73884),
            .I(N__73873));
    LocalMux I__17966 (
            .O(N__73881),
            .I(N__73868));
    Span4Mux_v I__17965 (
            .O(N__73876),
            .I(N__73868));
    Odrv4 I__17964 (
            .O(N__73873),
            .I(\c0.data_in_frame_20_0 ));
    Odrv4 I__17963 (
            .O(N__73868),
            .I(\c0.data_in_frame_20_0 ));
    CascadeMux I__17962 (
            .O(N__73863),
            .I(N__73858));
    CascadeMux I__17961 (
            .O(N__73862),
            .I(N__73855));
    CascadeMux I__17960 (
            .O(N__73861),
            .I(N__73851));
    InMux I__17959 (
            .O(N__73858),
            .I(N__73848));
    InMux I__17958 (
            .O(N__73855),
            .I(N__73843));
    InMux I__17957 (
            .O(N__73854),
            .I(N__73843));
    InMux I__17956 (
            .O(N__73851),
            .I(N__73840));
    LocalMux I__17955 (
            .O(N__73848),
            .I(N__73837));
    LocalMux I__17954 (
            .O(N__73843),
            .I(N__73834));
    LocalMux I__17953 (
            .O(N__73840),
            .I(N__73831));
    Span4Mux_v I__17952 (
            .O(N__73837),
            .I(N__73828));
    Span4Mux_h I__17951 (
            .O(N__73834),
            .I(N__73825));
    Span4Mux_h I__17950 (
            .O(N__73831),
            .I(N__73822));
    Span4Mux_h I__17949 (
            .O(N__73828),
            .I(N__73817));
    Span4Mux_h I__17948 (
            .O(N__73825),
            .I(N__73817));
    Span4Mux_h I__17947 (
            .O(N__73822),
            .I(N__73814));
    Odrv4 I__17946 (
            .O(N__73817),
            .I(\c0.data_in_frame_19_0 ));
    Odrv4 I__17945 (
            .O(N__73814),
            .I(\c0.data_in_frame_19_0 ));
    InMux I__17944 (
            .O(N__73809),
            .I(N__73806));
    LocalMux I__17943 (
            .O(N__73806),
            .I(N__73803));
    Span4Mux_h I__17942 (
            .O(N__73803),
            .I(N__73800));
    Odrv4 I__17941 (
            .O(N__73800),
            .I(\c0.n12_adj_4564 ));
    InMux I__17940 (
            .O(N__73797),
            .I(N__73793));
    InMux I__17939 (
            .O(N__73796),
            .I(N__73790));
    LocalMux I__17938 (
            .O(N__73793),
            .I(N__73787));
    LocalMux I__17937 (
            .O(N__73790),
            .I(N__73784));
    Span4Mux_v I__17936 (
            .O(N__73787),
            .I(N__73779));
    Span4Mux_h I__17935 (
            .O(N__73784),
            .I(N__73779));
    Odrv4 I__17934 (
            .O(N__73779),
            .I(\c0.n21404 ));
    CascadeMux I__17933 (
            .O(N__73776),
            .I(\c0.n6_adj_4462_cascade_ ));
    InMux I__17932 (
            .O(N__73773),
            .I(N__73769));
    InMux I__17931 (
            .O(N__73772),
            .I(N__73766));
    LocalMux I__17930 (
            .O(N__73769),
            .I(N__73763));
    LocalMux I__17929 (
            .O(N__73766),
            .I(N__73760));
    Span4Mux_v I__17928 (
            .O(N__73763),
            .I(N__73755));
    Span4Mux_h I__17927 (
            .O(N__73760),
            .I(N__73755));
    Odrv4 I__17926 (
            .O(N__73755),
            .I(\c0.n22562 ));
    CascadeMux I__17925 (
            .O(N__73752),
            .I(N__73747));
    InMux I__17924 (
            .O(N__73751),
            .I(N__73744));
    InMux I__17923 (
            .O(N__73750),
            .I(N__73741));
    InMux I__17922 (
            .O(N__73747),
            .I(N__73738));
    LocalMux I__17921 (
            .O(N__73744),
            .I(N__73735));
    LocalMux I__17920 (
            .O(N__73741),
            .I(N__73727));
    LocalMux I__17919 (
            .O(N__73738),
            .I(N__73727));
    Span4Mux_v I__17918 (
            .O(N__73735),
            .I(N__73727));
    InMux I__17917 (
            .O(N__73734),
            .I(N__73724));
    Odrv4 I__17916 (
            .O(N__73727),
            .I(data_in_frame_22_3));
    LocalMux I__17915 (
            .O(N__73724),
            .I(data_in_frame_22_3));
    CascadeMux I__17914 (
            .O(N__73719),
            .I(N__73711));
    InMux I__17913 (
            .O(N__73718),
            .I(N__73697));
    InMux I__17912 (
            .O(N__73717),
            .I(N__73697));
    InMux I__17911 (
            .O(N__73716),
            .I(N__73681));
    InMux I__17910 (
            .O(N__73715),
            .I(N__73670));
    InMux I__17909 (
            .O(N__73714),
            .I(N__73670));
    InMux I__17908 (
            .O(N__73711),
            .I(N__73670));
    InMux I__17907 (
            .O(N__73710),
            .I(N__73670));
    InMux I__17906 (
            .O(N__73709),
            .I(N__73670));
    InMux I__17905 (
            .O(N__73708),
            .I(N__73662));
    InMux I__17904 (
            .O(N__73707),
            .I(N__73659));
    InMux I__17903 (
            .O(N__73706),
            .I(N__73655));
    InMux I__17902 (
            .O(N__73705),
            .I(N__73652));
    InMux I__17901 (
            .O(N__73704),
            .I(N__73644));
    InMux I__17900 (
            .O(N__73703),
            .I(N__73644));
    InMux I__17899 (
            .O(N__73702),
            .I(N__73644));
    LocalMux I__17898 (
            .O(N__73697),
            .I(N__73641));
    InMux I__17897 (
            .O(N__73696),
            .I(N__73630));
    InMux I__17896 (
            .O(N__73695),
            .I(N__73630));
    InMux I__17895 (
            .O(N__73694),
            .I(N__73630));
    InMux I__17894 (
            .O(N__73693),
            .I(N__73630));
    InMux I__17893 (
            .O(N__73692),
            .I(N__73630));
    InMux I__17892 (
            .O(N__73691),
            .I(N__73623));
    InMux I__17891 (
            .O(N__73690),
            .I(N__73623));
    InMux I__17890 (
            .O(N__73689),
            .I(N__73623));
    InMux I__17889 (
            .O(N__73688),
            .I(N__73620));
    InMux I__17888 (
            .O(N__73687),
            .I(N__73615));
    InMux I__17887 (
            .O(N__73686),
            .I(N__73615));
    CascadeMux I__17886 (
            .O(N__73685),
            .I(N__73612));
    CascadeMux I__17885 (
            .O(N__73684),
            .I(N__73605));
    LocalMux I__17884 (
            .O(N__73681),
            .I(N__73602));
    LocalMux I__17883 (
            .O(N__73670),
            .I(N__73599));
    InMux I__17882 (
            .O(N__73669),
            .I(N__73590));
    InMux I__17881 (
            .O(N__73668),
            .I(N__73590));
    InMux I__17880 (
            .O(N__73667),
            .I(N__73587));
    InMux I__17879 (
            .O(N__73666),
            .I(N__73582));
    InMux I__17878 (
            .O(N__73665),
            .I(N__73582));
    LocalMux I__17877 (
            .O(N__73662),
            .I(N__73579));
    LocalMux I__17876 (
            .O(N__73659),
            .I(N__73576));
    InMux I__17875 (
            .O(N__73658),
            .I(N__73573));
    LocalMux I__17874 (
            .O(N__73655),
            .I(N__73570));
    LocalMux I__17873 (
            .O(N__73652),
            .I(N__73567));
    InMux I__17872 (
            .O(N__73651),
            .I(N__73564));
    LocalMux I__17871 (
            .O(N__73644),
            .I(N__73561));
    Span4Mux_v I__17870 (
            .O(N__73641),
            .I(N__73558));
    LocalMux I__17869 (
            .O(N__73630),
            .I(N__73551));
    LocalMux I__17868 (
            .O(N__73623),
            .I(N__73551));
    LocalMux I__17867 (
            .O(N__73620),
            .I(N__73551));
    LocalMux I__17866 (
            .O(N__73615),
            .I(N__73548));
    InMux I__17865 (
            .O(N__73612),
            .I(N__73543));
    InMux I__17864 (
            .O(N__73611),
            .I(N__73543));
    InMux I__17863 (
            .O(N__73610),
            .I(N__73534));
    InMux I__17862 (
            .O(N__73609),
            .I(N__73534));
    InMux I__17861 (
            .O(N__73608),
            .I(N__73534));
    InMux I__17860 (
            .O(N__73605),
            .I(N__73534));
    Span4Mux_h I__17859 (
            .O(N__73602),
            .I(N__73529));
    Span4Mux_v I__17858 (
            .O(N__73599),
            .I(N__73529));
    InMux I__17857 (
            .O(N__73598),
            .I(N__73526));
    InMux I__17856 (
            .O(N__73597),
            .I(N__73523));
    InMux I__17855 (
            .O(N__73596),
            .I(N__73513));
    InMux I__17854 (
            .O(N__73595),
            .I(N__73513));
    LocalMux I__17853 (
            .O(N__73590),
            .I(N__73506));
    LocalMux I__17852 (
            .O(N__73587),
            .I(N__73506));
    LocalMux I__17851 (
            .O(N__73582),
            .I(N__73506));
    Span4Mux_v I__17850 (
            .O(N__73579),
            .I(N__73503));
    Span4Mux_h I__17849 (
            .O(N__73576),
            .I(N__73500));
    LocalMux I__17848 (
            .O(N__73573),
            .I(N__73497));
    Span4Mux_h I__17847 (
            .O(N__73570),
            .I(N__73492));
    Span4Mux_v I__17846 (
            .O(N__73567),
            .I(N__73492));
    LocalMux I__17845 (
            .O(N__73564),
            .I(N__73489));
    Span4Mux_h I__17844 (
            .O(N__73561),
            .I(N__73484));
    Span4Mux_v I__17843 (
            .O(N__73558),
            .I(N__73484));
    Span4Mux_v I__17842 (
            .O(N__73551),
            .I(N__73479));
    Span4Mux_h I__17841 (
            .O(N__73548),
            .I(N__73479));
    LocalMux I__17840 (
            .O(N__73543),
            .I(N__73472));
    LocalMux I__17839 (
            .O(N__73534),
            .I(N__73472));
    Span4Mux_v I__17838 (
            .O(N__73529),
            .I(N__73472));
    LocalMux I__17837 (
            .O(N__73526),
            .I(N__73467));
    LocalMux I__17836 (
            .O(N__73523),
            .I(N__73467));
    InMux I__17835 (
            .O(N__73522),
            .I(N__73464));
    InMux I__17834 (
            .O(N__73521),
            .I(N__73461));
    InMux I__17833 (
            .O(N__73520),
            .I(N__73458));
    InMux I__17832 (
            .O(N__73519),
            .I(N__73453));
    InMux I__17831 (
            .O(N__73518),
            .I(N__73453));
    LocalMux I__17830 (
            .O(N__73513),
            .I(N__73450));
    Span12Mux_h I__17829 (
            .O(N__73506),
            .I(N__73447));
    Span4Mux_h I__17828 (
            .O(N__73503),
            .I(N__73444));
    Span4Mux_v I__17827 (
            .O(N__73500),
            .I(N__73441));
    Span4Mux_v I__17826 (
            .O(N__73497),
            .I(N__73436));
    Span4Mux_h I__17825 (
            .O(N__73492),
            .I(N__73436));
    Span4Mux_h I__17824 (
            .O(N__73489),
            .I(N__73431));
    Span4Mux_h I__17823 (
            .O(N__73484),
            .I(N__73431));
    Span4Mux_h I__17822 (
            .O(N__73479),
            .I(N__73424));
    Span4Mux_v I__17821 (
            .O(N__73472),
            .I(N__73424));
    Span4Mux_v I__17820 (
            .O(N__73467),
            .I(N__73424));
    LocalMux I__17819 (
            .O(N__73464),
            .I(\c0.n22112 ));
    LocalMux I__17818 (
            .O(N__73461),
            .I(\c0.n22112 ));
    LocalMux I__17817 (
            .O(N__73458),
            .I(\c0.n22112 ));
    LocalMux I__17816 (
            .O(N__73453),
            .I(\c0.n22112 ));
    Odrv12 I__17815 (
            .O(N__73450),
            .I(\c0.n22112 ));
    Odrv12 I__17814 (
            .O(N__73447),
            .I(\c0.n22112 ));
    Odrv4 I__17813 (
            .O(N__73444),
            .I(\c0.n22112 ));
    Odrv4 I__17812 (
            .O(N__73441),
            .I(\c0.n22112 ));
    Odrv4 I__17811 (
            .O(N__73436),
            .I(\c0.n22112 ));
    Odrv4 I__17810 (
            .O(N__73431),
            .I(\c0.n22112 ));
    Odrv4 I__17809 (
            .O(N__73424),
            .I(\c0.n22112 ));
    CascadeMux I__17808 (
            .O(N__73401),
            .I(N__73397));
    InMux I__17807 (
            .O(N__73400),
            .I(N__73393));
    InMux I__17806 (
            .O(N__73397),
            .I(N__73389));
    CascadeMux I__17805 (
            .O(N__73396),
            .I(N__73386));
    LocalMux I__17804 (
            .O(N__73393),
            .I(N__73383));
    InMux I__17803 (
            .O(N__73392),
            .I(N__73380));
    LocalMux I__17802 (
            .O(N__73389),
            .I(N__73377));
    InMux I__17801 (
            .O(N__73386),
            .I(N__73374));
    Span4Mux_h I__17800 (
            .O(N__73383),
            .I(N__73369));
    LocalMux I__17799 (
            .O(N__73380),
            .I(N__73369));
    Span4Mux_h I__17798 (
            .O(N__73377),
            .I(N__73366));
    LocalMux I__17797 (
            .O(N__73374),
            .I(N__73361));
    Span4Mux_v I__17796 (
            .O(N__73369),
            .I(N__73361));
    Odrv4 I__17795 (
            .O(N__73366),
            .I(\c0.data_in_frame_15_0 ));
    Odrv4 I__17794 (
            .O(N__73361),
            .I(\c0.data_in_frame_15_0 ));
    CascadeMux I__17793 (
            .O(N__73356),
            .I(N__73353));
    InMux I__17792 (
            .O(N__73353),
            .I(N__73350));
    LocalMux I__17791 (
            .O(N__73350),
            .I(N__73343));
    InMux I__17790 (
            .O(N__73349),
            .I(N__73338));
    InMux I__17789 (
            .O(N__73348),
            .I(N__73338));
    CascadeMux I__17788 (
            .O(N__73347),
            .I(N__73332));
    InMux I__17787 (
            .O(N__73346),
            .I(N__73327));
    Span4Mux_v I__17786 (
            .O(N__73343),
            .I(N__73321));
    LocalMux I__17785 (
            .O(N__73338),
            .I(N__73321));
    InMux I__17784 (
            .O(N__73337),
            .I(N__73316));
    InMux I__17783 (
            .O(N__73336),
            .I(N__73316));
    InMux I__17782 (
            .O(N__73335),
            .I(N__73313));
    InMux I__17781 (
            .O(N__73332),
            .I(N__73308));
    InMux I__17780 (
            .O(N__73331),
            .I(N__73308));
    InMux I__17779 (
            .O(N__73330),
            .I(N__73304));
    LocalMux I__17778 (
            .O(N__73327),
            .I(N__73301));
    InMux I__17777 (
            .O(N__73326),
            .I(N__73295));
    Span4Mux_v I__17776 (
            .O(N__73321),
            .I(N__73286));
    LocalMux I__17775 (
            .O(N__73316),
            .I(N__73283));
    LocalMux I__17774 (
            .O(N__73313),
            .I(N__73280));
    LocalMux I__17773 (
            .O(N__73308),
            .I(N__73277));
    CascadeMux I__17772 (
            .O(N__73307),
            .I(N__73273));
    LocalMux I__17771 (
            .O(N__73304),
            .I(N__73270));
    Span4Mux_h I__17770 (
            .O(N__73301),
            .I(N__73267));
    InMux I__17769 (
            .O(N__73300),
            .I(N__73264));
    InMux I__17768 (
            .O(N__73299),
            .I(N__73261));
    InMux I__17767 (
            .O(N__73298),
            .I(N__73258));
    LocalMux I__17766 (
            .O(N__73295),
            .I(N__73255));
    InMux I__17765 (
            .O(N__73294),
            .I(N__73250));
    InMux I__17764 (
            .O(N__73293),
            .I(N__73250));
    InMux I__17763 (
            .O(N__73292),
            .I(N__73245));
    InMux I__17762 (
            .O(N__73291),
            .I(N__73245));
    InMux I__17761 (
            .O(N__73290),
            .I(N__73242));
    InMux I__17760 (
            .O(N__73289),
            .I(N__73239));
    Span4Mux_h I__17759 (
            .O(N__73286),
            .I(N__73234));
    Span4Mux_v I__17758 (
            .O(N__73283),
            .I(N__73234));
    Span4Mux_h I__17757 (
            .O(N__73280),
            .I(N__73229));
    Span4Mux_v I__17756 (
            .O(N__73277),
            .I(N__73229));
    InMux I__17755 (
            .O(N__73276),
            .I(N__73226));
    InMux I__17754 (
            .O(N__73273),
            .I(N__73223));
    Span4Mux_h I__17753 (
            .O(N__73270),
            .I(N__73220));
    Span4Mux_v I__17752 (
            .O(N__73267),
            .I(N__73215));
    LocalMux I__17751 (
            .O(N__73264),
            .I(N__73215));
    LocalMux I__17750 (
            .O(N__73261),
            .I(N__73211));
    LocalMux I__17749 (
            .O(N__73258),
            .I(N__73202));
    Span4Mux_h I__17748 (
            .O(N__73255),
            .I(N__73202));
    LocalMux I__17747 (
            .O(N__73250),
            .I(N__73196));
    LocalMux I__17746 (
            .O(N__73245),
            .I(N__73196));
    LocalMux I__17745 (
            .O(N__73242),
            .I(N__73187));
    LocalMux I__17744 (
            .O(N__73239),
            .I(N__73187));
    Span4Mux_h I__17743 (
            .O(N__73234),
            .I(N__73187));
    Span4Mux_v I__17742 (
            .O(N__73229),
            .I(N__73187));
    LocalMux I__17741 (
            .O(N__73226),
            .I(N__73182));
    LocalMux I__17740 (
            .O(N__73223),
            .I(N__73182));
    Span4Mux_v I__17739 (
            .O(N__73220),
            .I(N__73179));
    Span4Mux_h I__17738 (
            .O(N__73215),
            .I(N__73176));
    InMux I__17737 (
            .O(N__73214),
            .I(N__73173));
    Span4Mux_h I__17736 (
            .O(N__73211),
            .I(N__73170));
    InMux I__17735 (
            .O(N__73210),
            .I(N__73167));
    InMux I__17734 (
            .O(N__73209),
            .I(N__73160));
    InMux I__17733 (
            .O(N__73208),
            .I(N__73160));
    InMux I__17732 (
            .O(N__73207),
            .I(N__73160));
    Span4Mux_h I__17731 (
            .O(N__73202),
            .I(N__73157));
    InMux I__17730 (
            .O(N__73201),
            .I(N__73150));
    Span4Mux_v I__17729 (
            .O(N__73196),
            .I(N__73147));
    Span4Mux_v I__17728 (
            .O(N__73187),
            .I(N__73144));
    Sp12to4 I__17727 (
            .O(N__73182),
            .I(N__73137));
    Sp12to4 I__17726 (
            .O(N__73179),
            .I(N__73137));
    Sp12to4 I__17725 (
            .O(N__73176),
            .I(N__73137));
    LocalMux I__17724 (
            .O(N__73173),
            .I(N__73134));
    Span4Mux_h I__17723 (
            .O(N__73170),
            .I(N__73131));
    LocalMux I__17722 (
            .O(N__73167),
            .I(N__73124));
    LocalMux I__17721 (
            .O(N__73160),
            .I(N__73124));
    Sp12to4 I__17720 (
            .O(N__73157),
            .I(N__73124));
    InMux I__17719 (
            .O(N__73156),
            .I(N__73121));
    InMux I__17718 (
            .O(N__73155),
            .I(N__73118));
    InMux I__17717 (
            .O(N__73154),
            .I(N__73113));
    InMux I__17716 (
            .O(N__73153),
            .I(N__73113));
    LocalMux I__17715 (
            .O(N__73150),
            .I(N__73110));
    Sp12to4 I__17714 (
            .O(N__73147),
            .I(N__73103));
    Sp12to4 I__17713 (
            .O(N__73144),
            .I(N__73103));
    Span12Mux_v I__17712 (
            .O(N__73137),
            .I(N__73103));
    Span12Mux_h I__17711 (
            .O(N__73134),
            .I(N__73096));
    Sp12to4 I__17710 (
            .O(N__73131),
            .I(N__73096));
    Span12Mux_v I__17709 (
            .O(N__73124),
            .I(N__73096));
    LocalMux I__17708 (
            .O(N__73121),
            .I(rx_data_6));
    LocalMux I__17707 (
            .O(N__73118),
            .I(rx_data_6));
    LocalMux I__17706 (
            .O(N__73113),
            .I(rx_data_6));
    Odrv4 I__17705 (
            .O(N__73110),
            .I(rx_data_6));
    Odrv12 I__17704 (
            .O(N__73103),
            .I(rx_data_6));
    Odrv12 I__17703 (
            .O(N__73096),
            .I(rx_data_6));
    CascadeMux I__17702 (
            .O(N__73083),
            .I(N__73078));
    CascadeMux I__17701 (
            .O(N__73082),
            .I(N__73075));
    InMux I__17700 (
            .O(N__73081),
            .I(N__73072));
    InMux I__17699 (
            .O(N__73078),
            .I(N__73067));
    InMux I__17698 (
            .O(N__73075),
            .I(N__73067));
    LocalMux I__17697 (
            .O(N__73072),
            .I(N__73064));
    LocalMux I__17696 (
            .O(N__73067),
            .I(data_in_frame_22_1));
    Odrv4 I__17695 (
            .O(N__73064),
            .I(data_in_frame_22_1));
    CascadeMux I__17694 (
            .O(N__73059),
            .I(N__73056));
    InMux I__17693 (
            .O(N__73056),
            .I(N__73052));
    InMux I__17692 (
            .O(N__73055),
            .I(N__73049));
    LocalMux I__17691 (
            .O(N__73052),
            .I(N__73046));
    LocalMux I__17690 (
            .O(N__73049),
            .I(N__73043));
    Odrv4 I__17689 (
            .O(N__73046),
            .I(\c0.data_in_frame_20_2 ));
    Odrv4 I__17688 (
            .O(N__73043),
            .I(\c0.data_in_frame_20_2 ));
    CascadeMux I__17687 (
            .O(N__73038),
            .I(N__73035));
    InMux I__17686 (
            .O(N__73035),
            .I(N__73030));
    InMux I__17685 (
            .O(N__73034),
            .I(N__73027));
    InMux I__17684 (
            .O(N__73033),
            .I(N__73024));
    LocalMux I__17683 (
            .O(N__73030),
            .I(N__73021));
    LocalMux I__17682 (
            .O(N__73027),
            .I(N__73015));
    LocalMux I__17681 (
            .O(N__73024),
            .I(N__73015));
    Span4Mux_h I__17680 (
            .O(N__73021),
            .I(N__73012));
    InMux I__17679 (
            .O(N__73020),
            .I(N__73009));
    Span4Mux_h I__17678 (
            .O(N__73015),
            .I(N__73006));
    Span4Mux_v I__17677 (
            .O(N__73012),
            .I(N__73003));
    LocalMux I__17676 (
            .O(N__73009),
            .I(\c0.data_in_frame_23_5 ));
    Odrv4 I__17675 (
            .O(N__73006),
            .I(\c0.data_in_frame_23_5 ));
    Odrv4 I__17674 (
            .O(N__73003),
            .I(\c0.data_in_frame_23_5 ));
    CascadeMux I__17673 (
            .O(N__72996),
            .I(N__72993));
    InMux I__17672 (
            .O(N__72993),
            .I(N__72986));
    CascadeMux I__17671 (
            .O(N__72992),
            .I(N__72983));
    InMux I__17670 (
            .O(N__72991),
            .I(N__72974));
    InMux I__17669 (
            .O(N__72990),
            .I(N__72971));
    InMux I__17668 (
            .O(N__72989),
            .I(N__72968));
    LocalMux I__17667 (
            .O(N__72986),
            .I(N__72961));
    InMux I__17666 (
            .O(N__72983),
            .I(N__72956));
    InMux I__17665 (
            .O(N__72982),
            .I(N__72956));
    InMux I__17664 (
            .O(N__72981),
            .I(N__72949));
    InMux I__17663 (
            .O(N__72980),
            .I(N__72949));
    InMux I__17662 (
            .O(N__72979),
            .I(N__72949));
    CascadeMux I__17661 (
            .O(N__72978),
            .I(N__72946));
    CascadeMux I__17660 (
            .O(N__72977),
            .I(N__72943));
    LocalMux I__17659 (
            .O(N__72974),
            .I(N__72932));
    LocalMux I__17658 (
            .O(N__72971),
            .I(N__72929));
    LocalMux I__17657 (
            .O(N__72968),
            .I(N__72926));
    CascadeMux I__17656 (
            .O(N__72967),
            .I(N__72920));
    CascadeMux I__17655 (
            .O(N__72966),
            .I(N__72917));
    InMux I__17654 (
            .O(N__72965),
            .I(N__72912));
    InMux I__17653 (
            .O(N__72964),
            .I(N__72912));
    Span4Mux_h I__17652 (
            .O(N__72961),
            .I(N__72909));
    LocalMux I__17651 (
            .O(N__72956),
            .I(N__72906));
    LocalMux I__17650 (
            .O(N__72949),
            .I(N__72903));
    InMux I__17649 (
            .O(N__72946),
            .I(N__72900));
    InMux I__17648 (
            .O(N__72943),
            .I(N__72893));
    InMux I__17647 (
            .O(N__72942),
            .I(N__72893));
    InMux I__17646 (
            .O(N__72941),
            .I(N__72890));
    InMux I__17645 (
            .O(N__72940),
            .I(N__72887));
    InMux I__17644 (
            .O(N__72939),
            .I(N__72884));
    InMux I__17643 (
            .O(N__72938),
            .I(N__72881));
    InMux I__17642 (
            .O(N__72937),
            .I(N__72875));
    InMux I__17641 (
            .O(N__72936),
            .I(N__72875));
    InMux I__17640 (
            .O(N__72935),
            .I(N__72872));
    Span4Mux_v I__17639 (
            .O(N__72932),
            .I(N__72869));
    Span4Mux_h I__17638 (
            .O(N__72929),
            .I(N__72866));
    Span4Mux_h I__17637 (
            .O(N__72926),
            .I(N__72863));
    InMux I__17636 (
            .O(N__72925),
            .I(N__72857));
    InMux I__17635 (
            .O(N__72924),
            .I(N__72848));
    InMux I__17634 (
            .O(N__72923),
            .I(N__72848));
    InMux I__17633 (
            .O(N__72920),
            .I(N__72848));
    InMux I__17632 (
            .O(N__72917),
            .I(N__72848));
    LocalMux I__17631 (
            .O(N__72912),
            .I(N__72845));
    Span4Mux_h I__17630 (
            .O(N__72909),
            .I(N__72838));
    Span4Mux_h I__17629 (
            .O(N__72906),
            .I(N__72838));
    Span4Mux_h I__17628 (
            .O(N__72903),
            .I(N__72838));
    LocalMux I__17627 (
            .O(N__72900),
            .I(N__72835));
    InMux I__17626 (
            .O(N__72899),
            .I(N__72832));
    InMux I__17625 (
            .O(N__72898),
            .I(N__72829));
    LocalMux I__17624 (
            .O(N__72893),
            .I(N__72826));
    LocalMux I__17623 (
            .O(N__72890),
            .I(N__72821));
    LocalMux I__17622 (
            .O(N__72887),
            .I(N__72821));
    LocalMux I__17621 (
            .O(N__72884),
            .I(N__72816));
    LocalMux I__17620 (
            .O(N__72881),
            .I(N__72816));
    InMux I__17619 (
            .O(N__72880),
            .I(N__72813));
    LocalMux I__17618 (
            .O(N__72875),
            .I(N__72810));
    LocalMux I__17617 (
            .O(N__72872),
            .I(N__72805));
    Span4Mux_v I__17616 (
            .O(N__72869),
            .I(N__72805));
    Span4Mux_v I__17615 (
            .O(N__72866),
            .I(N__72800));
    Span4Mux_v I__17614 (
            .O(N__72863),
            .I(N__72800));
    InMux I__17613 (
            .O(N__72862),
            .I(N__72797));
    InMux I__17612 (
            .O(N__72861),
            .I(N__72792));
    InMux I__17611 (
            .O(N__72860),
            .I(N__72792));
    LocalMux I__17610 (
            .O(N__72857),
            .I(N__72789));
    LocalMux I__17609 (
            .O(N__72848),
            .I(N__72786));
    Span4Mux_h I__17608 (
            .O(N__72845),
            .I(N__72781));
    Span4Mux_v I__17607 (
            .O(N__72838),
            .I(N__72781));
    Span4Mux_v I__17606 (
            .O(N__72835),
            .I(N__72774));
    LocalMux I__17605 (
            .O(N__72832),
            .I(N__72774));
    LocalMux I__17604 (
            .O(N__72829),
            .I(N__72774));
    Span4Mux_h I__17603 (
            .O(N__72826),
            .I(N__72771));
    Span4Mux_v I__17602 (
            .O(N__72821),
            .I(N__72768));
    Span4Mux_v I__17601 (
            .O(N__72816),
            .I(N__72765));
    LocalMux I__17600 (
            .O(N__72813),
            .I(N__72762));
    Span4Mux_v I__17599 (
            .O(N__72810),
            .I(N__72759));
    Span4Mux_h I__17598 (
            .O(N__72805),
            .I(N__72754));
    Span4Mux_v I__17597 (
            .O(N__72800),
            .I(N__72754));
    LocalMux I__17596 (
            .O(N__72797),
            .I(N__72751));
    LocalMux I__17595 (
            .O(N__72792),
            .I(N__72748));
    Span4Mux_h I__17594 (
            .O(N__72789),
            .I(N__72745));
    Span4Mux_h I__17593 (
            .O(N__72786),
            .I(N__72740));
    Span4Mux_v I__17592 (
            .O(N__72781),
            .I(N__72740));
    Span4Mux_h I__17591 (
            .O(N__72774),
            .I(N__72737));
    Sp12to4 I__17590 (
            .O(N__72771),
            .I(N__72734));
    Sp12to4 I__17589 (
            .O(N__72768),
            .I(N__72729));
    Sp12to4 I__17588 (
            .O(N__72765),
            .I(N__72729));
    Span4Mux_h I__17587 (
            .O(N__72762),
            .I(N__72722));
    Span4Mux_h I__17586 (
            .O(N__72759),
            .I(N__72722));
    Span4Mux_v I__17585 (
            .O(N__72754),
            .I(N__72722));
    Span12Mux_h I__17584 (
            .O(N__72751),
            .I(N__72717));
    Span12Mux_h I__17583 (
            .O(N__72748),
            .I(N__72717));
    Span4Mux_h I__17582 (
            .O(N__72745),
            .I(N__72712));
    Span4Mux_v I__17581 (
            .O(N__72740),
            .I(N__72712));
    Sp12to4 I__17580 (
            .O(N__72737),
            .I(N__72705));
    Span12Mux_v I__17579 (
            .O(N__72734),
            .I(N__72705));
    Span12Mux_h I__17578 (
            .O(N__72729),
            .I(N__72705));
    Span4Mux_v I__17577 (
            .O(N__72722),
            .I(N__72702));
    Odrv12 I__17576 (
            .O(N__72717),
            .I(\c0.n9_adj_4563 ));
    Odrv4 I__17575 (
            .O(N__72712),
            .I(\c0.n9_adj_4563 ));
    Odrv12 I__17574 (
            .O(N__72705),
            .I(\c0.n9_adj_4563 ));
    Odrv4 I__17573 (
            .O(N__72702),
            .I(\c0.n9_adj_4563 ));
    CascadeMux I__17572 (
            .O(N__72693),
            .I(N__72690));
    InMux I__17571 (
            .O(N__72690),
            .I(N__72686));
    InMux I__17570 (
            .O(N__72689),
            .I(N__72683));
    LocalMux I__17569 (
            .O(N__72686),
            .I(N__72678));
    LocalMux I__17568 (
            .O(N__72683),
            .I(N__72675));
    CascadeMux I__17567 (
            .O(N__72682),
            .I(N__72672));
    InMux I__17566 (
            .O(N__72681),
            .I(N__72669));
    Span4Mux_h I__17565 (
            .O(N__72678),
            .I(N__72666));
    Span4Mux_h I__17564 (
            .O(N__72675),
            .I(N__72663));
    InMux I__17563 (
            .O(N__72672),
            .I(N__72660));
    LocalMux I__17562 (
            .O(N__72669),
            .I(N__72657));
    Span4Mux_h I__17561 (
            .O(N__72666),
            .I(N__72654));
    Span4Mux_h I__17560 (
            .O(N__72663),
            .I(N__72651));
    LocalMux I__17559 (
            .O(N__72660),
            .I(\c0.data_in_frame_16_7 ));
    Odrv12 I__17558 (
            .O(N__72657),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__17557 (
            .O(N__72654),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__17556 (
            .O(N__72651),
            .I(\c0.data_in_frame_16_7 ));
    InMux I__17555 (
            .O(N__72642),
            .I(N__72639));
    LocalMux I__17554 (
            .O(N__72639),
            .I(N__72635));
    InMux I__17553 (
            .O(N__72638),
            .I(N__72632));
    Span4Mux_v I__17552 (
            .O(N__72635),
            .I(N__72626));
    LocalMux I__17551 (
            .O(N__72632),
            .I(N__72626));
    InMux I__17550 (
            .O(N__72631),
            .I(N__72623));
    Span4Mux_v I__17549 (
            .O(N__72626),
            .I(N__72620));
    LocalMux I__17548 (
            .O(N__72623),
            .I(N__72617));
    Odrv4 I__17547 (
            .O(N__72620),
            .I(\c0.n22_adj_4244 ));
    Odrv4 I__17546 (
            .O(N__72617),
            .I(\c0.n22_adj_4244 ));
    InMux I__17545 (
            .O(N__72612),
            .I(N__72609));
    LocalMux I__17544 (
            .O(N__72609),
            .I(\c0.n24_adj_4618 ));
    CascadeMux I__17543 (
            .O(N__72606),
            .I(N__72603));
    InMux I__17542 (
            .O(N__72603),
            .I(N__72600));
    LocalMux I__17541 (
            .O(N__72600),
            .I(N__72597));
    Odrv4 I__17540 (
            .O(N__72597),
            .I(\c0.n14_adj_4619 ));
    CascadeMux I__17539 (
            .O(N__72594),
            .I(N__72591));
    InMux I__17538 (
            .O(N__72591),
            .I(N__72588));
    LocalMux I__17537 (
            .O(N__72588),
            .I(N__72582));
    InMux I__17536 (
            .O(N__72587),
            .I(N__72578));
    CascadeMux I__17535 (
            .O(N__72586),
            .I(N__72574));
    CascadeMux I__17534 (
            .O(N__72585),
            .I(N__72571));
    Span4Mux_v I__17533 (
            .O(N__72582),
            .I(N__72567));
    InMux I__17532 (
            .O(N__72581),
            .I(N__72564));
    LocalMux I__17531 (
            .O(N__72578),
            .I(N__72560));
    InMux I__17530 (
            .O(N__72577),
            .I(N__72556));
    InMux I__17529 (
            .O(N__72574),
            .I(N__72553));
    InMux I__17528 (
            .O(N__72571),
            .I(N__72550));
    InMux I__17527 (
            .O(N__72570),
            .I(N__72547));
    Span4Mux_v I__17526 (
            .O(N__72567),
            .I(N__72542));
    LocalMux I__17525 (
            .O(N__72564),
            .I(N__72542));
    InMux I__17524 (
            .O(N__72563),
            .I(N__72539));
    Span4Mux_v I__17523 (
            .O(N__72560),
            .I(N__72536));
    InMux I__17522 (
            .O(N__72559),
            .I(N__72533));
    LocalMux I__17521 (
            .O(N__72556),
            .I(N__72530));
    LocalMux I__17520 (
            .O(N__72553),
            .I(N__72521));
    LocalMux I__17519 (
            .O(N__72550),
            .I(N__72521));
    LocalMux I__17518 (
            .O(N__72547),
            .I(N__72521));
    Span4Mux_v I__17517 (
            .O(N__72542),
            .I(N__72518));
    LocalMux I__17516 (
            .O(N__72539),
            .I(N__72515));
    Span4Mux_v I__17515 (
            .O(N__72536),
            .I(N__72508));
    LocalMux I__17514 (
            .O(N__72533),
            .I(N__72508));
    Span4Mux_h I__17513 (
            .O(N__72530),
            .I(N__72508));
    InMux I__17512 (
            .O(N__72529),
            .I(N__72503));
    InMux I__17511 (
            .O(N__72528),
            .I(N__72503));
    Span4Mux_h I__17510 (
            .O(N__72521),
            .I(N__72500));
    Odrv4 I__17509 (
            .O(N__72518),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__17508 (
            .O(N__72515),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__17507 (
            .O(N__72508),
            .I(\c0.data_in_frame_2_1 ));
    LocalMux I__17506 (
            .O(N__72503),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__17505 (
            .O(N__72500),
            .I(\c0.data_in_frame_2_1 ));
    InMux I__17504 (
            .O(N__72489),
            .I(N__72486));
    LocalMux I__17503 (
            .O(N__72486),
            .I(\c0.n22288 ));
    CascadeMux I__17502 (
            .O(N__72483),
            .I(N__72479));
    CascadeMux I__17501 (
            .O(N__72482),
            .I(N__72476));
    InMux I__17500 (
            .O(N__72479),
            .I(N__72473));
    InMux I__17499 (
            .O(N__72476),
            .I(N__72469));
    LocalMux I__17498 (
            .O(N__72473),
            .I(N__72465));
    InMux I__17497 (
            .O(N__72472),
            .I(N__72460));
    LocalMux I__17496 (
            .O(N__72469),
            .I(N__72457));
    InMux I__17495 (
            .O(N__72468),
            .I(N__72454));
    Span4Mux_h I__17494 (
            .O(N__72465),
            .I(N__72451));
    CascadeMux I__17493 (
            .O(N__72464),
            .I(N__72448));
    InMux I__17492 (
            .O(N__72463),
            .I(N__72445));
    LocalMux I__17491 (
            .O(N__72460),
            .I(N__72442));
    Span4Mux_v I__17490 (
            .O(N__72457),
            .I(N__72439));
    LocalMux I__17489 (
            .O(N__72454),
            .I(N__72436));
    Span4Mux_h I__17488 (
            .O(N__72451),
            .I(N__72433));
    InMux I__17487 (
            .O(N__72448),
            .I(N__72430));
    LocalMux I__17486 (
            .O(N__72445),
            .I(\c0.data_in_frame_13_2 ));
    Odrv4 I__17485 (
            .O(N__72442),
            .I(\c0.data_in_frame_13_2 ));
    Odrv4 I__17484 (
            .O(N__72439),
            .I(\c0.data_in_frame_13_2 ));
    Odrv4 I__17483 (
            .O(N__72436),
            .I(\c0.data_in_frame_13_2 ));
    Odrv4 I__17482 (
            .O(N__72433),
            .I(\c0.data_in_frame_13_2 ));
    LocalMux I__17481 (
            .O(N__72430),
            .I(\c0.data_in_frame_13_2 ));
    CascadeMux I__17480 (
            .O(N__72417),
            .I(\c0.n22288_cascade_ ));
    CascadeMux I__17479 (
            .O(N__72414),
            .I(N__72410));
    InMux I__17478 (
            .O(N__72413),
            .I(N__72407));
    InMux I__17477 (
            .O(N__72410),
            .I(N__72404));
    LocalMux I__17476 (
            .O(N__72407),
            .I(N__72401));
    LocalMux I__17475 (
            .O(N__72404),
            .I(N__72398));
    Span4Mux_h I__17474 (
            .O(N__72401),
            .I(N__72393));
    Span4Mux_v I__17473 (
            .O(N__72398),
            .I(N__72390));
    InMux I__17472 (
            .O(N__72397),
            .I(N__72387));
    InMux I__17471 (
            .O(N__72396),
            .I(N__72384));
    Span4Mux_v I__17470 (
            .O(N__72393),
            .I(N__72377));
    Span4Mux_h I__17469 (
            .O(N__72390),
            .I(N__72377));
    LocalMux I__17468 (
            .O(N__72387),
            .I(N__72377));
    LocalMux I__17467 (
            .O(N__72384),
            .I(\c0.n5807 ));
    Odrv4 I__17466 (
            .O(N__72377),
            .I(\c0.n5807 ));
    InMux I__17465 (
            .O(N__72372),
            .I(N__72367));
    InMux I__17464 (
            .O(N__72371),
            .I(N__72361));
    InMux I__17463 (
            .O(N__72370),
            .I(N__72361));
    LocalMux I__17462 (
            .O(N__72367),
            .I(N__72357));
    InMux I__17461 (
            .O(N__72366),
            .I(N__72354));
    LocalMux I__17460 (
            .O(N__72361),
            .I(N__72351));
    InMux I__17459 (
            .O(N__72360),
            .I(N__72348));
    Span4Mux_v I__17458 (
            .O(N__72357),
            .I(N__72342));
    LocalMux I__17457 (
            .O(N__72354),
            .I(N__72342));
    Span4Mux_v I__17456 (
            .O(N__72351),
            .I(N__72337));
    LocalMux I__17455 (
            .O(N__72348),
            .I(N__72337));
    InMux I__17454 (
            .O(N__72347),
            .I(N__72334));
    Span4Mux_v I__17453 (
            .O(N__72342),
            .I(N__72329));
    Span4Mux_h I__17452 (
            .O(N__72337),
            .I(N__72329));
    LocalMux I__17451 (
            .O(N__72334),
            .I(N__72326));
    Odrv4 I__17450 (
            .O(N__72329),
            .I(\c0.n14160 ));
    Odrv12 I__17449 (
            .O(N__72326),
            .I(\c0.n14160 ));
    InMux I__17448 (
            .O(N__72321),
            .I(N__72315));
    InMux I__17447 (
            .O(N__72320),
            .I(N__72310));
    InMux I__17446 (
            .O(N__72319),
            .I(N__72310));
    InMux I__17445 (
            .O(N__72318),
            .I(N__72306));
    LocalMux I__17444 (
            .O(N__72315),
            .I(N__72303));
    LocalMux I__17443 (
            .O(N__72310),
            .I(N__72300));
    CascadeMux I__17442 (
            .O(N__72309),
            .I(N__72296));
    LocalMux I__17441 (
            .O(N__72306),
            .I(N__72293));
    Span4Mux_v I__17440 (
            .O(N__72303),
            .I(N__72288));
    Span4Mux_h I__17439 (
            .O(N__72300),
            .I(N__72288));
    InMux I__17438 (
            .O(N__72299),
            .I(N__72285));
    InMux I__17437 (
            .O(N__72296),
            .I(N__72280));
    Span4Mux_h I__17436 (
            .O(N__72293),
            .I(N__72277));
    Span4Mux_v I__17435 (
            .O(N__72288),
            .I(N__72274));
    LocalMux I__17434 (
            .O(N__72285),
            .I(N__72271));
    InMux I__17433 (
            .O(N__72284),
            .I(N__72268));
    InMux I__17432 (
            .O(N__72283),
            .I(N__72265));
    LocalMux I__17431 (
            .O(N__72280),
            .I(\c0.data_in_frame_8_3 ));
    Odrv4 I__17430 (
            .O(N__72277),
            .I(\c0.data_in_frame_8_3 ));
    Odrv4 I__17429 (
            .O(N__72274),
            .I(\c0.data_in_frame_8_3 ));
    Odrv12 I__17428 (
            .O(N__72271),
            .I(\c0.data_in_frame_8_3 ));
    LocalMux I__17427 (
            .O(N__72268),
            .I(\c0.data_in_frame_8_3 ));
    LocalMux I__17426 (
            .O(N__72265),
            .I(\c0.data_in_frame_8_3 ));
    InMux I__17425 (
            .O(N__72252),
            .I(N__72246));
    InMux I__17424 (
            .O(N__72251),
            .I(N__72246));
    LocalMux I__17423 (
            .O(N__72246),
            .I(N__72243));
    Span4Mux_v I__17422 (
            .O(N__72243),
            .I(N__72239));
    InMux I__17421 (
            .O(N__72242),
            .I(N__72234));
    Span4Mux_h I__17420 (
            .O(N__72239),
            .I(N__72231));
    InMux I__17419 (
            .O(N__72238),
            .I(N__72226));
    InMux I__17418 (
            .O(N__72237),
            .I(N__72226));
    LocalMux I__17417 (
            .O(N__72234),
            .I(\c0.data_in_frame_17_4 ));
    Odrv4 I__17416 (
            .O(N__72231),
            .I(\c0.data_in_frame_17_4 ));
    LocalMux I__17415 (
            .O(N__72226),
            .I(\c0.data_in_frame_17_4 ));
    InMux I__17414 (
            .O(N__72219),
            .I(N__72216));
    LocalMux I__17413 (
            .O(N__72216),
            .I(N__72211));
    CascadeMux I__17412 (
            .O(N__72215),
            .I(N__72207));
    CascadeMux I__17411 (
            .O(N__72214),
            .I(N__72203));
    Span4Mux_v I__17410 (
            .O(N__72211),
            .I(N__72200));
    InMux I__17409 (
            .O(N__72210),
            .I(N__72197));
    InMux I__17408 (
            .O(N__72207),
            .I(N__72192));
    InMux I__17407 (
            .O(N__72206),
            .I(N__72187));
    InMux I__17406 (
            .O(N__72203),
            .I(N__72187));
    Span4Mux_h I__17405 (
            .O(N__72200),
            .I(N__72182));
    LocalMux I__17404 (
            .O(N__72197),
            .I(N__72182));
    InMux I__17403 (
            .O(N__72196),
            .I(N__72179));
    InMux I__17402 (
            .O(N__72195),
            .I(N__72176));
    LocalMux I__17401 (
            .O(N__72192),
            .I(\c0.data_in_frame_13_3 ));
    LocalMux I__17400 (
            .O(N__72187),
            .I(\c0.data_in_frame_13_3 ));
    Odrv4 I__17399 (
            .O(N__72182),
            .I(\c0.data_in_frame_13_3 ));
    LocalMux I__17398 (
            .O(N__72179),
            .I(\c0.data_in_frame_13_3 ));
    LocalMux I__17397 (
            .O(N__72176),
            .I(\c0.data_in_frame_13_3 ));
    InMux I__17396 (
            .O(N__72165),
            .I(N__72162));
    LocalMux I__17395 (
            .O(N__72162),
            .I(N__72158));
    InMux I__17394 (
            .O(N__72161),
            .I(N__72155));
    Span4Mux_h I__17393 (
            .O(N__72158),
            .I(N__72149));
    LocalMux I__17392 (
            .O(N__72155),
            .I(N__72146));
    InMux I__17391 (
            .O(N__72154),
            .I(N__72143));
    InMux I__17390 (
            .O(N__72153),
            .I(N__72138));
    InMux I__17389 (
            .O(N__72152),
            .I(N__72138));
    Span4Mux_h I__17388 (
            .O(N__72149),
            .I(N__72135));
    Span12Mux_v I__17387 (
            .O(N__72146),
            .I(N__72130));
    LocalMux I__17386 (
            .O(N__72143),
            .I(N__72130));
    LocalMux I__17385 (
            .O(N__72138),
            .I(\c0.n22319 ));
    Odrv4 I__17384 (
            .O(N__72135),
            .I(\c0.n22319 ));
    Odrv12 I__17383 (
            .O(N__72130),
            .I(\c0.n22319 ));
    InMux I__17382 (
            .O(N__72123),
            .I(N__72120));
    LocalMux I__17381 (
            .O(N__72120),
            .I(N__72117));
    Span4Mux_h I__17380 (
            .O(N__72117),
            .I(N__72114));
    Odrv4 I__17379 (
            .O(N__72114),
            .I(\c0.n4_adj_4586 ));
    InMux I__17378 (
            .O(N__72111),
            .I(N__72107));
    CascadeMux I__17377 (
            .O(N__72110),
            .I(N__72104));
    LocalMux I__17376 (
            .O(N__72107),
            .I(N__72100));
    InMux I__17375 (
            .O(N__72104),
            .I(N__72095));
    InMux I__17374 (
            .O(N__72103),
            .I(N__72095));
    Odrv4 I__17373 (
            .O(N__72100),
            .I(\c0.data_in_frame_16_0 ));
    LocalMux I__17372 (
            .O(N__72095),
            .I(\c0.data_in_frame_16_0 ));
    InMux I__17371 (
            .O(N__72090),
            .I(N__72085));
    InMux I__17370 (
            .O(N__72089),
            .I(N__72082));
    CascadeMux I__17369 (
            .O(N__72088),
            .I(N__72079));
    LocalMux I__17368 (
            .O(N__72085),
            .I(N__72075));
    LocalMux I__17367 (
            .O(N__72082),
            .I(N__72072));
    InMux I__17366 (
            .O(N__72079),
            .I(N__72067));
    InMux I__17365 (
            .O(N__72078),
            .I(N__72067));
    Odrv12 I__17364 (
            .O(N__72075),
            .I(\c0.data_in_frame_13_6 ));
    Odrv4 I__17363 (
            .O(N__72072),
            .I(\c0.data_in_frame_13_6 ));
    LocalMux I__17362 (
            .O(N__72067),
            .I(\c0.data_in_frame_13_6 ));
    CascadeMux I__17361 (
            .O(N__72060),
            .I(N__72057));
    InMux I__17360 (
            .O(N__72057),
            .I(N__72054));
    LocalMux I__17359 (
            .O(N__72054),
            .I(N__72051));
    Span12Mux_s11_h I__17358 (
            .O(N__72051),
            .I(N__72046));
    InMux I__17357 (
            .O(N__72050),
            .I(N__72041));
    InMux I__17356 (
            .O(N__72049),
            .I(N__72041));
    Odrv12 I__17355 (
            .O(N__72046),
            .I(\c0.data_in_frame_18_1 ));
    LocalMux I__17354 (
            .O(N__72041),
            .I(\c0.data_in_frame_18_1 ));
    InMux I__17353 (
            .O(N__72036),
            .I(N__72033));
    LocalMux I__17352 (
            .O(N__72033),
            .I(N__72029));
    InMux I__17351 (
            .O(N__72032),
            .I(N__72026));
    Odrv4 I__17350 (
            .O(N__72029),
            .I(\c0.n14081 ));
    LocalMux I__17349 (
            .O(N__72026),
            .I(\c0.n14081 ));
    InMux I__17348 (
            .O(N__72021),
            .I(N__72018));
    LocalMux I__17347 (
            .O(N__72018),
            .I(N__72014));
    InMux I__17346 (
            .O(N__72017),
            .I(N__72011));
    Odrv12 I__17345 (
            .O(N__72014),
            .I(\c0.n10_adj_4250 ));
    LocalMux I__17344 (
            .O(N__72011),
            .I(\c0.n10_adj_4250 ));
    CascadeMux I__17343 (
            .O(N__72006),
            .I(N__72003));
    InMux I__17342 (
            .O(N__72003),
            .I(N__71998));
    InMux I__17341 (
            .O(N__72002),
            .I(N__71995));
    InMux I__17340 (
            .O(N__72001),
            .I(N__71992));
    LocalMux I__17339 (
            .O(N__71998),
            .I(N__71989));
    LocalMux I__17338 (
            .O(N__71995),
            .I(N__71981));
    LocalMux I__17337 (
            .O(N__71992),
            .I(N__71981));
    Span4Mux_v I__17336 (
            .O(N__71989),
            .I(N__71981));
    InMux I__17335 (
            .O(N__71988),
            .I(N__71978));
    Span4Mux_h I__17334 (
            .O(N__71981),
            .I(N__71975));
    LocalMux I__17333 (
            .O(N__71978),
            .I(\c0.data_in_frame_16_4 ));
    Odrv4 I__17332 (
            .O(N__71975),
            .I(\c0.data_in_frame_16_4 ));
    CascadeMux I__17331 (
            .O(N__71970),
            .I(N__71963));
    CascadeMux I__17330 (
            .O(N__71969),
            .I(N__71960));
    InMux I__17329 (
            .O(N__71968),
            .I(N__71954));
    CascadeMux I__17328 (
            .O(N__71967),
            .I(N__71950));
    CascadeMux I__17327 (
            .O(N__71966),
            .I(N__71947));
    InMux I__17326 (
            .O(N__71963),
            .I(N__71940));
    InMux I__17325 (
            .O(N__71960),
            .I(N__71931));
    InMux I__17324 (
            .O(N__71959),
            .I(N__71931));
    InMux I__17323 (
            .O(N__71958),
            .I(N__71928));
    InMux I__17322 (
            .O(N__71957),
            .I(N__71925));
    LocalMux I__17321 (
            .O(N__71954),
            .I(N__71922));
    InMux I__17320 (
            .O(N__71953),
            .I(N__71918));
    InMux I__17319 (
            .O(N__71950),
            .I(N__71910));
    InMux I__17318 (
            .O(N__71947),
            .I(N__71907));
    CascadeMux I__17317 (
            .O(N__71946),
            .I(N__71903));
    InMux I__17316 (
            .O(N__71945),
            .I(N__71897));
    InMux I__17315 (
            .O(N__71944),
            .I(N__71897));
    InMux I__17314 (
            .O(N__71943),
            .I(N__71894));
    LocalMux I__17313 (
            .O(N__71940),
            .I(N__71891));
    InMux I__17312 (
            .O(N__71939),
            .I(N__71888));
    CascadeMux I__17311 (
            .O(N__71938),
            .I(N__71884));
    InMux I__17310 (
            .O(N__71937),
            .I(N__71879));
    InMux I__17309 (
            .O(N__71936),
            .I(N__71879));
    LocalMux I__17308 (
            .O(N__71931),
            .I(N__71876));
    LocalMux I__17307 (
            .O(N__71928),
            .I(N__71872));
    LocalMux I__17306 (
            .O(N__71925),
            .I(N__71867));
    Span4Mux_h I__17305 (
            .O(N__71922),
            .I(N__71867));
    CascadeMux I__17304 (
            .O(N__71921),
            .I(N__71863));
    LocalMux I__17303 (
            .O(N__71918),
            .I(N__71860));
    InMux I__17302 (
            .O(N__71917),
            .I(N__71855));
    InMux I__17301 (
            .O(N__71916),
            .I(N__71855));
    InMux I__17300 (
            .O(N__71915),
            .I(N__71850));
    InMux I__17299 (
            .O(N__71914),
            .I(N__71850));
    InMux I__17298 (
            .O(N__71913),
            .I(N__71847));
    LocalMux I__17297 (
            .O(N__71910),
            .I(N__71842));
    LocalMux I__17296 (
            .O(N__71907),
            .I(N__71842));
    InMux I__17295 (
            .O(N__71906),
            .I(N__71837));
    InMux I__17294 (
            .O(N__71903),
            .I(N__71837));
    InMux I__17293 (
            .O(N__71902),
            .I(N__71834));
    LocalMux I__17292 (
            .O(N__71897),
            .I(N__71831));
    LocalMux I__17291 (
            .O(N__71894),
            .I(N__71828));
    Span4Mux_h I__17290 (
            .O(N__71891),
            .I(N__71825));
    LocalMux I__17289 (
            .O(N__71888),
            .I(N__71822));
    InMux I__17288 (
            .O(N__71887),
            .I(N__71817));
    InMux I__17287 (
            .O(N__71884),
            .I(N__71817));
    LocalMux I__17286 (
            .O(N__71879),
            .I(N__71811));
    Span4Mux_v I__17285 (
            .O(N__71876),
            .I(N__71811));
    InMux I__17284 (
            .O(N__71875),
            .I(N__71808));
    Span4Mux_h I__17283 (
            .O(N__71872),
            .I(N__71805));
    Sp12to4 I__17282 (
            .O(N__71867),
            .I(N__71802));
    InMux I__17281 (
            .O(N__71866),
            .I(N__71799));
    InMux I__17280 (
            .O(N__71863),
            .I(N__71796));
    Span4Mux_v I__17279 (
            .O(N__71860),
            .I(N__71793));
    LocalMux I__17278 (
            .O(N__71855),
            .I(N__71790));
    LocalMux I__17277 (
            .O(N__71850),
            .I(N__71787));
    LocalMux I__17276 (
            .O(N__71847),
            .I(N__71782));
    Span4Mux_h I__17275 (
            .O(N__71842),
            .I(N__71782));
    LocalMux I__17274 (
            .O(N__71837),
            .I(N__71778));
    LocalMux I__17273 (
            .O(N__71834),
            .I(N__71773));
    Span4Mux_v I__17272 (
            .O(N__71831),
            .I(N__71773));
    Span4Mux_h I__17271 (
            .O(N__71828),
            .I(N__71768));
    Span4Mux_v I__17270 (
            .O(N__71825),
            .I(N__71768));
    Span4Mux_h I__17269 (
            .O(N__71822),
            .I(N__71763));
    LocalMux I__17268 (
            .O(N__71817),
            .I(N__71763));
    InMux I__17267 (
            .O(N__71816),
            .I(N__71758));
    Span4Mux_v I__17266 (
            .O(N__71811),
            .I(N__71753));
    LocalMux I__17265 (
            .O(N__71808),
            .I(N__71753));
    Sp12to4 I__17264 (
            .O(N__71805),
            .I(N__71744));
    Span12Mux_v I__17263 (
            .O(N__71802),
            .I(N__71744));
    LocalMux I__17262 (
            .O(N__71799),
            .I(N__71744));
    LocalMux I__17261 (
            .O(N__71796),
            .I(N__71744));
    Span4Mux_v I__17260 (
            .O(N__71793),
            .I(N__71741));
    Span4Mux_h I__17259 (
            .O(N__71790),
            .I(N__71734));
    Span4Mux_v I__17258 (
            .O(N__71787),
            .I(N__71734));
    Span4Mux_v I__17257 (
            .O(N__71782),
            .I(N__71734));
    InMux I__17256 (
            .O(N__71781),
            .I(N__71731));
    Span4Mux_v I__17255 (
            .O(N__71778),
            .I(N__71726));
    Span4Mux_v I__17254 (
            .O(N__71773),
            .I(N__71726));
    Sp12to4 I__17253 (
            .O(N__71768),
            .I(N__71723));
    Sp12to4 I__17252 (
            .O(N__71763),
            .I(N__71720));
    InMux I__17251 (
            .O(N__71762),
            .I(N__71715));
    InMux I__17250 (
            .O(N__71761),
            .I(N__71715));
    LocalMux I__17249 (
            .O(N__71758),
            .I(N__71712));
    Span4Mux_h I__17248 (
            .O(N__71753),
            .I(N__71709));
    Span12Mux_v I__17247 (
            .O(N__71744),
            .I(N__71706));
    Span4Mux_h I__17246 (
            .O(N__71741),
            .I(N__71701));
    Span4Mux_v I__17245 (
            .O(N__71734),
            .I(N__71701));
    LocalMux I__17244 (
            .O(N__71731),
            .I(N__71692));
    Sp12to4 I__17243 (
            .O(N__71726),
            .I(N__71692));
    Span12Mux_v I__17242 (
            .O(N__71723),
            .I(N__71692));
    Span12Mux_v I__17241 (
            .O(N__71720),
            .I(N__71692));
    LocalMux I__17240 (
            .O(N__71715),
            .I(rx_data_4));
    Odrv4 I__17239 (
            .O(N__71712),
            .I(rx_data_4));
    Odrv4 I__17238 (
            .O(N__71709),
            .I(rx_data_4));
    Odrv12 I__17237 (
            .O(N__71706),
            .I(rx_data_4));
    Odrv4 I__17236 (
            .O(N__71701),
            .I(rx_data_4));
    Odrv12 I__17235 (
            .O(N__71692),
            .I(rx_data_4));
    CascadeMux I__17234 (
            .O(N__71679),
            .I(N__71676));
    InMux I__17233 (
            .O(N__71676),
            .I(N__71670));
    InMux I__17232 (
            .O(N__71675),
            .I(N__71667));
    InMux I__17231 (
            .O(N__71674),
            .I(N__71662));
    InMux I__17230 (
            .O(N__71673),
            .I(N__71662));
    LocalMux I__17229 (
            .O(N__71670),
            .I(N__71659));
    LocalMux I__17228 (
            .O(N__71667),
            .I(N__71656));
    LocalMux I__17227 (
            .O(N__71662),
            .I(N__71653));
    Odrv4 I__17226 (
            .O(N__71659),
            .I(\c0.data_in_frame_13_4 ));
    Odrv4 I__17225 (
            .O(N__71656),
            .I(\c0.data_in_frame_13_4 ));
    Odrv4 I__17224 (
            .O(N__71653),
            .I(\c0.data_in_frame_13_4 ));
    InMux I__17223 (
            .O(N__71646),
            .I(N__71642));
    InMux I__17222 (
            .O(N__71645),
            .I(N__71639));
    LocalMux I__17221 (
            .O(N__71642),
            .I(N__71636));
    LocalMux I__17220 (
            .O(N__71639),
            .I(N__71632));
    Span4Mux_v I__17219 (
            .O(N__71636),
            .I(N__71628));
    CascadeMux I__17218 (
            .O(N__71635),
            .I(N__71624));
    Span4Mux_v I__17217 (
            .O(N__71632),
            .I(N__71621));
    CascadeMux I__17216 (
            .O(N__71631),
            .I(N__71618));
    Span4Mux_h I__17215 (
            .O(N__71628),
            .I(N__71615));
    InMux I__17214 (
            .O(N__71627),
            .I(N__71612));
    InMux I__17213 (
            .O(N__71624),
            .I(N__71609));
    Span4Mux_h I__17212 (
            .O(N__71621),
            .I(N__71606));
    InMux I__17211 (
            .O(N__71618),
            .I(N__71603));
    Sp12to4 I__17210 (
            .O(N__71615),
            .I(N__71598));
    LocalMux I__17209 (
            .O(N__71612),
            .I(N__71598));
    LocalMux I__17208 (
            .O(N__71609),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__17207 (
            .O(N__71606),
            .I(\c0.data_in_frame_19_5 ));
    LocalMux I__17206 (
            .O(N__71603),
            .I(\c0.data_in_frame_19_5 ));
    Odrv12 I__17205 (
            .O(N__71598),
            .I(\c0.data_in_frame_19_5 ));
    InMux I__17204 (
            .O(N__71589),
            .I(N__71585));
    InMux I__17203 (
            .O(N__71588),
            .I(N__71582));
    LocalMux I__17202 (
            .O(N__71585),
            .I(N__71579));
    LocalMux I__17201 (
            .O(N__71582),
            .I(N__71576));
    Span4Mux_h I__17200 (
            .O(N__71579),
            .I(N__71573));
    Span4Mux_v I__17199 (
            .O(N__71576),
            .I(N__71569));
    Span4Mux_h I__17198 (
            .O(N__71573),
            .I(N__71566));
    InMux I__17197 (
            .O(N__71572),
            .I(N__71563));
    Span4Mux_v I__17196 (
            .O(N__71569),
            .I(N__71560));
    Odrv4 I__17195 (
            .O(N__71566),
            .I(\c0.FRAME_MATCHER_i_18 ));
    LocalMux I__17194 (
            .O(N__71563),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__17193 (
            .O(N__71560),
            .I(\c0.FRAME_MATCHER_i_18 ));
    InMux I__17192 (
            .O(N__71553),
            .I(N__71549));
    InMux I__17191 (
            .O(N__71552),
            .I(N__71546));
    LocalMux I__17190 (
            .O(N__71549),
            .I(N__71539));
    LocalMux I__17189 (
            .O(N__71546),
            .I(N__71533));
    InMux I__17188 (
            .O(N__71545),
            .I(N__71530));
    InMux I__17187 (
            .O(N__71544),
            .I(N__71526));
    InMux I__17186 (
            .O(N__71543),
            .I(N__71523));
    InMux I__17185 (
            .O(N__71542),
            .I(N__71520));
    Span4Mux_h I__17184 (
            .O(N__71539),
            .I(N__71516));
    InMux I__17183 (
            .O(N__71538),
            .I(N__71513));
    InMux I__17182 (
            .O(N__71537),
            .I(N__71510));
    InMux I__17181 (
            .O(N__71536),
            .I(N__71507));
    Span4Mux_v I__17180 (
            .O(N__71533),
            .I(N__71499));
    LocalMux I__17179 (
            .O(N__71530),
            .I(N__71499));
    InMux I__17178 (
            .O(N__71529),
            .I(N__71496));
    LocalMux I__17177 (
            .O(N__71526),
            .I(N__71493));
    LocalMux I__17176 (
            .O(N__71523),
            .I(N__71490));
    LocalMux I__17175 (
            .O(N__71520),
            .I(N__71487));
    InMux I__17174 (
            .O(N__71519),
            .I(N__71484));
    Span4Mux_v I__17173 (
            .O(N__71516),
            .I(N__71477));
    LocalMux I__17172 (
            .O(N__71513),
            .I(N__71477));
    LocalMux I__17171 (
            .O(N__71510),
            .I(N__71474));
    LocalMux I__17170 (
            .O(N__71507),
            .I(N__71468));
    InMux I__17169 (
            .O(N__71506),
            .I(N__71465));
    InMux I__17168 (
            .O(N__71505),
            .I(N__71462));
    InMux I__17167 (
            .O(N__71504),
            .I(N__71459));
    Span4Mux_h I__17166 (
            .O(N__71499),
            .I(N__71451));
    LocalMux I__17165 (
            .O(N__71496),
            .I(N__71448));
    Span4Mux_h I__17164 (
            .O(N__71493),
            .I(N__71445));
    Span4Mux_v I__17163 (
            .O(N__71490),
            .I(N__71442));
    Span4Mux_v I__17162 (
            .O(N__71487),
            .I(N__71437));
    LocalMux I__17161 (
            .O(N__71484),
            .I(N__71437));
    InMux I__17160 (
            .O(N__71483),
            .I(N__71432));
    InMux I__17159 (
            .O(N__71482),
            .I(N__71432));
    Span4Mux_v I__17158 (
            .O(N__71477),
            .I(N__71429));
    Span4Mux_v I__17157 (
            .O(N__71474),
            .I(N__71425));
    InMux I__17156 (
            .O(N__71473),
            .I(N__71418));
    InMux I__17155 (
            .O(N__71472),
            .I(N__71418));
    InMux I__17154 (
            .O(N__71471),
            .I(N__71418));
    Span4Mux_h I__17153 (
            .O(N__71468),
            .I(N__71409));
    LocalMux I__17152 (
            .O(N__71465),
            .I(N__71409));
    LocalMux I__17151 (
            .O(N__71462),
            .I(N__71409));
    LocalMux I__17150 (
            .O(N__71459),
            .I(N__71409));
    InMux I__17149 (
            .O(N__71458),
            .I(N__71406));
    InMux I__17148 (
            .O(N__71457),
            .I(N__71403));
    InMux I__17147 (
            .O(N__71456),
            .I(N__71398));
    InMux I__17146 (
            .O(N__71455),
            .I(N__71398));
    InMux I__17145 (
            .O(N__71454),
            .I(N__71395));
    Sp12to4 I__17144 (
            .O(N__71451),
            .I(N__71391));
    Span12Mux_s11_h I__17143 (
            .O(N__71448),
            .I(N__71388));
    Span4Mux_h I__17142 (
            .O(N__71445),
            .I(N__71379));
    Span4Mux_h I__17141 (
            .O(N__71442),
            .I(N__71379));
    Span4Mux_v I__17140 (
            .O(N__71437),
            .I(N__71379));
    LocalMux I__17139 (
            .O(N__71432),
            .I(N__71379));
    Span4Mux_v I__17138 (
            .O(N__71429),
            .I(N__71376));
    InMux I__17137 (
            .O(N__71428),
            .I(N__71373));
    Span4Mux_v I__17136 (
            .O(N__71425),
            .I(N__71369));
    LocalMux I__17135 (
            .O(N__71418),
            .I(N__71366));
    Span4Mux_v I__17134 (
            .O(N__71409),
            .I(N__71355));
    LocalMux I__17133 (
            .O(N__71406),
            .I(N__71355));
    LocalMux I__17132 (
            .O(N__71403),
            .I(N__71355));
    LocalMux I__17131 (
            .O(N__71398),
            .I(N__71355));
    LocalMux I__17130 (
            .O(N__71395),
            .I(N__71355));
    InMux I__17129 (
            .O(N__71394),
            .I(N__71352));
    Span12Mux_v I__17128 (
            .O(N__71391),
            .I(N__71344));
    Span12Mux_v I__17127 (
            .O(N__71388),
            .I(N__71341));
    Span4Mux_v I__17126 (
            .O(N__71379),
            .I(N__71338));
    Span4Mux_v I__17125 (
            .O(N__71376),
            .I(N__71333));
    LocalMux I__17124 (
            .O(N__71373),
            .I(N__71333));
    InMux I__17123 (
            .O(N__71372),
            .I(N__71330));
    Span4Mux_h I__17122 (
            .O(N__71369),
            .I(N__71321));
    Span4Mux_v I__17121 (
            .O(N__71366),
            .I(N__71321));
    Span4Mux_v I__17120 (
            .O(N__71355),
            .I(N__71321));
    LocalMux I__17119 (
            .O(N__71352),
            .I(N__71321));
    InMux I__17118 (
            .O(N__71351),
            .I(N__71310));
    InMux I__17117 (
            .O(N__71350),
            .I(N__71310));
    InMux I__17116 (
            .O(N__71349),
            .I(N__71310));
    InMux I__17115 (
            .O(N__71348),
            .I(N__71310));
    InMux I__17114 (
            .O(N__71347),
            .I(N__71310));
    Odrv12 I__17113 (
            .O(N__71344),
            .I(\c0.n2119 ));
    Odrv12 I__17112 (
            .O(N__71341),
            .I(\c0.n2119 ));
    Odrv4 I__17111 (
            .O(N__71338),
            .I(\c0.n2119 ));
    Odrv4 I__17110 (
            .O(N__71333),
            .I(\c0.n2119 ));
    LocalMux I__17109 (
            .O(N__71330),
            .I(\c0.n2119 ));
    Odrv4 I__17108 (
            .O(N__71321),
            .I(\c0.n2119 ));
    LocalMux I__17107 (
            .O(N__71310),
            .I(\c0.n2119 ));
    SRMux I__17106 (
            .O(N__71295),
            .I(N__71292));
    LocalMux I__17105 (
            .O(N__71292),
            .I(N__71289));
    Span4Mux_v I__17104 (
            .O(N__71289),
            .I(N__71286));
    Span4Mux_h I__17103 (
            .O(N__71286),
            .I(N__71283));
    Odrv4 I__17102 (
            .O(N__71283),
            .I(\c0.n3_adj_4400 ));
    CascadeMux I__17101 (
            .O(N__71280),
            .I(N__71277));
    InMux I__17100 (
            .O(N__71277),
            .I(N__71274));
    LocalMux I__17099 (
            .O(N__71274),
            .I(N__71271));
    Span4Mux_v I__17098 (
            .O(N__71271),
            .I(N__71265));
    InMux I__17097 (
            .O(N__71270),
            .I(N__71260));
    InMux I__17096 (
            .O(N__71269),
            .I(N__71260));
    InMux I__17095 (
            .O(N__71268),
            .I(N__71257));
    Span4Mux_h I__17094 (
            .O(N__71265),
            .I(N__71254));
    LocalMux I__17093 (
            .O(N__71260),
            .I(\c0.data_in_frame_17_6 ));
    LocalMux I__17092 (
            .O(N__71257),
            .I(\c0.data_in_frame_17_6 ));
    Odrv4 I__17091 (
            .O(N__71254),
            .I(\c0.data_in_frame_17_6 ));
    InMux I__17090 (
            .O(N__71247),
            .I(N__71243));
    CascadeMux I__17089 (
            .O(N__71246),
            .I(N__71239));
    LocalMux I__17088 (
            .O(N__71243),
            .I(N__71236));
    InMux I__17087 (
            .O(N__71242),
            .I(N__71233));
    InMux I__17086 (
            .O(N__71239),
            .I(N__71230));
    Span4Mux_v I__17085 (
            .O(N__71236),
            .I(N__71225));
    LocalMux I__17084 (
            .O(N__71233),
            .I(N__71225));
    LocalMux I__17083 (
            .O(N__71230),
            .I(\c0.data_in_frame_15_5 ));
    Odrv4 I__17082 (
            .O(N__71225),
            .I(\c0.data_in_frame_15_5 ));
    CascadeMux I__17081 (
            .O(N__71220),
            .I(N__71216));
    InMux I__17080 (
            .O(N__71219),
            .I(N__71213));
    InMux I__17079 (
            .O(N__71216),
            .I(N__71210));
    LocalMux I__17078 (
            .O(N__71213),
            .I(N__71206));
    LocalMux I__17077 (
            .O(N__71210),
            .I(N__71203));
    InMux I__17076 (
            .O(N__71209),
            .I(N__71200));
    Span4Mux_h I__17075 (
            .O(N__71206),
            .I(N__71197));
    Span4Mux_v I__17074 (
            .O(N__71203),
            .I(N__71192));
    LocalMux I__17073 (
            .O(N__71200),
            .I(N__71192));
    Odrv4 I__17072 (
            .O(N__71197),
            .I(\c0.n31_adj_4701 ));
    Odrv4 I__17071 (
            .O(N__71192),
            .I(\c0.n31_adj_4701 ));
    CascadeMux I__17070 (
            .O(N__71187),
            .I(N__71184));
    InMux I__17069 (
            .O(N__71184),
            .I(N__71181));
    LocalMux I__17068 (
            .O(N__71181),
            .I(N__71178));
    Span4Mux_h I__17067 (
            .O(N__71178),
            .I(N__71172));
    InMux I__17066 (
            .O(N__71177),
            .I(N__71169));
    CascadeMux I__17065 (
            .O(N__71176),
            .I(N__71166));
    InMux I__17064 (
            .O(N__71175),
            .I(N__71163));
    Span4Mux_h I__17063 (
            .O(N__71172),
            .I(N__71158));
    LocalMux I__17062 (
            .O(N__71169),
            .I(N__71158));
    InMux I__17061 (
            .O(N__71166),
            .I(N__71155));
    LocalMux I__17060 (
            .O(N__71163),
            .I(\c0.n13474 ));
    Odrv4 I__17059 (
            .O(N__71158),
            .I(\c0.n13474 ));
    LocalMux I__17058 (
            .O(N__71155),
            .I(\c0.n13474 ));
    CascadeMux I__17057 (
            .O(N__71148),
            .I(N__71145));
    InMux I__17056 (
            .O(N__71145),
            .I(N__71142));
    LocalMux I__17055 (
            .O(N__71142),
            .I(N__71139));
    Span4Mux_h I__17054 (
            .O(N__71139),
            .I(N__71136));
    Odrv4 I__17053 (
            .O(N__71136),
            .I(\c0.n22650 ));
    InMux I__17052 (
            .O(N__71133),
            .I(N__71130));
    LocalMux I__17051 (
            .O(N__71130),
            .I(N__71127));
    Span4Mux_h I__17050 (
            .O(N__71127),
            .I(N__71123));
    InMux I__17049 (
            .O(N__71126),
            .I(N__71120));
    Span4Mux_h I__17048 (
            .O(N__71123),
            .I(N__71110));
    LocalMux I__17047 (
            .O(N__71120),
            .I(N__71107));
    InMux I__17046 (
            .O(N__71119),
            .I(N__71104));
    InMux I__17045 (
            .O(N__71118),
            .I(N__71101));
    InMux I__17044 (
            .O(N__71117),
            .I(N__71096));
    InMux I__17043 (
            .O(N__71116),
            .I(N__71088));
    InMux I__17042 (
            .O(N__71115),
            .I(N__71081));
    InMux I__17041 (
            .O(N__71114),
            .I(N__71081));
    InMux I__17040 (
            .O(N__71113),
            .I(N__71081));
    Span4Mux_v I__17039 (
            .O(N__71110),
            .I(N__71068));
    Span4Mux_h I__17038 (
            .O(N__71107),
            .I(N__71068));
    LocalMux I__17037 (
            .O(N__71104),
            .I(N__71068));
    LocalMux I__17036 (
            .O(N__71101),
            .I(N__71068));
    InMux I__17035 (
            .O(N__71100),
            .I(N__71065));
    InMux I__17034 (
            .O(N__71099),
            .I(N__71062));
    LocalMux I__17033 (
            .O(N__71096),
            .I(N__71059));
    InMux I__17032 (
            .O(N__71095),
            .I(N__71054));
    InMux I__17031 (
            .O(N__71094),
            .I(N__71054));
    InMux I__17030 (
            .O(N__71093),
            .I(N__71051));
    InMux I__17029 (
            .O(N__71092),
            .I(N__71046));
    InMux I__17028 (
            .O(N__71091),
            .I(N__71046));
    LocalMux I__17027 (
            .O(N__71088),
            .I(N__71041));
    LocalMux I__17026 (
            .O(N__71081),
            .I(N__71041));
    InMux I__17025 (
            .O(N__71080),
            .I(N__71036));
    InMux I__17024 (
            .O(N__71079),
            .I(N__71036));
    CascadeMux I__17023 (
            .O(N__71078),
            .I(N__71033));
    InMux I__17022 (
            .O(N__71077),
            .I(N__71027));
    Span4Mux_v I__17021 (
            .O(N__71068),
            .I(N__71024));
    LocalMux I__17020 (
            .O(N__71065),
            .I(N__71019));
    LocalMux I__17019 (
            .O(N__71062),
            .I(N__71019));
    Span4Mux_v I__17018 (
            .O(N__71059),
            .I(N__71016));
    LocalMux I__17017 (
            .O(N__71054),
            .I(N__71005));
    LocalMux I__17016 (
            .O(N__71051),
            .I(N__71005));
    LocalMux I__17015 (
            .O(N__71046),
            .I(N__71005));
    Span4Mux_v I__17014 (
            .O(N__71041),
            .I(N__71005));
    LocalMux I__17013 (
            .O(N__71036),
            .I(N__71005));
    InMux I__17012 (
            .O(N__71033),
            .I(N__71002));
    InMux I__17011 (
            .O(N__71032),
            .I(N__70999));
    InMux I__17010 (
            .O(N__71031),
            .I(N__70994));
    InMux I__17009 (
            .O(N__71030),
            .I(N__70994));
    LocalMux I__17008 (
            .O(N__71027),
            .I(N__70989));
    Span4Mux_h I__17007 (
            .O(N__71024),
            .I(N__70989));
    Span4Mux_v I__17006 (
            .O(N__71019),
            .I(N__70982));
    Span4Mux_h I__17005 (
            .O(N__71016),
            .I(N__70982));
    Span4Mux_v I__17004 (
            .O(N__71005),
            .I(N__70982));
    LocalMux I__17003 (
            .O(N__71002),
            .I(data_in_frame_1_7));
    LocalMux I__17002 (
            .O(N__70999),
            .I(data_in_frame_1_7));
    LocalMux I__17001 (
            .O(N__70994),
            .I(data_in_frame_1_7));
    Odrv4 I__17000 (
            .O(N__70989),
            .I(data_in_frame_1_7));
    Odrv4 I__16999 (
            .O(N__70982),
            .I(data_in_frame_1_7));
    CascadeMux I__16998 (
            .O(N__70971),
            .I(N__70968));
    InMux I__16997 (
            .O(N__70968),
            .I(N__70965));
    LocalMux I__16996 (
            .O(N__70965),
            .I(N__70962));
    Odrv4 I__16995 (
            .O(N__70962),
            .I(\c0.n30_adj_4747 ));
    InMux I__16994 (
            .O(N__70959),
            .I(N__70955));
    InMux I__16993 (
            .O(N__70958),
            .I(N__70952));
    LocalMux I__16992 (
            .O(N__70955),
            .I(N__70949));
    LocalMux I__16991 (
            .O(N__70952),
            .I(N__70946));
    Span4Mux_v I__16990 (
            .O(N__70949),
            .I(N__70943));
    Span4Mux_v I__16989 (
            .O(N__70946),
            .I(N__70940));
    Span4Mux_v I__16988 (
            .O(N__70943),
            .I(N__70937));
    Odrv4 I__16987 (
            .O(N__70940),
            .I(\c0.n6_adj_4632 ));
    Odrv4 I__16986 (
            .O(N__70937),
            .I(\c0.n6_adj_4632 ));
    InMux I__16985 (
            .O(N__70932),
            .I(N__70929));
    LocalMux I__16984 (
            .O(N__70929),
            .I(\c0.n5_adj_4631 ));
    InMux I__16983 (
            .O(N__70926),
            .I(N__70923));
    LocalMux I__16982 (
            .O(N__70923),
            .I(N__70919));
    InMux I__16981 (
            .O(N__70922),
            .I(N__70916));
    Span4Mux_h I__16980 (
            .O(N__70919),
            .I(N__70910));
    LocalMux I__16979 (
            .O(N__70916),
            .I(N__70910));
    InMux I__16978 (
            .O(N__70915),
            .I(N__70907));
    Span4Mux_v I__16977 (
            .O(N__70910),
            .I(N__70902));
    LocalMux I__16976 (
            .O(N__70907),
            .I(N__70902));
    Odrv4 I__16975 (
            .O(N__70902),
            .I(\c0.n23343 ));
    InMux I__16974 (
            .O(N__70899),
            .I(N__70896));
    LocalMux I__16973 (
            .O(N__70896),
            .I(N__70893));
    Sp12to4 I__16972 (
            .O(N__70893),
            .I(N__70890));
    Odrv12 I__16971 (
            .O(N__70890),
            .I(\c0.n25_adj_4633 ));
    InMux I__16970 (
            .O(N__70887),
            .I(N__70880));
    InMux I__16969 (
            .O(N__70886),
            .I(N__70880));
    InMux I__16968 (
            .O(N__70885),
            .I(N__70877));
    LocalMux I__16967 (
            .O(N__70880),
            .I(N__70873));
    LocalMux I__16966 (
            .O(N__70877),
            .I(N__70870));
    InMux I__16965 (
            .O(N__70876),
            .I(N__70867));
    Span4Mux_h I__16964 (
            .O(N__70873),
            .I(N__70864));
    Span12Mux_v I__16963 (
            .O(N__70870),
            .I(N__70861));
    LocalMux I__16962 (
            .O(N__70867),
            .I(\c0.data_in_frame_9_3 ));
    Odrv4 I__16961 (
            .O(N__70864),
            .I(\c0.data_in_frame_9_3 ));
    Odrv12 I__16960 (
            .O(N__70861),
            .I(\c0.data_in_frame_9_3 ));
    InMux I__16959 (
            .O(N__70854),
            .I(N__70851));
    LocalMux I__16958 (
            .O(N__70851),
            .I(N__70844));
    InMux I__16957 (
            .O(N__70850),
            .I(N__70841));
    InMux I__16956 (
            .O(N__70849),
            .I(N__70838));
    InMux I__16955 (
            .O(N__70848),
            .I(N__70835));
    InMux I__16954 (
            .O(N__70847),
            .I(N__70832));
    Span4Mux_h I__16953 (
            .O(N__70844),
            .I(N__70827));
    LocalMux I__16952 (
            .O(N__70841),
            .I(N__70827));
    LocalMux I__16951 (
            .O(N__70838),
            .I(\c0.data_in_frame_11_2 ));
    LocalMux I__16950 (
            .O(N__70835),
            .I(\c0.data_in_frame_11_2 ));
    LocalMux I__16949 (
            .O(N__70832),
            .I(\c0.data_in_frame_11_2 ));
    Odrv4 I__16948 (
            .O(N__70827),
            .I(\c0.data_in_frame_11_2 ));
    CascadeMux I__16947 (
            .O(N__70818),
            .I(N__70815));
    InMux I__16946 (
            .O(N__70815),
            .I(N__70812));
    LocalMux I__16945 (
            .O(N__70812),
            .I(N__70809));
    Span4Mux_v I__16944 (
            .O(N__70809),
            .I(N__70805));
    CascadeMux I__16943 (
            .O(N__70808),
            .I(N__70802));
    Span4Mux_h I__16942 (
            .O(N__70805),
            .I(N__70799));
    InMux I__16941 (
            .O(N__70802),
            .I(N__70796));
    Span4Mux_h I__16940 (
            .O(N__70799),
            .I(N__70793));
    LocalMux I__16939 (
            .O(N__70796),
            .I(\c0.data_in_frame_28_1 ));
    Odrv4 I__16938 (
            .O(N__70793),
            .I(\c0.data_in_frame_28_1 ));
    InMux I__16937 (
            .O(N__70788),
            .I(N__70784));
    CascadeMux I__16936 (
            .O(N__70787),
            .I(N__70781));
    LocalMux I__16935 (
            .O(N__70784),
            .I(N__70778));
    InMux I__16934 (
            .O(N__70781),
            .I(N__70775));
    Span4Mux_v I__16933 (
            .O(N__70778),
            .I(N__70771));
    LocalMux I__16932 (
            .O(N__70775),
            .I(N__70768));
    CascadeMux I__16931 (
            .O(N__70774),
            .I(N__70765));
    Span4Mux_h I__16930 (
            .O(N__70771),
            .I(N__70760));
    Span4Mux_v I__16929 (
            .O(N__70768),
            .I(N__70760));
    InMux I__16928 (
            .O(N__70765),
            .I(N__70757));
    Span4Mux_h I__16927 (
            .O(N__70760),
            .I(N__70754));
    LocalMux I__16926 (
            .O(N__70757),
            .I(\c0.data_in_frame_11_4 ));
    Odrv4 I__16925 (
            .O(N__70754),
            .I(\c0.data_in_frame_11_4 ));
    InMux I__16924 (
            .O(N__70749),
            .I(N__70746));
    LocalMux I__16923 (
            .O(N__70746),
            .I(N__70743));
    Span4Mux_h I__16922 (
            .O(N__70743),
            .I(N__70738));
    InMux I__16921 (
            .O(N__70742),
            .I(N__70735));
    CascadeMux I__16920 (
            .O(N__70741),
            .I(N__70732));
    Span4Mux_v I__16919 (
            .O(N__70738),
            .I(N__70727));
    LocalMux I__16918 (
            .O(N__70735),
            .I(N__70727));
    InMux I__16917 (
            .O(N__70732),
            .I(N__70724));
    Span4Mux_h I__16916 (
            .O(N__70727),
            .I(N__70721));
    LocalMux I__16915 (
            .O(N__70724),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__16914 (
            .O(N__70721),
            .I(\c0.data_in_frame_7_2 ));
    CascadeMux I__16913 (
            .O(N__70716),
            .I(N__70712));
    InMux I__16912 (
            .O(N__70715),
            .I(N__70709));
    InMux I__16911 (
            .O(N__70712),
            .I(N__70706));
    LocalMux I__16910 (
            .O(N__70709),
            .I(\c0.n9_adj_4220 ));
    LocalMux I__16909 (
            .O(N__70706),
            .I(\c0.n9_adj_4220 ));
    InMux I__16908 (
            .O(N__70701),
            .I(N__70698));
    LocalMux I__16907 (
            .O(N__70698),
            .I(N__70695));
    Span4Mux_v I__16906 (
            .O(N__70695),
            .I(N__70691));
    InMux I__16905 (
            .O(N__70694),
            .I(N__70688));
    Odrv4 I__16904 (
            .O(N__70691),
            .I(\c0.n7_adj_4226 ));
    LocalMux I__16903 (
            .O(N__70688),
            .I(\c0.n7_adj_4226 ));
    InMux I__16902 (
            .O(N__70683),
            .I(N__70680));
    LocalMux I__16901 (
            .O(N__70680),
            .I(\c0.n27_adj_4748 ));
    CascadeMux I__16900 (
            .O(N__70677),
            .I(N__70674));
    InMux I__16899 (
            .O(N__70674),
            .I(N__70669));
    CascadeMux I__16898 (
            .O(N__70673),
            .I(N__70666));
    InMux I__16897 (
            .O(N__70672),
            .I(N__70663));
    LocalMux I__16896 (
            .O(N__70669),
            .I(N__70660));
    InMux I__16895 (
            .O(N__70666),
            .I(N__70655));
    LocalMux I__16894 (
            .O(N__70663),
            .I(N__70652));
    Span4Mux_v I__16893 (
            .O(N__70660),
            .I(N__70649));
    InMux I__16892 (
            .O(N__70659),
            .I(N__70646));
    CascadeMux I__16891 (
            .O(N__70658),
            .I(N__70642));
    LocalMux I__16890 (
            .O(N__70655),
            .I(N__70637));
    Span4Mux_v I__16889 (
            .O(N__70652),
            .I(N__70637));
    Span4Mux_h I__16888 (
            .O(N__70649),
            .I(N__70632));
    LocalMux I__16887 (
            .O(N__70646),
            .I(N__70632));
    InMux I__16886 (
            .O(N__70645),
            .I(N__70627));
    InMux I__16885 (
            .O(N__70642),
            .I(N__70627));
    Odrv4 I__16884 (
            .O(N__70637),
            .I(\c0.data_in_frame_11_3 ));
    Odrv4 I__16883 (
            .O(N__70632),
            .I(\c0.data_in_frame_11_3 ));
    LocalMux I__16882 (
            .O(N__70627),
            .I(\c0.data_in_frame_11_3 ));
    InMux I__16881 (
            .O(N__70620),
            .I(N__70615));
    InMux I__16880 (
            .O(N__70619),
            .I(N__70612));
    InMux I__16879 (
            .O(N__70618),
            .I(N__70609));
    LocalMux I__16878 (
            .O(N__70615),
            .I(\c0.data_in_frame_9_0 ));
    LocalMux I__16877 (
            .O(N__70612),
            .I(\c0.data_in_frame_9_0 ));
    LocalMux I__16876 (
            .O(N__70609),
            .I(\c0.data_in_frame_9_0 ));
    InMux I__16875 (
            .O(N__70602),
            .I(N__70599));
    LocalMux I__16874 (
            .O(N__70599),
            .I(N__70595));
    CascadeMux I__16873 (
            .O(N__70598),
            .I(N__70592));
    Span4Mux_h I__16872 (
            .O(N__70595),
            .I(N__70588));
    InMux I__16871 (
            .O(N__70592),
            .I(N__70585));
    InMux I__16870 (
            .O(N__70591),
            .I(N__70582));
    Odrv4 I__16869 (
            .O(N__70588),
            .I(\c0.n4 ));
    LocalMux I__16868 (
            .O(N__70585),
            .I(\c0.n4 ));
    LocalMux I__16867 (
            .O(N__70582),
            .I(\c0.n4 ));
    InMux I__16866 (
            .O(N__70575),
            .I(N__70572));
    LocalMux I__16865 (
            .O(N__70572),
            .I(N__70568));
    CascadeMux I__16864 (
            .O(N__70571),
            .I(N__70565));
    Span4Mux_h I__16863 (
            .O(N__70568),
            .I(N__70562));
    InMux I__16862 (
            .O(N__70565),
            .I(N__70559));
    Span4Mux_v I__16861 (
            .O(N__70562),
            .I(N__70556));
    LocalMux I__16860 (
            .O(N__70559),
            .I(\c0.data_in_frame_28_3 ));
    Odrv4 I__16859 (
            .O(N__70556),
            .I(\c0.data_in_frame_28_3 ));
    InMux I__16858 (
            .O(N__70551),
            .I(N__70545));
    CascadeMux I__16857 (
            .O(N__70550),
            .I(N__70542));
    InMux I__16856 (
            .O(N__70549),
            .I(N__70537));
    InMux I__16855 (
            .O(N__70548),
            .I(N__70537));
    LocalMux I__16854 (
            .O(N__70545),
            .I(N__70534));
    InMux I__16853 (
            .O(N__70542),
            .I(N__70531));
    LocalMux I__16852 (
            .O(N__70537),
            .I(N__70528));
    Span4Mux_h I__16851 (
            .O(N__70534),
            .I(N__70524));
    LocalMux I__16850 (
            .O(N__70531),
            .I(N__70519));
    Span4Mux_v I__16849 (
            .O(N__70528),
            .I(N__70519));
    InMux I__16848 (
            .O(N__70527),
            .I(N__70516));
    Span4Mux_h I__16847 (
            .O(N__70524),
            .I(N__70513));
    Odrv4 I__16846 (
            .O(N__70519),
            .I(\c0.data_in_frame_12_3 ));
    LocalMux I__16845 (
            .O(N__70516),
            .I(\c0.data_in_frame_12_3 ));
    Odrv4 I__16844 (
            .O(N__70513),
            .I(\c0.data_in_frame_12_3 ));
    CascadeMux I__16843 (
            .O(N__70506),
            .I(N__70502));
    InMux I__16842 (
            .O(N__70505),
            .I(N__70499));
    InMux I__16841 (
            .O(N__70502),
            .I(N__70495));
    LocalMux I__16840 (
            .O(N__70499),
            .I(N__70492));
    InMux I__16839 (
            .O(N__70498),
            .I(N__70489));
    LocalMux I__16838 (
            .O(N__70495),
            .I(\c0.data_in_frame_15_6 ));
    Odrv4 I__16837 (
            .O(N__70492),
            .I(\c0.data_in_frame_15_6 ));
    LocalMux I__16836 (
            .O(N__70489),
            .I(\c0.data_in_frame_15_6 ));
    CascadeMux I__16835 (
            .O(N__70482),
            .I(N__70479));
    InMux I__16834 (
            .O(N__70479),
            .I(N__70476));
    LocalMux I__16833 (
            .O(N__70476),
            .I(N__70473));
    Span4Mux_h I__16832 (
            .O(N__70473),
            .I(N__70470));
    Span4Mux_h I__16831 (
            .O(N__70470),
            .I(N__70466));
    InMux I__16830 (
            .O(N__70469),
            .I(N__70463));
    Odrv4 I__16829 (
            .O(N__70466),
            .I(\c0.n22379 ));
    LocalMux I__16828 (
            .O(N__70463),
            .I(\c0.n22379 ));
    CascadeMux I__16827 (
            .O(N__70458),
            .I(N__70455));
    InMux I__16826 (
            .O(N__70455),
            .I(N__70452));
    LocalMux I__16825 (
            .O(N__70452),
            .I(\c0.n6_adj_4559 ));
    CascadeMux I__16824 (
            .O(N__70449),
            .I(N__70446));
    InMux I__16823 (
            .O(N__70446),
            .I(N__70440));
    InMux I__16822 (
            .O(N__70445),
            .I(N__70432));
    InMux I__16821 (
            .O(N__70444),
            .I(N__70432));
    InMux I__16820 (
            .O(N__70443),
            .I(N__70432));
    LocalMux I__16819 (
            .O(N__70440),
            .I(N__70429));
    InMux I__16818 (
            .O(N__70439),
            .I(N__70426));
    LocalMux I__16817 (
            .O(N__70432),
            .I(N__70422));
    Span4Mux_v I__16816 (
            .O(N__70429),
            .I(N__70417));
    LocalMux I__16815 (
            .O(N__70426),
            .I(N__70417));
    InMux I__16814 (
            .O(N__70425),
            .I(N__70414));
    Span4Mux_h I__16813 (
            .O(N__70422),
            .I(N__70411));
    Span4Mux_h I__16812 (
            .O(N__70417),
            .I(N__70408));
    LocalMux I__16811 (
            .O(N__70414),
            .I(\c0.data_in_frame_9_5 ));
    Odrv4 I__16810 (
            .O(N__70411),
            .I(\c0.data_in_frame_9_5 ));
    Odrv4 I__16809 (
            .O(N__70408),
            .I(\c0.data_in_frame_9_5 ));
    InMux I__16808 (
            .O(N__70401),
            .I(N__70397));
    InMux I__16807 (
            .O(N__70400),
            .I(N__70394));
    LocalMux I__16806 (
            .O(N__70397),
            .I(N__70391));
    LocalMux I__16805 (
            .O(N__70394),
            .I(N__70388));
    Span4Mux_v I__16804 (
            .O(N__70391),
            .I(N__70384));
    Span12Mux_h I__16803 (
            .O(N__70388),
            .I(N__70381));
    InMux I__16802 (
            .O(N__70387),
            .I(N__70378));
    Sp12to4 I__16801 (
            .O(N__70384),
            .I(N__70373));
    Span12Mux_v I__16800 (
            .O(N__70381),
            .I(N__70373));
    LocalMux I__16799 (
            .O(N__70378),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv12 I__16798 (
            .O(N__70373),
            .I(\c0.FRAME_MATCHER_i_13 ));
    SRMux I__16797 (
            .O(N__70368),
            .I(N__70365));
    LocalMux I__16796 (
            .O(N__70365),
            .I(N__70362));
    Span4Mux_v I__16795 (
            .O(N__70362),
            .I(N__70359));
    Span4Mux_h I__16794 (
            .O(N__70359),
            .I(N__70356));
    Odrv4 I__16793 (
            .O(N__70356),
            .I(\c0.n3_adj_4410 ));
    InMux I__16792 (
            .O(N__70353),
            .I(N__70349));
    InMux I__16791 (
            .O(N__70352),
            .I(N__70344));
    LocalMux I__16790 (
            .O(N__70349),
            .I(N__70341));
    InMux I__16789 (
            .O(N__70348),
            .I(N__70338));
    CascadeMux I__16788 (
            .O(N__70347),
            .I(N__70335));
    LocalMux I__16787 (
            .O(N__70344),
            .I(N__70332));
    Span4Mux_h I__16786 (
            .O(N__70341),
            .I(N__70329));
    LocalMux I__16785 (
            .O(N__70338),
            .I(N__70325));
    InMux I__16784 (
            .O(N__70335),
            .I(N__70322));
    Span4Mux_h I__16783 (
            .O(N__70332),
            .I(N__70319));
    Span4Mux_h I__16782 (
            .O(N__70329),
            .I(N__70316));
    InMux I__16781 (
            .O(N__70328),
            .I(N__70313));
    Span4Mux_h I__16780 (
            .O(N__70325),
            .I(N__70310));
    LocalMux I__16779 (
            .O(N__70322),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__16778 (
            .O(N__70319),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__16777 (
            .O(N__70316),
            .I(\c0.data_in_frame_7_4 ));
    LocalMux I__16776 (
            .O(N__70313),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__16775 (
            .O(N__70310),
            .I(\c0.data_in_frame_7_4 ));
    InMux I__16774 (
            .O(N__70299),
            .I(N__70294));
    InMux I__16773 (
            .O(N__70298),
            .I(N__70291));
    InMux I__16772 (
            .O(N__70297),
            .I(N__70288));
    LocalMux I__16771 (
            .O(N__70294),
            .I(N__70285));
    LocalMux I__16770 (
            .O(N__70291),
            .I(N__70281));
    LocalMux I__16769 (
            .O(N__70288),
            .I(N__70278));
    Span4Mux_v I__16768 (
            .O(N__70285),
            .I(N__70274));
    InMux I__16767 (
            .O(N__70284),
            .I(N__70271));
    Span4Mux_v I__16766 (
            .O(N__70281),
            .I(N__70268));
    Span4Mux_v I__16765 (
            .O(N__70278),
            .I(N__70265));
    CascadeMux I__16764 (
            .O(N__70277),
            .I(N__70261));
    Span4Mux_h I__16763 (
            .O(N__70274),
            .I(N__70258));
    LocalMux I__16762 (
            .O(N__70271),
            .I(N__70253));
    Span4Mux_h I__16761 (
            .O(N__70268),
            .I(N__70253));
    Span4Mux_h I__16760 (
            .O(N__70265),
            .I(N__70250));
    InMux I__16759 (
            .O(N__70264),
            .I(N__70247));
    InMux I__16758 (
            .O(N__70261),
            .I(N__70244));
    Odrv4 I__16757 (
            .O(N__70258),
            .I(data_in_frame_5_1));
    Odrv4 I__16756 (
            .O(N__70253),
            .I(data_in_frame_5_1));
    Odrv4 I__16755 (
            .O(N__70250),
            .I(data_in_frame_5_1));
    LocalMux I__16754 (
            .O(N__70247),
            .I(data_in_frame_5_1));
    LocalMux I__16753 (
            .O(N__70244),
            .I(data_in_frame_5_1));
    InMux I__16752 (
            .O(N__70233),
            .I(N__70230));
    LocalMux I__16751 (
            .O(N__70230),
            .I(N__70226));
    InMux I__16750 (
            .O(N__70229),
            .I(N__70222));
    Span4Mux_h I__16749 (
            .O(N__70226),
            .I(N__70219));
    InMux I__16748 (
            .O(N__70225),
            .I(N__70216));
    LocalMux I__16747 (
            .O(N__70222),
            .I(N__70212));
    Span4Mux_h I__16746 (
            .O(N__70219),
            .I(N__70209));
    LocalMux I__16745 (
            .O(N__70216),
            .I(N__70206));
    InMux I__16744 (
            .O(N__70215),
            .I(N__70203));
    Odrv12 I__16743 (
            .O(N__70212),
            .I(\c0.n40_adj_4288 ));
    Odrv4 I__16742 (
            .O(N__70209),
            .I(\c0.n40_adj_4288 ));
    Odrv4 I__16741 (
            .O(N__70206),
            .I(\c0.n40_adj_4288 ));
    LocalMux I__16740 (
            .O(N__70203),
            .I(\c0.n40_adj_4288 ));
    InMux I__16739 (
            .O(N__70194),
            .I(N__70188));
    InMux I__16738 (
            .O(N__70193),
            .I(N__70188));
    LocalMux I__16737 (
            .O(N__70188),
            .I(N__70183));
    InMux I__16736 (
            .O(N__70187),
            .I(N__70180));
    CascadeMux I__16735 (
            .O(N__70186),
            .I(N__70175));
    Span4Mux_v I__16734 (
            .O(N__70183),
            .I(N__70159));
    LocalMux I__16733 (
            .O(N__70180),
            .I(N__70159));
    InMux I__16732 (
            .O(N__70179),
            .I(N__70156));
    InMux I__16731 (
            .O(N__70178),
            .I(N__70131));
    InMux I__16730 (
            .O(N__70175),
            .I(N__70131));
    InMux I__16729 (
            .O(N__70174),
            .I(N__70131));
    InMux I__16728 (
            .O(N__70173),
            .I(N__70128));
    InMux I__16727 (
            .O(N__70172),
            .I(N__70121));
    InMux I__16726 (
            .O(N__70171),
            .I(N__70121));
    InMux I__16725 (
            .O(N__70170),
            .I(N__70121));
    InMux I__16724 (
            .O(N__70169),
            .I(N__70116));
    InMux I__16723 (
            .O(N__70168),
            .I(N__70116));
    InMux I__16722 (
            .O(N__70167),
            .I(N__70107));
    InMux I__16721 (
            .O(N__70166),
            .I(N__70107));
    InMux I__16720 (
            .O(N__70165),
            .I(N__70107));
    InMux I__16719 (
            .O(N__70164),
            .I(N__70107));
    Span4Mux_h I__16718 (
            .O(N__70159),
            .I(N__70102));
    LocalMux I__16717 (
            .O(N__70156),
            .I(N__70102));
    InMux I__16716 (
            .O(N__70155),
            .I(N__70097));
    InMux I__16715 (
            .O(N__70154),
            .I(N__70097));
    InMux I__16714 (
            .O(N__70153),
            .I(N__70094));
    InMux I__16713 (
            .O(N__70152),
            .I(N__70091));
    InMux I__16712 (
            .O(N__70151),
            .I(N__70088));
    CascadeMux I__16711 (
            .O(N__70150),
            .I(N__70084));
    InMux I__16710 (
            .O(N__70149),
            .I(N__70075));
    InMux I__16709 (
            .O(N__70148),
            .I(N__70070));
    InMux I__16708 (
            .O(N__70147),
            .I(N__70070));
    InMux I__16707 (
            .O(N__70146),
            .I(N__70063));
    InMux I__16706 (
            .O(N__70145),
            .I(N__70063));
    InMux I__16705 (
            .O(N__70144),
            .I(N__70063));
    InMux I__16704 (
            .O(N__70143),
            .I(N__70058));
    InMux I__16703 (
            .O(N__70142),
            .I(N__70058));
    InMux I__16702 (
            .O(N__70141),
            .I(N__70055));
    InMux I__16701 (
            .O(N__70140),
            .I(N__70048));
    InMux I__16700 (
            .O(N__70139),
            .I(N__70048));
    InMux I__16699 (
            .O(N__70138),
            .I(N__70048));
    LocalMux I__16698 (
            .O(N__70131),
            .I(N__70045));
    LocalMux I__16697 (
            .O(N__70128),
            .I(N__70038));
    LocalMux I__16696 (
            .O(N__70121),
            .I(N__70038));
    LocalMux I__16695 (
            .O(N__70116),
            .I(N__70038));
    LocalMux I__16694 (
            .O(N__70107),
            .I(N__70031));
    Span4Mux_h I__16693 (
            .O(N__70102),
            .I(N__70031));
    LocalMux I__16692 (
            .O(N__70097),
            .I(N__70031));
    LocalMux I__16691 (
            .O(N__70094),
            .I(N__70024));
    LocalMux I__16690 (
            .O(N__70091),
            .I(N__70024));
    LocalMux I__16689 (
            .O(N__70088),
            .I(N__70024));
    CascadeMux I__16688 (
            .O(N__70087),
            .I(N__70019));
    InMux I__16687 (
            .O(N__70084),
            .I(N__70005));
    InMux I__16686 (
            .O(N__70083),
            .I(N__70005));
    InMux I__16685 (
            .O(N__70082),
            .I(N__70005));
    InMux I__16684 (
            .O(N__70081),
            .I(N__70005));
    InMux I__16683 (
            .O(N__70080),
            .I(N__69998));
    InMux I__16682 (
            .O(N__70079),
            .I(N__69998));
    InMux I__16681 (
            .O(N__70078),
            .I(N__69998));
    LocalMux I__16680 (
            .O(N__70075),
            .I(N__69993));
    LocalMux I__16679 (
            .O(N__70070),
            .I(N__69993));
    LocalMux I__16678 (
            .O(N__70063),
            .I(N__69988));
    LocalMux I__16677 (
            .O(N__70058),
            .I(N__69988));
    LocalMux I__16676 (
            .O(N__70055),
            .I(N__69979));
    LocalMux I__16675 (
            .O(N__70048),
            .I(N__69979));
    Span4Mux_h I__16674 (
            .O(N__70045),
            .I(N__69979));
    Span4Mux_v I__16673 (
            .O(N__70038),
            .I(N__69979));
    Span4Mux_v I__16672 (
            .O(N__70031),
            .I(N__69974));
    Span4Mux_v I__16671 (
            .O(N__70024),
            .I(N__69974));
    InMux I__16670 (
            .O(N__70023),
            .I(N__69969));
    InMux I__16669 (
            .O(N__70022),
            .I(N__69969));
    InMux I__16668 (
            .O(N__70019),
            .I(N__69966));
    InMux I__16667 (
            .O(N__70018),
            .I(N__69963));
    InMux I__16666 (
            .O(N__70017),
            .I(N__69954));
    InMux I__16665 (
            .O(N__70016),
            .I(N__69954));
    InMux I__16664 (
            .O(N__70015),
            .I(N__69954));
    InMux I__16663 (
            .O(N__70014),
            .I(N__69954));
    LocalMux I__16662 (
            .O(N__70005),
            .I(N__69951));
    LocalMux I__16661 (
            .O(N__69998),
            .I(N__69946));
    Span4Mux_v I__16660 (
            .O(N__69993),
            .I(N__69946));
    Span4Mux_h I__16659 (
            .O(N__69988),
            .I(N__69941));
    Span4Mux_h I__16658 (
            .O(N__69979),
            .I(N__69941));
    Sp12to4 I__16657 (
            .O(N__69974),
            .I(N__69938));
    LocalMux I__16656 (
            .O(N__69969),
            .I(N__69935));
    LocalMux I__16655 (
            .O(N__69966),
            .I(N__69928));
    LocalMux I__16654 (
            .O(N__69963),
            .I(N__69928));
    LocalMux I__16653 (
            .O(N__69954),
            .I(N__69928));
    Span4Mux_v I__16652 (
            .O(N__69951),
            .I(N__69925));
    Span4Mux_h I__16651 (
            .O(N__69946),
            .I(N__69920));
    Span4Mux_v I__16650 (
            .O(N__69941),
            .I(N__69920));
    Span12Mux_h I__16649 (
            .O(N__69938),
            .I(N__69917));
    Span4Mux_v I__16648 (
            .O(N__69935),
            .I(N__69912));
    Span4Mux_h I__16647 (
            .O(N__69928),
            .I(N__69912));
    Odrv4 I__16646 (
            .O(N__69925),
            .I(\c0.n22120 ));
    Odrv4 I__16645 (
            .O(N__69920),
            .I(\c0.n22120 ));
    Odrv12 I__16644 (
            .O(N__69917),
            .I(\c0.n22120 ));
    Odrv4 I__16643 (
            .O(N__69912),
            .I(\c0.n22120 ));
    InMux I__16642 (
            .O(N__69903),
            .I(N__69899));
    CascadeMux I__16641 (
            .O(N__69902),
            .I(N__69895));
    LocalMux I__16640 (
            .O(N__69899),
            .I(N__69891));
    InMux I__16639 (
            .O(N__69898),
            .I(N__69888));
    InMux I__16638 (
            .O(N__69895),
            .I(N__69885));
    InMux I__16637 (
            .O(N__69894),
            .I(N__69881));
    Span4Mux_h I__16636 (
            .O(N__69891),
            .I(N__69878));
    LocalMux I__16635 (
            .O(N__69888),
            .I(N__69873));
    LocalMux I__16634 (
            .O(N__69885),
            .I(N__69873));
    CascadeMux I__16633 (
            .O(N__69884),
            .I(N__69870));
    LocalMux I__16632 (
            .O(N__69881),
            .I(N__69867));
    Span4Mux_v I__16631 (
            .O(N__69878),
            .I(N__69862));
    Span4Mux_v I__16630 (
            .O(N__69873),
            .I(N__69862));
    InMux I__16629 (
            .O(N__69870),
            .I(N__69857));
    Span4Mux_v I__16628 (
            .O(N__69867),
            .I(N__69852));
    Span4Mux_h I__16627 (
            .O(N__69862),
            .I(N__69852));
    InMux I__16626 (
            .O(N__69861),
            .I(N__69847));
    InMux I__16625 (
            .O(N__69860),
            .I(N__69847));
    LocalMux I__16624 (
            .O(N__69857),
            .I(N__69844));
    Odrv4 I__16623 (
            .O(N__69852),
            .I(\c0.data_in_frame_7_3 ));
    LocalMux I__16622 (
            .O(N__69847),
            .I(\c0.data_in_frame_7_3 ));
    Odrv4 I__16621 (
            .O(N__69844),
            .I(\c0.data_in_frame_7_3 ));
    InMux I__16620 (
            .O(N__69837),
            .I(N__69834));
    LocalMux I__16619 (
            .O(N__69834),
            .I(N__69829));
    CascadeMux I__16618 (
            .O(N__69833),
            .I(N__69826));
    CascadeMux I__16617 (
            .O(N__69832),
            .I(N__69822));
    Span4Mux_h I__16616 (
            .O(N__69829),
            .I(N__69819));
    InMux I__16615 (
            .O(N__69826),
            .I(N__69814));
    InMux I__16614 (
            .O(N__69825),
            .I(N__69814));
    InMux I__16613 (
            .O(N__69822),
            .I(N__69811));
    Odrv4 I__16612 (
            .O(N__69819),
            .I(\c0.data_in_frame_12_0 ));
    LocalMux I__16611 (
            .O(N__69814),
            .I(\c0.data_in_frame_12_0 ));
    LocalMux I__16610 (
            .O(N__69811),
            .I(\c0.data_in_frame_12_0 ));
    InMux I__16609 (
            .O(N__69804),
            .I(N__69801));
    LocalMux I__16608 (
            .O(N__69801),
            .I(N__69797));
    InMux I__16607 (
            .O(N__69800),
            .I(N__69794));
    Span4Mux_v I__16606 (
            .O(N__69797),
            .I(N__69789));
    LocalMux I__16605 (
            .O(N__69794),
            .I(N__69785));
    InMux I__16604 (
            .O(N__69793),
            .I(N__69780));
    InMux I__16603 (
            .O(N__69792),
            .I(N__69780));
    Span4Mux_h I__16602 (
            .O(N__69789),
            .I(N__69777));
    InMux I__16601 (
            .O(N__69788),
            .I(N__69774));
    Odrv12 I__16600 (
            .O(N__69785),
            .I(\c0.data_in_frame_12_1 ));
    LocalMux I__16599 (
            .O(N__69780),
            .I(\c0.data_in_frame_12_1 ));
    Odrv4 I__16598 (
            .O(N__69777),
            .I(\c0.data_in_frame_12_1 ));
    LocalMux I__16597 (
            .O(N__69774),
            .I(\c0.data_in_frame_12_1 ));
    InMux I__16596 (
            .O(N__69765),
            .I(N__69762));
    LocalMux I__16595 (
            .O(N__69762),
            .I(N__69755));
    InMux I__16594 (
            .O(N__69761),
            .I(N__69752));
    InMux I__16593 (
            .O(N__69760),
            .I(N__69747));
    InMux I__16592 (
            .O(N__69759),
            .I(N__69747));
    InMux I__16591 (
            .O(N__69758),
            .I(N__69744));
    Span4Mux_h I__16590 (
            .O(N__69755),
            .I(N__69741));
    LocalMux I__16589 (
            .O(N__69752),
            .I(N__69738));
    LocalMux I__16588 (
            .O(N__69747),
            .I(N__69735));
    LocalMux I__16587 (
            .O(N__69744),
            .I(N__69732));
    Span4Mux_h I__16586 (
            .O(N__69741),
            .I(N__69729));
    Span4Mux_v I__16585 (
            .O(N__69738),
            .I(N__69725));
    Span4Mux_v I__16584 (
            .O(N__69735),
            .I(N__69720));
    Span4Mux_h I__16583 (
            .O(N__69732),
            .I(N__69720));
    Span4Mux_v I__16582 (
            .O(N__69729),
            .I(N__69717));
    InMux I__16581 (
            .O(N__69728),
            .I(N__69714));
    Span4Mux_h I__16580 (
            .O(N__69725),
            .I(N__69709));
    Span4Mux_v I__16579 (
            .O(N__69720),
            .I(N__69709));
    Odrv4 I__16578 (
            .O(N__69717),
            .I(\c0.n39 ));
    LocalMux I__16577 (
            .O(N__69714),
            .I(\c0.n39 ));
    Odrv4 I__16576 (
            .O(N__69709),
            .I(\c0.n39 ));
    InMux I__16575 (
            .O(N__69702),
            .I(N__69697));
    InMux I__16574 (
            .O(N__69701),
            .I(N__69694));
    InMux I__16573 (
            .O(N__69700),
            .I(N__69690));
    LocalMux I__16572 (
            .O(N__69697),
            .I(N__69687));
    LocalMux I__16571 (
            .O(N__69694),
            .I(N__69684));
    InMux I__16570 (
            .O(N__69693),
            .I(N__69681));
    LocalMux I__16569 (
            .O(N__69690),
            .I(N__69672));
    Span4Mux_h I__16568 (
            .O(N__69687),
            .I(N__69672));
    Span4Mux_v I__16567 (
            .O(N__69684),
            .I(N__69672));
    LocalMux I__16566 (
            .O(N__69681),
            .I(N__69672));
    Odrv4 I__16565 (
            .O(N__69672),
            .I(\c0.n61 ));
    CascadeMux I__16564 (
            .O(N__69669),
            .I(N__69666));
    InMux I__16563 (
            .O(N__69666),
            .I(N__69663));
    LocalMux I__16562 (
            .O(N__69663),
            .I(N__69660));
    Span4Mux_v I__16561 (
            .O(N__69660),
            .I(N__69657));
    Span4Mux_h I__16560 (
            .O(N__69657),
            .I(N__69654));
    Span4Mux_h I__16559 (
            .O(N__69654),
            .I(N__69651));
    Odrv4 I__16558 (
            .O(N__69651),
            .I(\c0.n13253 ));
    CascadeMux I__16557 (
            .O(N__69648),
            .I(\c0.n13253_cascade_ ));
    CascadeMux I__16556 (
            .O(N__69645),
            .I(N__69641));
    InMux I__16555 (
            .O(N__69644),
            .I(N__69637));
    InMux I__16554 (
            .O(N__69641),
            .I(N__69634));
    CascadeMux I__16553 (
            .O(N__69640),
            .I(N__69631));
    LocalMux I__16552 (
            .O(N__69637),
            .I(N__69627));
    LocalMux I__16551 (
            .O(N__69634),
            .I(N__69624));
    InMux I__16550 (
            .O(N__69631),
            .I(N__69619));
    InMux I__16549 (
            .O(N__69630),
            .I(N__69619));
    Span4Mux_h I__16548 (
            .O(N__69627),
            .I(N__69616));
    Odrv4 I__16547 (
            .O(N__69624),
            .I(\c0.n22518 ));
    LocalMux I__16546 (
            .O(N__69619),
            .I(\c0.n22518 ));
    Odrv4 I__16545 (
            .O(N__69616),
            .I(\c0.n22518 ));
    InMux I__16544 (
            .O(N__69609),
            .I(N__69605));
    InMux I__16543 (
            .O(N__69608),
            .I(N__69602));
    LocalMux I__16542 (
            .O(N__69605),
            .I(N__69599));
    LocalMux I__16541 (
            .O(N__69602),
            .I(N__69596));
    Span4Mux_v I__16540 (
            .O(N__69599),
            .I(N__69593));
    Sp12to4 I__16539 (
            .O(N__69596),
            .I(N__69590));
    Odrv4 I__16538 (
            .O(N__69593),
            .I(\c0.n22828 ));
    Odrv12 I__16537 (
            .O(N__69590),
            .I(\c0.n22828 ));
    InMux I__16536 (
            .O(N__69585),
            .I(N__69577));
    InMux I__16535 (
            .O(N__69584),
            .I(N__69574));
    InMux I__16534 (
            .O(N__69583),
            .I(N__69567));
    InMux I__16533 (
            .O(N__69582),
            .I(N__69567));
    InMux I__16532 (
            .O(N__69581),
            .I(N__69567));
    InMux I__16531 (
            .O(N__69580),
            .I(N__69564));
    LocalMux I__16530 (
            .O(N__69577),
            .I(N__69561));
    LocalMux I__16529 (
            .O(N__69574),
            .I(N__69558));
    LocalMux I__16528 (
            .O(N__69567),
            .I(N__69554));
    LocalMux I__16527 (
            .O(N__69564),
            .I(N__69551));
    Span4Mux_h I__16526 (
            .O(N__69561),
            .I(N__69543));
    Span4Mux_h I__16525 (
            .O(N__69558),
            .I(N__69540));
    InMux I__16524 (
            .O(N__69557),
            .I(N__69537));
    Span4Mux_v I__16523 (
            .O(N__69554),
            .I(N__69532));
    Span4Mux_h I__16522 (
            .O(N__69551),
            .I(N__69532));
    InMux I__16521 (
            .O(N__69550),
            .I(N__69525));
    InMux I__16520 (
            .O(N__69549),
            .I(N__69525));
    InMux I__16519 (
            .O(N__69548),
            .I(N__69525));
    InMux I__16518 (
            .O(N__69547),
            .I(N__69522));
    InMux I__16517 (
            .O(N__69546),
            .I(N__69519));
    Odrv4 I__16516 (
            .O(N__69543),
            .I(\c0.data_in_frame_0_0 ));
    Odrv4 I__16515 (
            .O(N__69540),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__16514 (
            .O(N__69537),
            .I(\c0.data_in_frame_0_0 ));
    Odrv4 I__16513 (
            .O(N__69532),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__16512 (
            .O(N__69525),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__16511 (
            .O(N__69522),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__16510 (
            .O(N__69519),
            .I(\c0.data_in_frame_0_0 ));
    CascadeMux I__16509 (
            .O(N__69504),
            .I(N__69501));
    InMux I__16508 (
            .O(N__69501),
            .I(N__69495));
    InMux I__16507 (
            .O(N__69500),
            .I(N__69495));
    LocalMux I__16506 (
            .O(N__69495),
            .I(\c0.n22701 ));
    InMux I__16505 (
            .O(N__69492),
            .I(N__69488));
    InMux I__16504 (
            .O(N__69491),
            .I(N__69485));
    LocalMux I__16503 (
            .O(N__69488),
            .I(N__69482));
    LocalMux I__16502 (
            .O(N__69485),
            .I(N__69475));
    Span4Mux_h I__16501 (
            .O(N__69482),
            .I(N__69475));
    InMux I__16500 (
            .O(N__69481),
            .I(N__69472));
    InMux I__16499 (
            .O(N__69480),
            .I(N__69469));
    Odrv4 I__16498 (
            .O(N__69475),
            .I(\c0.n5_adj_4323 ));
    LocalMux I__16497 (
            .O(N__69472),
            .I(\c0.n5_adj_4323 ));
    LocalMux I__16496 (
            .O(N__69469),
            .I(\c0.n5_adj_4323 ));
    InMux I__16495 (
            .O(N__69462),
            .I(N__69454));
    InMux I__16494 (
            .O(N__69461),
            .I(N__69454));
    InMux I__16493 (
            .O(N__69460),
            .I(N__69451));
    InMux I__16492 (
            .O(N__69459),
            .I(N__69447));
    LocalMux I__16491 (
            .O(N__69454),
            .I(N__69444));
    LocalMux I__16490 (
            .O(N__69451),
            .I(N__69441));
    InMux I__16489 (
            .O(N__69450),
            .I(N__69438));
    LocalMux I__16488 (
            .O(N__69447),
            .I(N__69434));
    Span4Mux_h I__16487 (
            .O(N__69444),
            .I(N__69431));
    Span4Mux_v I__16486 (
            .O(N__69441),
            .I(N__69426));
    LocalMux I__16485 (
            .O(N__69438),
            .I(N__69426));
    InMux I__16484 (
            .O(N__69437),
            .I(N__69423));
    Span4Mux_h I__16483 (
            .O(N__69434),
            .I(N__69420));
    Span4Mux_v I__16482 (
            .O(N__69431),
            .I(N__69415));
    Span4Mux_h I__16481 (
            .O(N__69426),
            .I(N__69415));
    LocalMux I__16480 (
            .O(N__69423),
            .I(N__69412));
    Span4Mux_v I__16479 (
            .O(N__69420),
            .I(N__69407));
    Span4Mux_h I__16478 (
            .O(N__69415),
            .I(N__69402));
    Span4Mux_v I__16477 (
            .O(N__69412),
            .I(N__69402));
    InMux I__16476 (
            .O(N__69411),
            .I(N__69399));
    InMux I__16475 (
            .O(N__69410),
            .I(N__69396));
    Odrv4 I__16474 (
            .O(N__69407),
            .I(n22101));
    Odrv4 I__16473 (
            .O(N__69402),
            .I(n22101));
    LocalMux I__16472 (
            .O(N__69399),
            .I(n22101));
    LocalMux I__16471 (
            .O(N__69396),
            .I(n22101));
    CascadeMux I__16470 (
            .O(N__69387),
            .I(\c0.n9_cascade_ ));
    CascadeMux I__16469 (
            .O(N__69384),
            .I(N__69381));
    InMux I__16468 (
            .O(N__69381),
            .I(N__69377));
    InMux I__16467 (
            .O(N__69380),
            .I(N__69373));
    LocalMux I__16466 (
            .O(N__69377),
            .I(N__69370));
    InMux I__16465 (
            .O(N__69376),
            .I(N__69367));
    LocalMux I__16464 (
            .O(N__69373),
            .I(N__69364));
    Span4Mux_v I__16463 (
            .O(N__69370),
            .I(N__69355));
    LocalMux I__16462 (
            .O(N__69367),
            .I(N__69355));
    Span4Mux_v I__16461 (
            .O(N__69364),
            .I(N__69355));
    CascadeMux I__16460 (
            .O(N__69363),
            .I(N__69351));
    CascadeMux I__16459 (
            .O(N__69362),
            .I(N__69348));
    Span4Mux_v I__16458 (
            .O(N__69355),
            .I(N__69345));
    InMux I__16457 (
            .O(N__69354),
            .I(N__69342));
    InMux I__16456 (
            .O(N__69351),
            .I(N__69337));
    InMux I__16455 (
            .O(N__69348),
            .I(N__69337));
    Odrv4 I__16454 (
            .O(N__69345),
            .I(\c0.data_in_frame_9_1 ));
    LocalMux I__16453 (
            .O(N__69342),
            .I(\c0.data_in_frame_9_1 ));
    LocalMux I__16452 (
            .O(N__69337),
            .I(\c0.data_in_frame_9_1 ));
    InMux I__16451 (
            .O(N__69330),
            .I(N__69326));
    InMux I__16450 (
            .O(N__69329),
            .I(N__69322));
    LocalMux I__16449 (
            .O(N__69326),
            .I(N__69317));
    CascadeMux I__16448 (
            .O(N__69325),
            .I(N__69314));
    LocalMux I__16447 (
            .O(N__69322),
            .I(N__69310));
    InMux I__16446 (
            .O(N__69321),
            .I(N__69305));
    InMux I__16445 (
            .O(N__69320),
            .I(N__69305));
    Span4Mux_h I__16444 (
            .O(N__69317),
            .I(N__69302));
    InMux I__16443 (
            .O(N__69314),
            .I(N__69298));
    InMux I__16442 (
            .O(N__69313),
            .I(N__69295));
    Span4Mux_h I__16441 (
            .O(N__69310),
            .I(N__69288));
    LocalMux I__16440 (
            .O(N__69305),
            .I(N__69288));
    Span4Mux_v I__16439 (
            .O(N__69302),
            .I(N__69288));
    InMux I__16438 (
            .O(N__69301),
            .I(N__69285));
    LocalMux I__16437 (
            .O(N__69298),
            .I(\c0.data_in_frame_8_6 ));
    LocalMux I__16436 (
            .O(N__69295),
            .I(\c0.data_in_frame_8_6 ));
    Odrv4 I__16435 (
            .O(N__69288),
            .I(\c0.data_in_frame_8_6 ));
    LocalMux I__16434 (
            .O(N__69285),
            .I(\c0.data_in_frame_8_6 ));
    CascadeMux I__16433 (
            .O(N__69276),
            .I(N__69272));
    InMux I__16432 (
            .O(N__69275),
            .I(N__69267));
    InMux I__16431 (
            .O(N__69272),
            .I(N__69267));
    LocalMux I__16430 (
            .O(N__69267),
            .I(\c0.data_in_frame_18_0 ));
    InMux I__16429 (
            .O(N__69264),
            .I(N__69255));
    InMux I__16428 (
            .O(N__69263),
            .I(N__69255));
    InMux I__16427 (
            .O(N__69262),
            .I(N__69255));
    LocalMux I__16426 (
            .O(N__69255),
            .I(data_in_frame_6_5));
    CascadeMux I__16425 (
            .O(N__69252),
            .I(N__69249));
    InMux I__16424 (
            .O(N__69249),
            .I(N__69246));
    LocalMux I__16423 (
            .O(N__69246),
            .I(N__69243));
    Span4Mux_h I__16422 (
            .O(N__69243),
            .I(N__69240));
    Odrv4 I__16421 (
            .O(N__69240),
            .I(\c0.n19_adj_4620 ));
    InMux I__16420 (
            .O(N__69237),
            .I(N__69228));
    InMux I__16419 (
            .O(N__69236),
            .I(N__69228));
    InMux I__16418 (
            .O(N__69235),
            .I(N__69228));
    LocalMux I__16417 (
            .O(N__69228),
            .I(N__69220));
    InMux I__16416 (
            .O(N__69227),
            .I(N__69215));
    InMux I__16415 (
            .O(N__69226),
            .I(N__69215));
    CascadeMux I__16414 (
            .O(N__69225),
            .I(N__69212));
    InMux I__16413 (
            .O(N__69224),
            .I(N__69205));
    InMux I__16412 (
            .O(N__69223),
            .I(N__69205));
    Span4Mux_v I__16411 (
            .O(N__69220),
            .I(N__69201));
    LocalMux I__16410 (
            .O(N__69215),
            .I(N__69196));
    InMux I__16409 (
            .O(N__69212),
            .I(N__69191));
    InMux I__16408 (
            .O(N__69211),
            .I(N__69186));
    InMux I__16407 (
            .O(N__69210),
            .I(N__69186));
    LocalMux I__16406 (
            .O(N__69205),
            .I(N__69177));
    InMux I__16405 (
            .O(N__69204),
            .I(N__69174));
    Span4Mux_v I__16404 (
            .O(N__69201),
            .I(N__69171));
    CascadeMux I__16403 (
            .O(N__69200),
            .I(N__69167));
    CascadeMux I__16402 (
            .O(N__69199),
            .I(N__69163));
    Span4Mux_v I__16401 (
            .O(N__69196),
            .I(N__69158));
    InMux I__16400 (
            .O(N__69195),
            .I(N__69151));
    InMux I__16399 (
            .O(N__69194),
            .I(N__69151));
    LocalMux I__16398 (
            .O(N__69191),
            .I(N__69147));
    LocalMux I__16397 (
            .O(N__69186),
            .I(N__69144));
    InMux I__16396 (
            .O(N__69185),
            .I(N__69141));
    InMux I__16395 (
            .O(N__69184),
            .I(N__69136));
    InMux I__16394 (
            .O(N__69183),
            .I(N__69136));
    InMux I__16393 (
            .O(N__69182),
            .I(N__69129));
    InMux I__16392 (
            .O(N__69181),
            .I(N__69129));
    InMux I__16391 (
            .O(N__69180),
            .I(N__69129));
    Span4Mux_h I__16390 (
            .O(N__69177),
            .I(N__69124));
    LocalMux I__16389 (
            .O(N__69174),
            .I(N__69124));
    Span4Mux_h I__16388 (
            .O(N__69171),
            .I(N__69121));
    CascadeMux I__16387 (
            .O(N__69170),
            .I(N__69118));
    InMux I__16386 (
            .O(N__69167),
            .I(N__69112));
    InMux I__16385 (
            .O(N__69166),
            .I(N__69112));
    InMux I__16384 (
            .O(N__69163),
            .I(N__69109));
    InMux I__16383 (
            .O(N__69162),
            .I(N__69104));
    InMux I__16382 (
            .O(N__69161),
            .I(N__69104));
    Sp12to4 I__16381 (
            .O(N__69158),
            .I(N__69101));
    InMux I__16380 (
            .O(N__69157),
            .I(N__69098));
    InMux I__16379 (
            .O(N__69156),
            .I(N__69095));
    LocalMux I__16378 (
            .O(N__69151),
            .I(N__69092));
    InMux I__16377 (
            .O(N__69150),
            .I(N__69088));
    Span4Mux_v I__16376 (
            .O(N__69147),
            .I(N__69085));
    Span4Mux_v I__16375 (
            .O(N__69144),
            .I(N__69078));
    LocalMux I__16374 (
            .O(N__69141),
            .I(N__69078));
    LocalMux I__16373 (
            .O(N__69136),
            .I(N__69078));
    LocalMux I__16372 (
            .O(N__69129),
            .I(N__69075));
    Span4Mux_h I__16371 (
            .O(N__69124),
            .I(N__69072));
    Sp12to4 I__16370 (
            .O(N__69121),
            .I(N__69069));
    InMux I__16369 (
            .O(N__69118),
            .I(N__69065));
    InMux I__16368 (
            .O(N__69117),
            .I(N__69062));
    LocalMux I__16367 (
            .O(N__69112),
            .I(N__69059));
    LocalMux I__16366 (
            .O(N__69109),
            .I(N__69050));
    LocalMux I__16365 (
            .O(N__69104),
            .I(N__69050));
    Span12Mux_s9_v I__16364 (
            .O(N__69101),
            .I(N__69050));
    LocalMux I__16363 (
            .O(N__69098),
            .I(N__69050));
    LocalMux I__16362 (
            .O(N__69095),
            .I(N__69047));
    Span4Mux_h I__16361 (
            .O(N__69092),
            .I(N__69044));
    InMux I__16360 (
            .O(N__69091),
            .I(N__69041));
    LocalMux I__16359 (
            .O(N__69088),
            .I(N__69038));
    Span4Mux_h I__16358 (
            .O(N__69085),
            .I(N__69035));
    Span4Mux_h I__16357 (
            .O(N__69078),
            .I(N__69032));
    Sp12to4 I__16356 (
            .O(N__69075),
            .I(N__69025));
    Sp12to4 I__16355 (
            .O(N__69072),
            .I(N__69025));
    Span12Mux_h I__16354 (
            .O(N__69069),
            .I(N__69025));
    InMux I__16353 (
            .O(N__69068),
            .I(N__69022));
    LocalMux I__16352 (
            .O(N__69065),
            .I(N__69019));
    LocalMux I__16351 (
            .O(N__69062),
            .I(N__69012));
    Span12Mux_s10_v I__16350 (
            .O(N__69059),
            .I(N__69012));
    Span12Mux_v I__16349 (
            .O(N__69050),
            .I(N__69012));
    Span4Mux_h I__16348 (
            .O(N__69047),
            .I(N__69007));
    Span4Mux_v I__16347 (
            .O(N__69044),
            .I(N__69007));
    LocalMux I__16346 (
            .O(N__69041),
            .I(N__69000));
    Span4Mux_v I__16345 (
            .O(N__69038),
            .I(N__69000));
    Span4Mux_v I__16344 (
            .O(N__69035),
            .I(N__69000));
    Sp12to4 I__16343 (
            .O(N__69032),
            .I(N__68995));
    Span12Mux_v I__16342 (
            .O(N__69025),
            .I(N__68995));
    LocalMux I__16341 (
            .O(N__69022),
            .I(\c0.n9 ));
    Odrv4 I__16340 (
            .O(N__69019),
            .I(\c0.n9 ));
    Odrv12 I__16339 (
            .O(N__69012),
            .I(\c0.n9 ));
    Odrv4 I__16338 (
            .O(N__69007),
            .I(\c0.n9 ));
    Odrv4 I__16337 (
            .O(N__69000),
            .I(\c0.n9 ));
    Odrv12 I__16336 (
            .O(N__68995),
            .I(\c0.n9 ));
    InMux I__16335 (
            .O(N__68982),
            .I(N__68979));
    LocalMux I__16334 (
            .O(N__68979),
            .I(N__68976));
    Span4Mux_v I__16333 (
            .O(N__68976),
            .I(N__68973));
    Odrv4 I__16332 (
            .O(N__68973),
            .I(\c0.n22392 ));
    InMux I__16331 (
            .O(N__68970),
            .I(N__68966));
    CascadeMux I__16330 (
            .O(N__68969),
            .I(N__68963));
    LocalMux I__16329 (
            .O(N__68966),
            .I(N__68960));
    InMux I__16328 (
            .O(N__68963),
            .I(N__68954));
    Span4Mux_h I__16327 (
            .O(N__68960),
            .I(N__68951));
    InMux I__16326 (
            .O(N__68959),
            .I(N__68948));
    InMux I__16325 (
            .O(N__68958),
            .I(N__68945));
    InMux I__16324 (
            .O(N__68957),
            .I(N__68942));
    LocalMux I__16323 (
            .O(N__68954),
            .I(\c0.data_in_frame_4_3 ));
    Odrv4 I__16322 (
            .O(N__68951),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__16321 (
            .O(N__68948),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__16320 (
            .O(N__68945),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__16319 (
            .O(N__68942),
            .I(\c0.data_in_frame_4_3 ));
    CascadeMux I__16318 (
            .O(N__68931),
            .I(\c0.n6_adj_4687_cascade_ ));
    InMux I__16317 (
            .O(N__68928),
            .I(N__68924));
    CascadeMux I__16316 (
            .O(N__68927),
            .I(N__68920));
    LocalMux I__16315 (
            .O(N__68924),
            .I(N__68917));
    InMux I__16314 (
            .O(N__68923),
            .I(N__68914));
    InMux I__16313 (
            .O(N__68920),
            .I(N__68911));
    Span4Mux_v I__16312 (
            .O(N__68917),
            .I(N__68908));
    LocalMux I__16311 (
            .O(N__68914),
            .I(\c0.n23274 ));
    LocalMux I__16310 (
            .O(N__68911),
            .I(\c0.n23274 ));
    Odrv4 I__16309 (
            .O(N__68908),
            .I(\c0.n23274 ));
    InMux I__16308 (
            .O(N__68901),
            .I(N__68895));
    InMux I__16307 (
            .O(N__68900),
            .I(N__68895));
    LocalMux I__16306 (
            .O(N__68895),
            .I(\c0.n23282 ));
    CascadeMux I__16305 (
            .O(N__68892),
            .I(\c0.n23274_cascade_ ));
    InMux I__16304 (
            .O(N__68889),
            .I(N__68886));
    LocalMux I__16303 (
            .O(N__68886),
            .I(\c0.n20_adj_4316 ));
    InMux I__16302 (
            .O(N__68883),
            .I(N__68880));
    LocalMux I__16301 (
            .O(N__68880),
            .I(N__68876));
    CascadeMux I__16300 (
            .O(N__68879),
            .I(N__68873));
    Span4Mux_v I__16299 (
            .O(N__68876),
            .I(N__68870));
    InMux I__16298 (
            .O(N__68873),
            .I(N__68867));
    Span4Mux_h I__16297 (
            .O(N__68870),
            .I(N__68864));
    LocalMux I__16296 (
            .O(N__68867),
            .I(N__68861));
    Span4Mux_v I__16295 (
            .O(N__68864),
            .I(N__68858));
    Span12Mux_h I__16294 (
            .O(N__68861),
            .I(N__68855));
    Odrv4 I__16293 (
            .O(N__68858),
            .I(\c0.n29_adj_4287 ));
    Odrv12 I__16292 (
            .O(N__68855),
            .I(\c0.n29_adj_4287 ));
    InMux I__16291 (
            .O(N__68850),
            .I(N__68837));
    InMux I__16290 (
            .O(N__68849),
            .I(N__68832));
    InMux I__16289 (
            .O(N__68848),
            .I(N__68832));
    InMux I__16288 (
            .O(N__68847),
            .I(N__68829));
    InMux I__16287 (
            .O(N__68846),
            .I(N__68826));
    InMux I__16286 (
            .O(N__68845),
            .I(N__68821));
    InMux I__16285 (
            .O(N__68844),
            .I(N__68821));
    InMux I__16284 (
            .O(N__68843),
            .I(N__68814));
    InMux I__16283 (
            .O(N__68842),
            .I(N__68814));
    InMux I__16282 (
            .O(N__68841),
            .I(N__68814));
    InMux I__16281 (
            .O(N__68840),
            .I(N__68811));
    LocalMux I__16280 (
            .O(N__68837),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__16279 (
            .O(N__68832),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__16278 (
            .O(N__68829),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__16277 (
            .O(N__68826),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__16276 (
            .O(N__68821),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__16275 (
            .O(N__68814),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__16274 (
            .O(N__68811),
            .I(\c0.data_in_frame_0_2 ));
    CascadeMux I__16273 (
            .O(N__68796),
            .I(N__68790));
    InMux I__16272 (
            .O(N__68795),
            .I(N__68787));
    InMux I__16271 (
            .O(N__68794),
            .I(N__68782));
    InMux I__16270 (
            .O(N__68793),
            .I(N__68782));
    InMux I__16269 (
            .O(N__68790),
            .I(N__68777));
    LocalMux I__16268 (
            .O(N__68787),
            .I(N__68774));
    LocalMux I__16267 (
            .O(N__68782),
            .I(N__68771));
    InMux I__16266 (
            .O(N__68781),
            .I(N__68766));
    InMux I__16265 (
            .O(N__68780),
            .I(N__68766));
    LocalMux I__16264 (
            .O(N__68777),
            .I(\c0.data_in_frame_2_3 ));
    Odrv4 I__16263 (
            .O(N__68774),
            .I(\c0.data_in_frame_2_3 ));
    Odrv4 I__16262 (
            .O(N__68771),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__16261 (
            .O(N__68766),
            .I(\c0.data_in_frame_2_3 ));
    InMux I__16260 (
            .O(N__68757),
            .I(N__68753));
    CascadeMux I__16259 (
            .O(N__68756),
            .I(N__68746));
    LocalMux I__16258 (
            .O(N__68753),
            .I(N__68743));
    InMux I__16257 (
            .O(N__68752),
            .I(N__68740));
    InMux I__16256 (
            .O(N__68751),
            .I(N__68737));
    InMux I__16255 (
            .O(N__68750),
            .I(N__68734));
    CascadeMux I__16254 (
            .O(N__68749),
            .I(N__68729));
    InMux I__16253 (
            .O(N__68746),
            .I(N__68723));
    Span4Mux_h I__16252 (
            .O(N__68743),
            .I(N__68716));
    LocalMux I__16251 (
            .O(N__68740),
            .I(N__68716));
    LocalMux I__16250 (
            .O(N__68737),
            .I(N__68716));
    LocalMux I__16249 (
            .O(N__68734),
            .I(N__68713));
    InMux I__16248 (
            .O(N__68733),
            .I(N__68710));
    InMux I__16247 (
            .O(N__68732),
            .I(N__68707));
    InMux I__16246 (
            .O(N__68729),
            .I(N__68702));
    InMux I__16245 (
            .O(N__68728),
            .I(N__68702));
    InMux I__16244 (
            .O(N__68727),
            .I(N__68699));
    InMux I__16243 (
            .O(N__68726),
            .I(N__68696));
    LocalMux I__16242 (
            .O(N__68723),
            .I(\c0.data_in_frame_0_1 ));
    Odrv4 I__16241 (
            .O(N__68716),
            .I(\c0.data_in_frame_0_1 ));
    Odrv4 I__16240 (
            .O(N__68713),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__16239 (
            .O(N__68710),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__16238 (
            .O(N__68707),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__16237 (
            .O(N__68702),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__16236 (
            .O(N__68699),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__16235 (
            .O(N__68696),
            .I(\c0.data_in_frame_0_1 ));
    InMux I__16234 (
            .O(N__68679),
            .I(N__68672));
    InMux I__16233 (
            .O(N__68678),
            .I(N__68672));
    InMux I__16232 (
            .O(N__68677),
            .I(N__68666));
    LocalMux I__16231 (
            .O(N__68672),
            .I(N__68663));
    InMux I__16230 (
            .O(N__68671),
            .I(N__68660));
    InMux I__16229 (
            .O(N__68670),
            .I(N__68655));
    InMux I__16228 (
            .O(N__68669),
            .I(N__68655));
    LocalMux I__16227 (
            .O(N__68666),
            .I(\c0.data_in_frame_4_4 ));
    Odrv12 I__16226 (
            .O(N__68663),
            .I(\c0.data_in_frame_4_4 ));
    LocalMux I__16225 (
            .O(N__68660),
            .I(\c0.data_in_frame_4_4 ));
    LocalMux I__16224 (
            .O(N__68655),
            .I(\c0.data_in_frame_4_4 ));
    InMux I__16223 (
            .O(N__68646),
            .I(N__68642));
    InMux I__16222 (
            .O(N__68645),
            .I(N__68639));
    LocalMux I__16221 (
            .O(N__68642),
            .I(\c0.n23276 ));
    LocalMux I__16220 (
            .O(N__68639),
            .I(\c0.n23276 ));
    InMux I__16219 (
            .O(N__68634),
            .I(N__68628));
    InMux I__16218 (
            .O(N__68633),
            .I(N__68628));
    LocalMux I__16217 (
            .O(N__68628),
            .I(N__68625));
    Span4Mux_v I__16216 (
            .O(N__68625),
            .I(N__68619));
    InMux I__16215 (
            .O(N__68624),
            .I(N__68612));
    InMux I__16214 (
            .O(N__68623),
            .I(N__68612));
    InMux I__16213 (
            .O(N__68622),
            .I(N__68612));
    Odrv4 I__16212 (
            .O(N__68619),
            .I(\c0.n22322 ));
    LocalMux I__16211 (
            .O(N__68612),
            .I(\c0.n22322 ));
    CascadeMux I__16210 (
            .O(N__68607),
            .I(\c0.n23276_cascade_ ));
    InMux I__16209 (
            .O(N__68604),
            .I(N__68601));
    LocalMux I__16208 (
            .O(N__68601),
            .I(N__68597));
    InMux I__16207 (
            .O(N__68600),
            .I(N__68594));
    Span4Mux_v I__16206 (
            .O(N__68597),
            .I(N__68588));
    LocalMux I__16205 (
            .O(N__68594),
            .I(N__68588));
    InMux I__16204 (
            .O(N__68593),
            .I(N__68585));
    Span4Mux_h I__16203 (
            .O(N__68588),
            .I(N__68582));
    LocalMux I__16202 (
            .O(N__68585),
            .I(N__68579));
    Span4Mux_h I__16201 (
            .O(N__68582),
            .I(N__68576));
    Odrv4 I__16200 (
            .O(N__68579),
            .I(\c0.n25 ));
    Odrv4 I__16199 (
            .O(N__68576),
            .I(\c0.n25 ));
    InMux I__16198 (
            .O(N__68571),
            .I(N__68567));
    InMux I__16197 (
            .O(N__68570),
            .I(N__68564));
    LocalMux I__16196 (
            .O(N__68567),
            .I(\c0.n24_adj_4213 ));
    LocalMux I__16195 (
            .O(N__68564),
            .I(\c0.n24_adj_4213 ));
    CascadeMux I__16194 (
            .O(N__68559),
            .I(\c0.n8_cascade_ ));
    InMux I__16193 (
            .O(N__68556),
            .I(N__68552));
    CascadeMux I__16192 (
            .O(N__68555),
            .I(N__68549));
    LocalMux I__16191 (
            .O(N__68552),
            .I(N__68546));
    InMux I__16190 (
            .O(N__68549),
            .I(N__68539));
    Span4Mux_h I__16189 (
            .O(N__68546),
            .I(N__68536));
    InMux I__16188 (
            .O(N__68545),
            .I(N__68533));
    InMux I__16187 (
            .O(N__68544),
            .I(N__68528));
    CascadeMux I__16186 (
            .O(N__68543),
            .I(N__68524));
    CascadeMux I__16185 (
            .O(N__68542),
            .I(N__68521));
    LocalMux I__16184 (
            .O(N__68539),
            .I(N__68518));
    Span4Mux_v I__16183 (
            .O(N__68536),
            .I(N__68513));
    LocalMux I__16182 (
            .O(N__68533),
            .I(N__68513));
    InMux I__16181 (
            .O(N__68532),
            .I(N__68507));
    InMux I__16180 (
            .O(N__68531),
            .I(N__68504));
    LocalMux I__16179 (
            .O(N__68528),
            .I(N__68501));
    InMux I__16178 (
            .O(N__68527),
            .I(N__68498));
    InMux I__16177 (
            .O(N__68524),
            .I(N__68490));
    InMux I__16176 (
            .O(N__68521),
            .I(N__68490));
    Span4Mux_v I__16175 (
            .O(N__68518),
            .I(N__68485));
    Span4Mux_v I__16174 (
            .O(N__68513),
            .I(N__68485));
    InMux I__16173 (
            .O(N__68512),
            .I(N__68482));
    InMux I__16172 (
            .O(N__68511),
            .I(N__68477));
    InMux I__16171 (
            .O(N__68510),
            .I(N__68477));
    LocalMux I__16170 (
            .O(N__68507),
            .I(N__68472));
    LocalMux I__16169 (
            .O(N__68504),
            .I(N__68472));
    Span4Mux_v I__16168 (
            .O(N__68501),
            .I(N__68467));
    LocalMux I__16167 (
            .O(N__68498),
            .I(N__68467));
    InMux I__16166 (
            .O(N__68497),
            .I(N__68464));
    InMux I__16165 (
            .O(N__68496),
            .I(N__68459));
    InMux I__16164 (
            .O(N__68495),
            .I(N__68459));
    LocalMux I__16163 (
            .O(N__68490),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__16162 (
            .O(N__68485),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__16161 (
            .O(N__68482),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__16160 (
            .O(N__68477),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__16159 (
            .O(N__68472),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__16158 (
            .O(N__68467),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__16157 (
            .O(N__68464),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__16156 (
            .O(N__68459),
            .I(\c0.data_in_frame_0_4 ));
    InMux I__16155 (
            .O(N__68442),
            .I(N__68438));
    InMux I__16154 (
            .O(N__68441),
            .I(N__68434));
    LocalMux I__16153 (
            .O(N__68438),
            .I(N__68429));
    InMux I__16152 (
            .O(N__68437),
            .I(N__68426));
    LocalMux I__16151 (
            .O(N__68434),
            .I(N__68423));
    InMux I__16150 (
            .O(N__68433),
            .I(N__68419));
    InMux I__16149 (
            .O(N__68432),
            .I(N__68416));
    Span4Mux_h I__16148 (
            .O(N__68429),
            .I(N__68411));
    LocalMux I__16147 (
            .O(N__68426),
            .I(N__68411));
    Span4Mux_v I__16146 (
            .O(N__68423),
            .I(N__68408));
    InMux I__16145 (
            .O(N__68422),
            .I(N__68405));
    LocalMux I__16144 (
            .O(N__68419),
            .I(N__68402));
    LocalMux I__16143 (
            .O(N__68416),
            .I(N__68399));
    Span4Mux_h I__16142 (
            .O(N__68411),
            .I(N__68396));
    Sp12to4 I__16141 (
            .O(N__68408),
            .I(N__68390));
    LocalMux I__16140 (
            .O(N__68405),
            .I(N__68390));
    Span12Mux_h I__16139 (
            .O(N__68402),
            .I(N__68387));
    Span4Mux_h I__16138 (
            .O(N__68399),
            .I(N__68382));
    Span4Mux_h I__16137 (
            .O(N__68396),
            .I(N__68382));
    InMux I__16136 (
            .O(N__68395),
            .I(N__68379));
    Odrv12 I__16135 (
            .O(N__68390),
            .I(n22121));
    Odrv12 I__16134 (
            .O(N__68387),
            .I(n22121));
    Odrv4 I__16133 (
            .O(N__68382),
            .I(n22121));
    LocalMux I__16132 (
            .O(N__68379),
            .I(n22121));
    InMux I__16131 (
            .O(N__68370),
            .I(N__68367));
    LocalMux I__16130 (
            .O(N__68367),
            .I(N__68362));
    InMux I__16129 (
            .O(N__68366),
            .I(N__68359));
    InMux I__16128 (
            .O(N__68365),
            .I(N__68356));
    Span4Mux_v I__16127 (
            .O(N__68362),
            .I(N__68353));
    LocalMux I__16126 (
            .O(N__68359),
            .I(N__68350));
    LocalMux I__16125 (
            .O(N__68356),
            .I(N__68346));
    Span4Mux_h I__16124 (
            .O(N__68353),
            .I(N__68343));
    Span4Mux_v I__16123 (
            .O(N__68350),
            .I(N__68340));
    InMux I__16122 (
            .O(N__68349),
            .I(N__68337));
    Span12Mux_h I__16121 (
            .O(N__68346),
            .I(N__68334));
    Span4Mux_h I__16120 (
            .O(N__68343),
            .I(N__68331));
    Span4Mux_h I__16119 (
            .O(N__68340),
            .I(N__68328));
    LocalMux I__16118 (
            .O(N__68337),
            .I(\c0.data_in_frame_26_3 ));
    Odrv12 I__16117 (
            .O(N__68334),
            .I(\c0.data_in_frame_26_3 ));
    Odrv4 I__16116 (
            .O(N__68331),
            .I(\c0.data_in_frame_26_3 ));
    Odrv4 I__16115 (
            .O(N__68328),
            .I(\c0.data_in_frame_26_3 ));
    CascadeMux I__16114 (
            .O(N__68319),
            .I(\c0.n22362_cascade_ ));
    InMux I__16113 (
            .O(N__68316),
            .I(N__68313));
    LocalMux I__16112 (
            .O(N__68313),
            .I(N__68308));
    InMux I__16111 (
            .O(N__68312),
            .I(N__68305));
    InMux I__16110 (
            .O(N__68311),
            .I(N__68302));
    Odrv4 I__16109 (
            .O(N__68308),
            .I(\c0.n12559 ));
    LocalMux I__16108 (
            .O(N__68305),
            .I(\c0.n12559 ));
    LocalMux I__16107 (
            .O(N__68302),
            .I(\c0.n12559 ));
    CascadeMux I__16106 (
            .O(N__68295),
            .I(N__68292));
    InMux I__16105 (
            .O(N__68292),
            .I(N__68289));
    LocalMux I__16104 (
            .O(N__68289),
            .I(N__68286));
    Span4Mux_h I__16103 (
            .O(N__68286),
            .I(N__68283));
    Odrv4 I__16102 (
            .O(N__68283),
            .I(\c0.n13_adj_4527 ));
    InMux I__16101 (
            .O(N__68280),
            .I(N__68275));
    InMux I__16100 (
            .O(N__68279),
            .I(N__68270));
    InMux I__16099 (
            .O(N__68278),
            .I(N__68270));
    LocalMux I__16098 (
            .O(N__68275),
            .I(N__68267));
    LocalMux I__16097 (
            .O(N__68270),
            .I(\c0.n20802 ));
    Odrv4 I__16096 (
            .O(N__68267),
            .I(\c0.n20802 ));
    InMux I__16095 (
            .O(N__68262),
            .I(N__68258));
    InMux I__16094 (
            .O(N__68261),
            .I(N__68255));
    LocalMux I__16093 (
            .O(N__68258),
            .I(N__68252));
    LocalMux I__16092 (
            .O(N__68255),
            .I(\c0.n20358 ));
    Odrv12 I__16091 (
            .O(N__68252),
            .I(\c0.n20358 ));
    InMux I__16090 (
            .O(N__68247),
            .I(N__68244));
    LocalMux I__16089 (
            .O(N__68244),
            .I(\c0.n12_adj_4491 ));
    CascadeMux I__16088 (
            .O(N__68241),
            .I(N__68237));
    InMux I__16087 (
            .O(N__68240),
            .I(N__68232));
    InMux I__16086 (
            .O(N__68237),
            .I(N__68232));
    LocalMux I__16085 (
            .O(N__68232),
            .I(\c0.data_in_frame_28_6 ));
    InMux I__16084 (
            .O(N__68229),
            .I(N__68223));
    InMux I__16083 (
            .O(N__68228),
            .I(N__68223));
    LocalMux I__16082 (
            .O(N__68223),
            .I(N__68220));
    Odrv4 I__16081 (
            .O(N__68220),
            .I(\c0.data_in_frame_28_4 ));
    InMux I__16080 (
            .O(N__68217),
            .I(N__68212));
    CascadeMux I__16079 (
            .O(N__68216),
            .I(N__68209));
    InMux I__16078 (
            .O(N__68215),
            .I(N__68206));
    LocalMux I__16077 (
            .O(N__68212),
            .I(N__68203));
    InMux I__16076 (
            .O(N__68209),
            .I(N__68200));
    LocalMux I__16075 (
            .O(N__68206),
            .I(N__68197));
    Odrv12 I__16074 (
            .O(N__68203),
            .I(\c0.n13904 ));
    LocalMux I__16073 (
            .O(N__68200),
            .I(\c0.n13904 ));
    Odrv4 I__16072 (
            .O(N__68197),
            .I(\c0.n13904 ));
    InMux I__16071 (
            .O(N__68190),
            .I(N__68186));
    InMux I__16070 (
            .O(N__68189),
            .I(N__68183));
    LocalMux I__16069 (
            .O(N__68186),
            .I(N__68180));
    LocalMux I__16068 (
            .O(N__68183),
            .I(N__68177));
    Span4Mux_h I__16067 (
            .O(N__68180),
            .I(N__68174));
    Sp12to4 I__16066 (
            .O(N__68177),
            .I(N__68171));
    Span4Mux_v I__16065 (
            .O(N__68174),
            .I(N__68168));
    Odrv12 I__16064 (
            .O(N__68171),
            .I(\c0.n28_adj_4286 ));
    Odrv4 I__16063 (
            .O(N__68168),
            .I(\c0.n28_adj_4286 ));
    InMux I__16062 (
            .O(N__68163),
            .I(N__68157));
    InMux I__16061 (
            .O(N__68162),
            .I(N__68150));
    InMux I__16060 (
            .O(N__68161),
            .I(N__68150));
    InMux I__16059 (
            .O(N__68160),
            .I(N__68150));
    LocalMux I__16058 (
            .O(N__68157),
            .I(data_in_frame_5_0));
    LocalMux I__16057 (
            .O(N__68150),
            .I(data_in_frame_5_0));
    InMux I__16056 (
            .O(N__68145),
            .I(N__68142));
    LocalMux I__16055 (
            .O(N__68142),
            .I(N__68137));
    InMux I__16054 (
            .O(N__68141),
            .I(N__68132));
    InMux I__16053 (
            .O(N__68140),
            .I(N__68132));
    Odrv4 I__16052 (
            .O(N__68137),
            .I(\c0.n23302 ));
    LocalMux I__16051 (
            .O(N__68132),
            .I(\c0.n23302 ));
    InMux I__16050 (
            .O(N__68127),
            .I(N__68123));
    InMux I__16049 (
            .O(N__68126),
            .I(N__68117));
    LocalMux I__16048 (
            .O(N__68123),
            .I(N__68114));
    InMux I__16047 (
            .O(N__68122),
            .I(N__68111));
    CascadeMux I__16046 (
            .O(N__68121),
            .I(N__68105));
    InMux I__16045 (
            .O(N__68120),
            .I(N__68102));
    LocalMux I__16044 (
            .O(N__68117),
            .I(N__68097));
    Span4Mux_v I__16043 (
            .O(N__68114),
            .I(N__68097));
    LocalMux I__16042 (
            .O(N__68111),
            .I(N__68090));
    InMux I__16041 (
            .O(N__68110),
            .I(N__68083));
    InMux I__16040 (
            .O(N__68109),
            .I(N__68083));
    InMux I__16039 (
            .O(N__68108),
            .I(N__68083));
    InMux I__16038 (
            .O(N__68105),
            .I(N__68078));
    LocalMux I__16037 (
            .O(N__68102),
            .I(N__68073));
    Span4Mux_h I__16036 (
            .O(N__68097),
            .I(N__68073));
    InMux I__16035 (
            .O(N__68096),
            .I(N__68068));
    InMux I__16034 (
            .O(N__68095),
            .I(N__68068));
    InMux I__16033 (
            .O(N__68094),
            .I(N__68063));
    InMux I__16032 (
            .O(N__68093),
            .I(N__68063));
    Span4Mux_h I__16031 (
            .O(N__68090),
            .I(N__68058));
    LocalMux I__16030 (
            .O(N__68083),
            .I(N__68058));
    InMux I__16029 (
            .O(N__68082),
            .I(N__68053));
    InMux I__16028 (
            .O(N__68081),
            .I(N__68053));
    LocalMux I__16027 (
            .O(N__68078),
            .I(\c0.data_in_frame_0_3 ));
    Odrv4 I__16026 (
            .O(N__68073),
            .I(\c0.data_in_frame_0_3 ));
    LocalMux I__16025 (
            .O(N__68068),
            .I(\c0.data_in_frame_0_3 ));
    LocalMux I__16024 (
            .O(N__68063),
            .I(\c0.data_in_frame_0_3 ));
    Odrv4 I__16023 (
            .O(N__68058),
            .I(\c0.data_in_frame_0_3 ));
    LocalMux I__16022 (
            .O(N__68053),
            .I(\c0.data_in_frame_0_3 ));
    CascadeMux I__16021 (
            .O(N__68040),
            .I(N__68035));
    CascadeMux I__16020 (
            .O(N__68039),
            .I(N__68031));
    InMux I__16019 (
            .O(N__68038),
            .I(N__68025));
    InMux I__16018 (
            .O(N__68035),
            .I(N__68022));
    InMux I__16017 (
            .O(N__68034),
            .I(N__68019));
    InMux I__16016 (
            .O(N__68031),
            .I(N__68014));
    InMux I__16015 (
            .O(N__68030),
            .I(N__68014));
    InMux I__16014 (
            .O(N__68029),
            .I(N__68009));
    InMux I__16013 (
            .O(N__68028),
            .I(N__68009));
    LocalMux I__16012 (
            .O(N__68025),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__16011 (
            .O(N__68022),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__16010 (
            .O(N__68019),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__16009 (
            .O(N__68014),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__16008 (
            .O(N__68009),
            .I(\c0.data_in_frame_2_4 ));
    InMux I__16007 (
            .O(N__67998),
            .I(N__67995));
    LocalMux I__16006 (
            .O(N__67995),
            .I(N__67992));
    Span12Mux_h I__16005 (
            .O(N__67992),
            .I(N__67989));
    Odrv12 I__16004 (
            .O(N__67989),
            .I(\c0.n42_adj_4746 ));
    InMux I__16003 (
            .O(N__67986),
            .I(N__67981));
    InMux I__16002 (
            .O(N__67985),
            .I(N__67978));
    CascadeMux I__16001 (
            .O(N__67984),
            .I(N__67975));
    LocalMux I__16000 (
            .O(N__67981),
            .I(N__67972));
    LocalMux I__15999 (
            .O(N__67978),
            .I(N__67969));
    InMux I__15998 (
            .O(N__67975),
            .I(N__67964));
    Span4Mux_v I__15997 (
            .O(N__67972),
            .I(N__67959));
    Span4Mux_h I__15996 (
            .O(N__67969),
            .I(N__67959));
    InMux I__15995 (
            .O(N__67968),
            .I(N__67956));
    InMux I__15994 (
            .O(N__67967),
            .I(N__67953));
    LocalMux I__15993 (
            .O(N__67964),
            .I(\c0.data_in_frame_7_1 ));
    Odrv4 I__15992 (
            .O(N__67959),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__15991 (
            .O(N__67956),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__15990 (
            .O(N__67953),
            .I(\c0.data_in_frame_7_1 ));
    CascadeMux I__15989 (
            .O(N__67944),
            .I(N__67938));
    CascadeMux I__15988 (
            .O(N__67943),
            .I(N__67935));
    InMux I__15987 (
            .O(N__67942),
            .I(N__67931));
    InMux I__15986 (
            .O(N__67941),
            .I(N__67928));
    InMux I__15985 (
            .O(N__67938),
            .I(N__67925));
    InMux I__15984 (
            .O(N__67935),
            .I(N__67922));
    InMux I__15983 (
            .O(N__67934),
            .I(N__67919));
    LocalMux I__15982 (
            .O(N__67931),
            .I(N__67916));
    LocalMux I__15981 (
            .O(N__67928),
            .I(N__67911));
    LocalMux I__15980 (
            .O(N__67925),
            .I(N__67908));
    LocalMux I__15979 (
            .O(N__67922),
            .I(N__67903));
    LocalMux I__15978 (
            .O(N__67919),
            .I(N__67903));
    Span4Mux_h I__15977 (
            .O(N__67916),
            .I(N__67900));
    InMux I__15976 (
            .O(N__67915),
            .I(N__67895));
    InMux I__15975 (
            .O(N__67914),
            .I(N__67895));
    Odrv4 I__15974 (
            .O(N__67911),
            .I(\c0.data_in_frame_2_5 ));
    Odrv4 I__15973 (
            .O(N__67908),
            .I(\c0.data_in_frame_2_5 ));
    Odrv4 I__15972 (
            .O(N__67903),
            .I(\c0.data_in_frame_2_5 ));
    Odrv4 I__15971 (
            .O(N__67900),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__15970 (
            .O(N__67895),
            .I(\c0.data_in_frame_2_5 ));
    InMux I__15969 (
            .O(N__67884),
            .I(N__67880));
    InMux I__15968 (
            .O(N__67883),
            .I(N__67877));
    LocalMux I__15967 (
            .O(N__67880),
            .I(N__67874));
    LocalMux I__15966 (
            .O(N__67877),
            .I(N__67870));
    Span4Mux_v I__15965 (
            .O(N__67874),
            .I(N__67867));
    CascadeMux I__15964 (
            .O(N__67873),
            .I(N__67864));
    Span4Mux_v I__15963 (
            .O(N__67870),
            .I(N__67859));
    Sp12to4 I__15962 (
            .O(N__67867),
            .I(N__67856));
    InMux I__15961 (
            .O(N__67864),
            .I(N__67853));
    CascadeMux I__15960 (
            .O(N__67863),
            .I(N__67850));
    InMux I__15959 (
            .O(N__67862),
            .I(N__67847));
    Span4Mux_h I__15958 (
            .O(N__67859),
            .I(N__67844));
    Span12Mux_h I__15957 (
            .O(N__67856),
            .I(N__67841));
    LocalMux I__15956 (
            .O(N__67853),
            .I(N__67838));
    InMux I__15955 (
            .O(N__67850),
            .I(N__67835));
    LocalMux I__15954 (
            .O(N__67847),
            .I(\c0.data_in_frame_27_2 ));
    Odrv4 I__15953 (
            .O(N__67844),
            .I(\c0.data_in_frame_27_2 ));
    Odrv12 I__15952 (
            .O(N__67841),
            .I(\c0.data_in_frame_27_2 ));
    Odrv12 I__15951 (
            .O(N__67838),
            .I(\c0.data_in_frame_27_2 ));
    LocalMux I__15950 (
            .O(N__67835),
            .I(\c0.data_in_frame_27_2 ));
    InMux I__15949 (
            .O(N__67824),
            .I(N__67821));
    LocalMux I__15948 (
            .O(N__67821),
            .I(N__67816));
    InMux I__15947 (
            .O(N__67820),
            .I(N__67813));
    InMux I__15946 (
            .O(N__67819),
            .I(N__67810));
    Span4Mux_v I__15945 (
            .O(N__67816),
            .I(N__67805));
    LocalMux I__15944 (
            .O(N__67813),
            .I(N__67805));
    LocalMux I__15943 (
            .O(N__67810),
            .I(N__67802));
    Odrv4 I__15942 (
            .O(N__67805),
            .I(\c0.n25_adj_4469 ));
    Odrv4 I__15941 (
            .O(N__67802),
            .I(\c0.n25_adj_4469 ));
    InMux I__15940 (
            .O(N__67797),
            .I(N__67794));
    LocalMux I__15939 (
            .O(N__67794),
            .I(N__67789));
    InMux I__15938 (
            .O(N__67793),
            .I(N__67786));
    InMux I__15937 (
            .O(N__67792),
            .I(N__67783));
    Span4Mux_h I__15936 (
            .O(N__67789),
            .I(N__67780));
    LocalMux I__15935 (
            .O(N__67786),
            .I(\c0.n26_adj_4470 ));
    LocalMux I__15934 (
            .O(N__67783),
            .I(\c0.n26_adj_4470 ));
    Odrv4 I__15933 (
            .O(N__67780),
            .I(\c0.n26_adj_4470 ));
    InMux I__15932 (
            .O(N__67773),
            .I(N__67770));
    LocalMux I__15931 (
            .O(N__67770),
            .I(\c0.n39_adj_4467 ));
    InMux I__15930 (
            .O(N__67767),
            .I(N__67764));
    LocalMux I__15929 (
            .O(N__67764),
            .I(\c0.n38_adj_4468 ));
    InMux I__15928 (
            .O(N__67761),
            .I(N__67758));
    LocalMux I__15927 (
            .O(N__67758),
            .I(N__67755));
    Odrv4 I__15926 (
            .O(N__67755),
            .I(\c0.n37_adj_4473 ));
    CascadeMux I__15925 (
            .O(N__67752),
            .I(\c0.n44_adj_4471_cascade_ ));
    InMux I__15924 (
            .O(N__67749),
            .I(N__67745));
    InMux I__15923 (
            .O(N__67748),
            .I(N__67742));
    LocalMux I__15922 (
            .O(N__67745),
            .I(N__67739));
    LocalMux I__15921 (
            .O(N__67742),
            .I(N__67736));
    Span4Mux_v I__15920 (
            .O(N__67739),
            .I(N__67733));
    Span4Mux_v I__15919 (
            .O(N__67736),
            .I(N__67730));
    Odrv4 I__15918 (
            .O(N__67733),
            .I(\c0.n45_adj_4476 ));
    Odrv4 I__15917 (
            .O(N__67730),
            .I(\c0.n45_adj_4476 ));
    InMux I__15916 (
            .O(N__67725),
            .I(N__67722));
    LocalMux I__15915 (
            .O(N__67722),
            .I(N__67719));
    Odrv12 I__15914 (
            .O(N__67719),
            .I(\c0.n14_adj_4529 ));
    InMux I__15913 (
            .O(N__67716),
            .I(N__67713));
    LocalMux I__15912 (
            .O(N__67713),
            .I(N__67710));
    Span4Mux_h I__15911 (
            .O(N__67710),
            .I(N__67707));
    Span4Mux_v I__15910 (
            .O(N__67707),
            .I(N__67703));
    InMux I__15909 (
            .O(N__67706),
            .I(N__67700));
    Odrv4 I__15908 (
            .O(N__67703),
            .I(\c0.n15_adj_4508 ));
    LocalMux I__15907 (
            .O(N__67700),
            .I(\c0.n15_adj_4508 ));
    CascadeMux I__15906 (
            .O(N__67695),
            .I(\c0.n24362_cascade_ ));
    InMux I__15905 (
            .O(N__67692),
            .I(N__67689));
    LocalMux I__15904 (
            .O(N__67689),
            .I(N__67686));
    Span4Mux_h I__15903 (
            .O(N__67686),
            .I(N__67683));
    Odrv4 I__15902 (
            .O(N__67683),
            .I(\c0.n18_adj_4475 ));
    InMux I__15901 (
            .O(N__67680),
            .I(N__67677));
    LocalMux I__15900 (
            .O(N__67677),
            .I(N__67674));
    Span4Mux_v I__15899 (
            .O(N__67674),
            .I(N__67671));
    Span4Mux_h I__15898 (
            .O(N__67671),
            .I(N__67668));
    Odrv4 I__15897 (
            .O(N__67668),
            .I(\c0.n26_adj_4530 ));
    InMux I__15896 (
            .O(N__67665),
            .I(N__67661));
    InMux I__15895 (
            .O(N__67664),
            .I(N__67658));
    LocalMux I__15894 (
            .O(N__67661),
            .I(N__67652));
    LocalMux I__15893 (
            .O(N__67658),
            .I(N__67652));
    InMux I__15892 (
            .O(N__67657),
            .I(N__67649));
    Span4Mux_v I__15891 (
            .O(N__67652),
            .I(N__67645));
    LocalMux I__15890 (
            .O(N__67649),
            .I(N__67641));
    InMux I__15889 (
            .O(N__67648),
            .I(N__67637));
    Span4Mux_h I__15888 (
            .O(N__67645),
            .I(N__67634));
    InMux I__15887 (
            .O(N__67644),
            .I(N__67631));
    Span4Mux_h I__15886 (
            .O(N__67641),
            .I(N__67628));
    InMux I__15885 (
            .O(N__67640),
            .I(N__67625));
    LocalMux I__15884 (
            .O(N__67637),
            .I(N__67622));
    Span4Mux_v I__15883 (
            .O(N__67634),
            .I(N__67617));
    LocalMux I__15882 (
            .O(N__67631),
            .I(N__67614));
    Span4Mux_h I__15881 (
            .O(N__67628),
            .I(N__67607));
    LocalMux I__15880 (
            .O(N__67625),
            .I(N__67607));
    Span4Mux_h I__15879 (
            .O(N__67622),
            .I(N__67607));
    InMux I__15878 (
            .O(N__67621),
            .I(N__67602));
    InMux I__15877 (
            .O(N__67620),
            .I(N__67602));
    Odrv4 I__15876 (
            .O(N__67617),
            .I(n22103));
    Odrv4 I__15875 (
            .O(N__67614),
            .I(n22103));
    Odrv4 I__15874 (
            .O(N__67607),
            .I(n22103));
    LocalMux I__15873 (
            .O(N__67602),
            .I(n22103));
    InMux I__15872 (
            .O(N__67593),
            .I(N__67588));
    InMux I__15871 (
            .O(N__67592),
            .I(N__67585));
    InMux I__15870 (
            .O(N__67591),
            .I(N__67582));
    LocalMux I__15869 (
            .O(N__67588),
            .I(N__67577));
    LocalMux I__15868 (
            .O(N__67585),
            .I(N__67577));
    LocalMux I__15867 (
            .O(N__67582),
            .I(N__67574));
    Span4Mux_v I__15866 (
            .O(N__67577),
            .I(N__67571));
    Odrv4 I__15865 (
            .O(N__67574),
            .I(\c0.n22632 ));
    Odrv4 I__15864 (
            .O(N__67571),
            .I(\c0.n22632 ));
    CascadeMux I__15863 (
            .O(N__67566),
            .I(\c0.n22632_cascade_ ));
    InMux I__15862 (
            .O(N__67563),
            .I(N__67560));
    LocalMux I__15861 (
            .O(N__67560),
            .I(N__67556));
    InMux I__15860 (
            .O(N__67559),
            .I(N__67553));
    Span4Mux_v I__15859 (
            .O(N__67556),
            .I(N__67544));
    LocalMux I__15858 (
            .O(N__67553),
            .I(N__67544));
    InMux I__15857 (
            .O(N__67552),
            .I(N__67539));
    InMux I__15856 (
            .O(N__67551),
            .I(N__67539));
    InMux I__15855 (
            .O(N__67550),
            .I(N__67536));
    InMux I__15854 (
            .O(N__67549),
            .I(N__67533));
    Span4Mux_h I__15853 (
            .O(N__67544),
            .I(N__67529));
    LocalMux I__15852 (
            .O(N__67539),
            .I(N__67522));
    LocalMux I__15851 (
            .O(N__67536),
            .I(N__67522));
    LocalMux I__15850 (
            .O(N__67533),
            .I(N__67522));
    InMux I__15849 (
            .O(N__67532),
            .I(N__67519));
    Span4Mux_h I__15848 (
            .O(N__67529),
            .I(N__67516));
    Span12Mux_h I__15847 (
            .O(N__67522),
            .I(N__67513));
    LocalMux I__15846 (
            .O(N__67519),
            .I(\c0.data_in_frame_24_2 ));
    Odrv4 I__15845 (
            .O(N__67516),
            .I(\c0.data_in_frame_24_2 ));
    Odrv12 I__15844 (
            .O(N__67513),
            .I(\c0.data_in_frame_24_2 ));
    InMux I__15843 (
            .O(N__67506),
            .I(N__67502));
    InMux I__15842 (
            .O(N__67505),
            .I(N__67496));
    LocalMux I__15841 (
            .O(N__67502),
            .I(N__67493));
    InMux I__15840 (
            .O(N__67501),
            .I(N__67488));
    InMux I__15839 (
            .O(N__67500),
            .I(N__67483));
    InMux I__15838 (
            .O(N__67499),
            .I(N__67483));
    LocalMux I__15837 (
            .O(N__67496),
            .I(N__67480));
    Span4Mux_h I__15836 (
            .O(N__67493),
            .I(N__67477));
    InMux I__15835 (
            .O(N__67492),
            .I(N__67472));
    InMux I__15834 (
            .O(N__67491),
            .I(N__67472));
    LocalMux I__15833 (
            .O(N__67488),
            .I(\c0.n21316 ));
    LocalMux I__15832 (
            .O(N__67483),
            .I(\c0.n21316 ));
    Odrv12 I__15831 (
            .O(N__67480),
            .I(\c0.n21316 ));
    Odrv4 I__15830 (
            .O(N__67477),
            .I(\c0.n21316 ));
    LocalMux I__15829 (
            .O(N__67472),
            .I(\c0.n21316 ));
    InMux I__15828 (
            .O(N__67461),
            .I(N__67458));
    LocalMux I__15827 (
            .O(N__67458),
            .I(\c0.n39_adj_4487 ));
    CascadeMux I__15826 (
            .O(N__67455),
            .I(\c0.n30_adj_4489_cascade_ ));
    InMux I__15825 (
            .O(N__67452),
            .I(N__67449));
    LocalMux I__15824 (
            .O(N__67449),
            .I(\c0.n23209 ));
    CascadeMux I__15823 (
            .O(N__67446),
            .I(\c0.n45_adj_4490_cascade_ ));
    InMux I__15822 (
            .O(N__67443),
            .I(N__67440));
    LocalMux I__15821 (
            .O(N__67440),
            .I(N__67437));
    Odrv4 I__15820 (
            .O(N__67437),
            .I(\c0.n44_adj_4501 ));
    InMux I__15819 (
            .O(N__67434),
            .I(N__67431));
    LocalMux I__15818 (
            .O(N__67431),
            .I(N__67428));
    Span4Mux_h I__15817 (
            .O(N__67428),
            .I(N__67425));
    Odrv4 I__15816 (
            .O(N__67425),
            .I(\c0.n11_adj_4505 ));
    CascadeMux I__15815 (
            .O(N__67422),
            .I(\c0.n48_adj_4503_cascade_ ));
    InMux I__15814 (
            .O(N__67419),
            .I(N__67416));
    LocalMux I__15813 (
            .O(N__67416),
            .I(N__67412));
    CascadeMux I__15812 (
            .O(N__67415),
            .I(N__67409));
    Span4Mux_h I__15811 (
            .O(N__67412),
            .I(N__67406));
    InMux I__15810 (
            .O(N__67409),
            .I(N__67403));
    Odrv4 I__15809 (
            .O(N__67406),
            .I(\c0.n28_adj_4504 ));
    LocalMux I__15808 (
            .O(N__67403),
            .I(\c0.n28_adj_4504 ));
    InMux I__15807 (
            .O(N__67398),
            .I(N__67395));
    LocalMux I__15806 (
            .O(N__67395),
            .I(N__67392));
    Span4Mux_v I__15805 (
            .O(N__67392),
            .I(N__67389));
    Odrv4 I__15804 (
            .O(N__67389),
            .I(\c0.n24573 ));
    InMux I__15803 (
            .O(N__67386),
            .I(N__67383));
    LocalMux I__15802 (
            .O(N__67383),
            .I(\c0.n41_adj_4488 ));
    InMux I__15801 (
            .O(N__67380),
            .I(N__67377));
    LocalMux I__15800 (
            .O(N__67377),
            .I(N__67373));
    InMux I__15799 (
            .O(N__67376),
            .I(N__67370));
    Span4Mux_v I__15798 (
            .O(N__67373),
            .I(N__67365));
    LocalMux I__15797 (
            .O(N__67370),
            .I(N__67365));
    Odrv4 I__15796 (
            .O(N__67365),
            .I(\c0.n17_adj_4354 ));
    InMux I__15795 (
            .O(N__67362),
            .I(N__67358));
    InMux I__15794 (
            .O(N__67361),
            .I(N__67355));
    LocalMux I__15793 (
            .O(N__67358),
            .I(N__67352));
    LocalMux I__15792 (
            .O(N__67355),
            .I(N__67348));
    Span4Mux_h I__15791 (
            .O(N__67352),
            .I(N__67345));
    InMux I__15790 (
            .O(N__67351),
            .I(N__67342));
    Odrv4 I__15789 (
            .O(N__67348),
            .I(\c0.n28_adj_4343 ));
    Odrv4 I__15788 (
            .O(N__67345),
            .I(\c0.n28_adj_4343 ));
    LocalMux I__15787 (
            .O(N__67342),
            .I(\c0.n28_adj_4343 ));
    InMux I__15786 (
            .O(N__67335),
            .I(N__67332));
    LocalMux I__15785 (
            .O(N__67332),
            .I(\c0.n27_adj_4502 ));
    CascadeMux I__15784 (
            .O(N__67329),
            .I(N__67324));
    InMux I__15783 (
            .O(N__67328),
            .I(N__67321));
    CascadeMux I__15782 (
            .O(N__67327),
            .I(N__67318));
    InMux I__15781 (
            .O(N__67324),
            .I(N__67315));
    LocalMux I__15780 (
            .O(N__67321),
            .I(N__67310));
    InMux I__15779 (
            .O(N__67318),
            .I(N__67307));
    LocalMux I__15778 (
            .O(N__67315),
            .I(N__67304));
    InMux I__15777 (
            .O(N__67314),
            .I(N__67301));
    InMux I__15776 (
            .O(N__67313),
            .I(N__67298));
    Span4Mux_h I__15775 (
            .O(N__67310),
            .I(N__67287));
    LocalMux I__15774 (
            .O(N__67307),
            .I(N__67287));
    Span4Mux_h I__15773 (
            .O(N__67304),
            .I(N__67287));
    LocalMux I__15772 (
            .O(N__67301),
            .I(N__67287));
    LocalMux I__15771 (
            .O(N__67298),
            .I(N__67284));
    InMux I__15770 (
            .O(N__67297),
            .I(N__67281));
    InMux I__15769 (
            .O(N__67296),
            .I(N__67278));
    Span4Mux_h I__15768 (
            .O(N__67287),
            .I(N__67275));
    Span12Mux_h I__15767 (
            .O(N__67284),
            .I(N__67272));
    LocalMux I__15766 (
            .O(N__67281),
            .I(N__67269));
    LocalMux I__15765 (
            .O(N__67278),
            .I(\c0.data_in_frame_26_7 ));
    Odrv4 I__15764 (
            .O(N__67275),
            .I(\c0.data_in_frame_26_7 ));
    Odrv12 I__15763 (
            .O(N__67272),
            .I(\c0.data_in_frame_26_7 ));
    Odrv12 I__15762 (
            .O(N__67269),
            .I(\c0.data_in_frame_26_7 ));
    InMux I__15761 (
            .O(N__67260),
            .I(N__67257));
    LocalMux I__15760 (
            .O(N__67257),
            .I(N__67252));
    InMux I__15759 (
            .O(N__67256),
            .I(N__67243));
    InMux I__15758 (
            .O(N__67255),
            .I(N__67243));
    Span4Mux_v I__15757 (
            .O(N__67252),
            .I(N__67240));
    InMux I__15756 (
            .O(N__67251),
            .I(N__67235));
    InMux I__15755 (
            .O(N__67250),
            .I(N__67235));
    InMux I__15754 (
            .O(N__67249),
            .I(N__67230));
    InMux I__15753 (
            .O(N__67248),
            .I(N__67230));
    LocalMux I__15752 (
            .O(N__67243),
            .I(N__67223));
    Sp12to4 I__15751 (
            .O(N__67240),
            .I(N__67223));
    LocalMux I__15750 (
            .O(N__67235),
            .I(N__67223));
    LocalMux I__15749 (
            .O(N__67230),
            .I(\c0.data_in_frame_24_4 ));
    Odrv12 I__15748 (
            .O(N__67223),
            .I(\c0.data_in_frame_24_4 ));
    CascadeMux I__15747 (
            .O(N__67218),
            .I(N__67215));
    InMux I__15746 (
            .O(N__67215),
            .I(N__67209));
    InMux I__15745 (
            .O(N__67214),
            .I(N__67204));
    InMux I__15744 (
            .O(N__67213),
            .I(N__67204));
    InMux I__15743 (
            .O(N__67212),
            .I(N__67201));
    LocalMux I__15742 (
            .O(N__67209),
            .I(data_in_frame_21_6));
    LocalMux I__15741 (
            .O(N__67204),
            .I(data_in_frame_21_6));
    LocalMux I__15740 (
            .O(N__67201),
            .I(data_in_frame_21_6));
    InMux I__15739 (
            .O(N__67194),
            .I(N__67190));
    InMux I__15738 (
            .O(N__67193),
            .I(N__67187));
    LocalMux I__15737 (
            .O(N__67190),
            .I(N__67184));
    LocalMux I__15736 (
            .O(N__67187),
            .I(N__67181));
    Span4Mux_v I__15735 (
            .O(N__67184),
            .I(N__67177));
    Span4Mux_v I__15734 (
            .O(N__67181),
            .I(N__67174));
    InMux I__15733 (
            .O(N__67180),
            .I(N__67171));
    Odrv4 I__15732 (
            .O(N__67177),
            .I(\c0.n21301 ));
    Odrv4 I__15731 (
            .O(N__67174),
            .I(\c0.n21301 ));
    LocalMux I__15730 (
            .O(N__67171),
            .I(\c0.n21301 ));
    InMux I__15729 (
            .O(N__67164),
            .I(N__67160));
    InMux I__15728 (
            .O(N__67163),
            .I(N__67157));
    LocalMux I__15727 (
            .O(N__67160),
            .I(\c0.n23_adj_4582 ));
    LocalMux I__15726 (
            .O(N__67157),
            .I(\c0.n23_adj_4582 ));
    CascadeMux I__15725 (
            .O(N__67152),
            .I(N__67144));
    InMux I__15724 (
            .O(N__67151),
            .I(N__67141));
    CascadeMux I__15723 (
            .O(N__67150),
            .I(N__67137));
    InMux I__15722 (
            .O(N__67149),
            .I(N__67128));
    InMux I__15721 (
            .O(N__67148),
            .I(N__67128));
    InMux I__15720 (
            .O(N__67147),
            .I(N__67128));
    InMux I__15719 (
            .O(N__67144),
            .I(N__67128));
    LocalMux I__15718 (
            .O(N__67141),
            .I(N__67125));
    InMux I__15717 (
            .O(N__67140),
            .I(N__67122));
    InMux I__15716 (
            .O(N__67137),
            .I(N__67118));
    LocalMux I__15715 (
            .O(N__67128),
            .I(N__67115));
    Span4Mux_v I__15714 (
            .O(N__67125),
            .I(N__67112));
    LocalMux I__15713 (
            .O(N__67122),
            .I(N__67109));
    InMux I__15712 (
            .O(N__67121),
            .I(N__67106));
    LocalMux I__15711 (
            .O(N__67118),
            .I(N__67099));
    Span4Mux_v I__15710 (
            .O(N__67115),
            .I(N__67099));
    Span4Mux_h I__15709 (
            .O(N__67112),
            .I(N__67099));
    Span4Mux_v I__15708 (
            .O(N__67109),
            .I(N__67096));
    LocalMux I__15707 (
            .O(N__67106),
            .I(\c0.data_in_frame_24_6 ));
    Odrv4 I__15706 (
            .O(N__67099),
            .I(\c0.data_in_frame_24_6 ));
    Odrv4 I__15705 (
            .O(N__67096),
            .I(\c0.data_in_frame_24_6 ));
    InMux I__15704 (
            .O(N__67089),
            .I(N__67086));
    LocalMux I__15703 (
            .O(N__67086),
            .I(N__67083));
    Span4Mux_h I__15702 (
            .O(N__67083),
            .I(N__67079));
    InMux I__15701 (
            .O(N__67082),
            .I(N__67076));
    Odrv4 I__15700 (
            .O(N__67079),
            .I(\c0.n22495 ));
    LocalMux I__15699 (
            .O(N__67076),
            .I(\c0.n22495 ));
    CascadeMux I__15698 (
            .O(N__67071),
            .I(N__67067));
    InMux I__15697 (
            .O(N__67070),
            .I(N__67064));
    InMux I__15696 (
            .O(N__67067),
            .I(N__67061));
    LocalMux I__15695 (
            .O(N__67064),
            .I(\c0.data_in_frame_20_1 ));
    LocalMux I__15694 (
            .O(N__67061),
            .I(\c0.data_in_frame_20_1 ));
    InMux I__15693 (
            .O(N__67056),
            .I(N__67052));
    InMux I__15692 (
            .O(N__67055),
            .I(N__67049));
    LocalMux I__15691 (
            .O(N__67052),
            .I(N__67046));
    LocalMux I__15690 (
            .O(N__67049),
            .I(N__67043));
    Odrv4 I__15689 (
            .O(N__67046),
            .I(\c0.n58_adj_4355 ));
    Odrv4 I__15688 (
            .O(N__67043),
            .I(\c0.n58_adj_4355 ));
    InMux I__15687 (
            .O(N__67038),
            .I(N__67034));
    InMux I__15686 (
            .O(N__67037),
            .I(N__67030));
    LocalMux I__15685 (
            .O(N__67034),
            .I(N__67027));
    InMux I__15684 (
            .O(N__67033),
            .I(N__67024));
    LocalMux I__15683 (
            .O(N__67030),
            .I(N__67021));
    Span4Mux_h I__15682 (
            .O(N__67027),
            .I(N__67018));
    LocalMux I__15681 (
            .O(N__67024),
            .I(N__67015));
    Span4Mux_v I__15680 (
            .O(N__67021),
            .I(N__67012));
    Odrv4 I__15679 (
            .O(N__67018),
            .I(\c0.n59_adj_4351 ));
    Odrv12 I__15678 (
            .O(N__67015),
            .I(\c0.n59_adj_4351 ));
    Odrv4 I__15677 (
            .O(N__67012),
            .I(\c0.n59_adj_4351 ));
    InMux I__15676 (
            .O(N__67005),
            .I(N__67002));
    LocalMux I__15675 (
            .O(N__67002),
            .I(N__66999));
    Span4Mux_v I__15674 (
            .O(N__66999),
            .I(N__66995));
    InMux I__15673 (
            .O(N__66998),
            .I(N__66992));
    Odrv4 I__15672 (
            .O(N__66995),
            .I(\c0.n28_adj_4363 ));
    LocalMux I__15671 (
            .O(N__66992),
            .I(\c0.n28_adj_4363 ));
    InMux I__15670 (
            .O(N__66987),
            .I(N__66979));
    InMux I__15669 (
            .O(N__66986),
            .I(N__66979));
    InMux I__15668 (
            .O(N__66985),
            .I(N__66976));
    InMux I__15667 (
            .O(N__66984),
            .I(N__66973));
    LocalMux I__15666 (
            .O(N__66979),
            .I(N__66970));
    LocalMux I__15665 (
            .O(N__66976),
            .I(N__66965));
    LocalMux I__15664 (
            .O(N__66973),
            .I(N__66965));
    Span4Mux_v I__15663 (
            .O(N__66970),
            .I(N__66962));
    Odrv4 I__15662 (
            .O(N__66965),
            .I(\c0.n23691 ));
    Odrv4 I__15661 (
            .O(N__66962),
            .I(\c0.n23691 ));
    CascadeMux I__15660 (
            .O(N__66957),
            .I(N__66954));
    InMux I__15659 (
            .O(N__66954),
            .I(N__66951));
    LocalMux I__15658 (
            .O(N__66951),
            .I(N__66947));
    InMux I__15657 (
            .O(N__66950),
            .I(N__66944));
    Span4Mux_h I__15656 (
            .O(N__66947),
            .I(N__66939));
    LocalMux I__15655 (
            .O(N__66944),
            .I(N__66939));
    Span4Mux_h I__15654 (
            .O(N__66939),
            .I(N__66936));
    Span4Mux_h I__15653 (
            .O(N__66936),
            .I(N__66933));
    Odrv4 I__15652 (
            .O(N__66933),
            .I(\c0.n22577 ));
    InMux I__15651 (
            .O(N__66930),
            .I(N__66926));
    InMux I__15650 (
            .O(N__66929),
            .I(N__66923));
    LocalMux I__15649 (
            .O(N__66926),
            .I(N__66920));
    LocalMux I__15648 (
            .O(N__66923),
            .I(N__66916));
    Span4Mux_h I__15647 (
            .O(N__66920),
            .I(N__66913));
    InMux I__15646 (
            .O(N__66919),
            .I(N__66910));
    Odrv12 I__15645 (
            .O(N__66916),
            .I(\c0.n21414 ));
    Odrv4 I__15644 (
            .O(N__66913),
            .I(\c0.n21414 ));
    LocalMux I__15643 (
            .O(N__66910),
            .I(\c0.n21414 ));
    CascadeMux I__15642 (
            .O(N__66903),
            .I(\c0.n10_adj_4524_cascade_ ));
    CascadeMux I__15641 (
            .O(N__66900),
            .I(N__66894));
    InMux I__15640 (
            .O(N__66899),
            .I(N__66890));
    InMux I__15639 (
            .O(N__66898),
            .I(N__66887));
    InMux I__15638 (
            .O(N__66897),
            .I(N__66884));
    InMux I__15637 (
            .O(N__66894),
            .I(N__66881));
    InMux I__15636 (
            .O(N__66893),
            .I(N__66878));
    LocalMux I__15635 (
            .O(N__66890),
            .I(N__66875));
    LocalMux I__15634 (
            .O(N__66887),
            .I(N__66872));
    LocalMux I__15633 (
            .O(N__66884),
            .I(N__66864));
    LocalMux I__15632 (
            .O(N__66881),
            .I(N__66864));
    LocalMux I__15631 (
            .O(N__66878),
            .I(N__66864));
    Span4Mux_v I__15630 (
            .O(N__66875),
            .I(N__66858));
    Span4Mux_h I__15629 (
            .O(N__66872),
            .I(N__66858));
    InMux I__15628 (
            .O(N__66871),
            .I(N__66855));
    Span4Mux_v I__15627 (
            .O(N__66864),
            .I(N__66852));
    InMux I__15626 (
            .O(N__66863),
            .I(N__66849));
    Span4Mux_v I__15625 (
            .O(N__66858),
            .I(N__66846));
    LocalMux I__15624 (
            .O(N__66855),
            .I(N__66841));
    Span4Mux_h I__15623 (
            .O(N__66852),
            .I(N__66841));
    LocalMux I__15622 (
            .O(N__66849),
            .I(N__66838));
    Odrv4 I__15621 (
            .O(N__66846),
            .I(\c0.n13797 ));
    Odrv4 I__15620 (
            .O(N__66841),
            .I(\c0.n13797 ));
    Odrv4 I__15619 (
            .O(N__66838),
            .I(\c0.n13797 ));
    InMux I__15618 (
            .O(N__66831),
            .I(N__66828));
    LocalMux I__15617 (
            .O(N__66828),
            .I(N__66824));
    InMux I__15616 (
            .O(N__66827),
            .I(N__66821));
    Span4Mux_v I__15615 (
            .O(N__66824),
            .I(N__66818));
    LocalMux I__15614 (
            .O(N__66821),
            .I(\c0.n24576 ));
    Odrv4 I__15613 (
            .O(N__66818),
            .I(\c0.n24576 ));
    InMux I__15612 (
            .O(N__66813),
            .I(N__66808));
    InMux I__15611 (
            .O(N__66812),
            .I(N__66802));
    InMux I__15610 (
            .O(N__66811),
            .I(N__66802));
    LocalMux I__15609 (
            .O(N__66808),
            .I(N__66799));
    CascadeMux I__15608 (
            .O(N__66807),
            .I(N__66796));
    LocalMux I__15607 (
            .O(N__66802),
            .I(N__66793));
    Span4Mux_h I__15606 (
            .O(N__66799),
            .I(N__66790));
    InMux I__15605 (
            .O(N__66796),
            .I(N__66787));
    Span4Mux_h I__15604 (
            .O(N__66793),
            .I(N__66784));
    Span4Mux_h I__15603 (
            .O(N__66790),
            .I(N__66781));
    LocalMux I__15602 (
            .O(N__66787),
            .I(N__66776));
    Span4Mux_h I__15601 (
            .O(N__66784),
            .I(N__66776));
    Odrv4 I__15600 (
            .O(N__66781),
            .I(\c0.data_in_frame_26_2 ));
    Odrv4 I__15599 (
            .O(N__66776),
            .I(\c0.data_in_frame_26_2 ));
    CascadeMux I__15598 (
            .O(N__66771),
            .I(\c0.n24576_cascade_ ));
    InMux I__15597 (
            .O(N__66768),
            .I(N__66765));
    LocalMux I__15596 (
            .O(N__66765),
            .I(N__66762));
    Span4Mux_v I__15595 (
            .O(N__66762),
            .I(N__66759));
    Odrv4 I__15594 (
            .O(N__66759),
            .I(\c0.n14_adj_4519 ));
    InMux I__15593 (
            .O(N__66756),
            .I(N__66753));
    LocalMux I__15592 (
            .O(N__66753),
            .I(N__66747));
    InMux I__15591 (
            .O(N__66752),
            .I(N__66743));
    InMux I__15590 (
            .O(N__66751),
            .I(N__66740));
    InMux I__15589 (
            .O(N__66750),
            .I(N__66737));
    Span4Mux_h I__15588 (
            .O(N__66747),
            .I(N__66734));
    InMux I__15587 (
            .O(N__66746),
            .I(N__66731));
    LocalMux I__15586 (
            .O(N__66743),
            .I(N__66724));
    LocalMux I__15585 (
            .O(N__66740),
            .I(N__66724));
    LocalMux I__15584 (
            .O(N__66737),
            .I(N__66724));
    Span4Mux_h I__15583 (
            .O(N__66734),
            .I(N__66721));
    LocalMux I__15582 (
            .O(N__66731),
            .I(data_in_frame_21_4));
    Odrv12 I__15581 (
            .O(N__66724),
            .I(data_in_frame_21_4));
    Odrv4 I__15580 (
            .O(N__66721),
            .I(data_in_frame_21_4));
    InMux I__15579 (
            .O(N__66714),
            .I(N__66711));
    LocalMux I__15578 (
            .O(N__66711),
            .I(N__66706));
    InMux I__15577 (
            .O(N__66710),
            .I(N__66703));
    InMux I__15576 (
            .O(N__66709),
            .I(N__66700));
    Span4Mux_h I__15575 (
            .O(N__66706),
            .I(N__66697));
    LocalMux I__15574 (
            .O(N__66703),
            .I(N__66694));
    LocalMux I__15573 (
            .O(N__66700),
            .I(\c0.n23733 ));
    Odrv4 I__15572 (
            .O(N__66697),
            .I(\c0.n23733 ));
    Odrv4 I__15571 (
            .O(N__66694),
            .I(\c0.n23733 ));
    InMux I__15570 (
            .O(N__66687),
            .I(N__66684));
    LocalMux I__15569 (
            .O(N__66684),
            .I(\c0.n22686 ));
    InMux I__15568 (
            .O(N__66681),
            .I(N__66678));
    LocalMux I__15567 (
            .O(N__66678),
            .I(N__66675));
    Span4Mux_v I__15566 (
            .O(N__66675),
            .I(N__66672));
    Odrv4 I__15565 (
            .O(N__66672),
            .I(\c0.n5_adj_4472 ));
    CascadeMux I__15564 (
            .O(N__66669),
            .I(\c0.n22686_cascade_ ));
    InMux I__15563 (
            .O(N__66666),
            .I(N__66663));
    LocalMux I__15562 (
            .O(N__66663),
            .I(N__66658));
    InMux I__15561 (
            .O(N__66662),
            .I(N__66655));
    InMux I__15560 (
            .O(N__66661),
            .I(N__66651));
    Span4Mux_v I__15559 (
            .O(N__66658),
            .I(N__66647));
    LocalMux I__15558 (
            .O(N__66655),
            .I(N__66644));
    InMux I__15557 (
            .O(N__66654),
            .I(N__66641));
    LocalMux I__15556 (
            .O(N__66651),
            .I(N__66638));
    InMux I__15555 (
            .O(N__66650),
            .I(N__66634));
    Span4Mux_h I__15554 (
            .O(N__66647),
            .I(N__66629));
    Span4Mux_v I__15553 (
            .O(N__66644),
            .I(N__66629));
    LocalMux I__15552 (
            .O(N__66641),
            .I(N__66624));
    Span4Mux_h I__15551 (
            .O(N__66638),
            .I(N__66624));
    InMux I__15550 (
            .O(N__66637),
            .I(N__66621));
    LocalMux I__15549 (
            .O(N__66634),
            .I(\c0.data_in_frame_18_3 ));
    Odrv4 I__15548 (
            .O(N__66629),
            .I(\c0.data_in_frame_18_3 ));
    Odrv4 I__15547 (
            .O(N__66624),
            .I(\c0.data_in_frame_18_3 ));
    LocalMux I__15546 (
            .O(N__66621),
            .I(\c0.data_in_frame_18_3 ));
    InMux I__15545 (
            .O(N__66612),
            .I(N__66609));
    LocalMux I__15544 (
            .O(N__66609),
            .I(N__66605));
    InMux I__15543 (
            .O(N__66608),
            .I(N__66602));
    Odrv4 I__15542 (
            .O(N__66605),
            .I(\c0.n5_adj_4335 ));
    LocalMux I__15541 (
            .O(N__66602),
            .I(\c0.n5_adj_4335 ));
    InMux I__15540 (
            .O(N__66597),
            .I(N__66594));
    LocalMux I__15539 (
            .O(N__66594),
            .I(N__66590));
    InMux I__15538 (
            .O(N__66593),
            .I(N__66587));
    Span4Mux_h I__15537 (
            .O(N__66590),
            .I(N__66584));
    LocalMux I__15536 (
            .O(N__66587),
            .I(\c0.n4_adj_4568 ));
    Odrv4 I__15535 (
            .O(N__66584),
            .I(\c0.n4_adj_4568 ));
    InMux I__15534 (
            .O(N__66579),
            .I(N__66576));
    LocalMux I__15533 (
            .O(N__66576),
            .I(N__66573));
    Odrv12 I__15532 (
            .O(N__66573),
            .I(\c0.n15_adj_4569 ));
    InMux I__15531 (
            .O(N__66570),
            .I(N__66566));
    InMux I__15530 (
            .O(N__66569),
            .I(N__66562));
    LocalMux I__15529 (
            .O(N__66566),
            .I(N__66559));
    InMux I__15528 (
            .O(N__66565),
            .I(N__66556));
    LocalMux I__15527 (
            .O(N__66562),
            .I(N__66553));
    Span4Mux_h I__15526 (
            .O(N__66559),
            .I(N__66549));
    LocalMux I__15525 (
            .O(N__66556),
            .I(N__66546));
    Span4Mux_v I__15524 (
            .O(N__66553),
            .I(N__66543));
    InMux I__15523 (
            .O(N__66552),
            .I(N__66540));
    Span4Mux_h I__15522 (
            .O(N__66549),
            .I(N__66537));
    Span4Mux_v I__15521 (
            .O(N__66546),
            .I(N__66532));
    Span4Mux_h I__15520 (
            .O(N__66543),
            .I(N__66532));
    LocalMux I__15519 (
            .O(N__66540),
            .I(\c0.data_in_frame_18_7 ));
    Odrv4 I__15518 (
            .O(N__66537),
            .I(\c0.data_in_frame_18_7 ));
    Odrv4 I__15517 (
            .O(N__66532),
            .I(\c0.data_in_frame_18_7 ));
    InMux I__15516 (
            .O(N__66525),
            .I(N__66522));
    LocalMux I__15515 (
            .O(N__66522),
            .I(N__66518));
    CascadeMux I__15514 (
            .O(N__66521),
            .I(N__66514));
    Span12Mux_v I__15513 (
            .O(N__66518),
            .I(N__66511));
    InMux I__15512 (
            .O(N__66517),
            .I(N__66506));
    InMux I__15511 (
            .O(N__66514),
            .I(N__66506));
    Odrv12 I__15510 (
            .O(N__66511),
            .I(data_in_frame_22_5));
    LocalMux I__15509 (
            .O(N__66506),
            .I(data_in_frame_22_5));
    CascadeMux I__15508 (
            .O(N__66501),
            .I(N__66497));
    CascadeMux I__15507 (
            .O(N__66500),
            .I(N__66492));
    InMux I__15506 (
            .O(N__66497),
            .I(N__66487));
    InMux I__15505 (
            .O(N__66496),
            .I(N__66487));
    InMux I__15504 (
            .O(N__66495),
            .I(N__66484));
    InMux I__15503 (
            .O(N__66492),
            .I(N__66481));
    LocalMux I__15502 (
            .O(N__66487),
            .I(N__66478));
    LocalMux I__15501 (
            .O(N__66484),
            .I(N__66475));
    LocalMux I__15500 (
            .O(N__66481),
            .I(N__66470));
    Span4Mux_h I__15499 (
            .O(N__66478),
            .I(N__66470));
    Odrv4 I__15498 (
            .O(N__66475),
            .I(\c0.data_in_frame_17_5 ));
    Odrv4 I__15497 (
            .O(N__66470),
            .I(\c0.data_in_frame_17_5 ));
    InMux I__15496 (
            .O(N__66465),
            .I(N__66461));
    InMux I__15495 (
            .O(N__66464),
            .I(N__66458));
    LocalMux I__15494 (
            .O(N__66461),
            .I(N__66455));
    LocalMux I__15493 (
            .O(N__66458),
            .I(N__66452));
    Span4Mux_v I__15492 (
            .O(N__66455),
            .I(N__66447));
    Span4Mux_h I__15491 (
            .O(N__66452),
            .I(N__66447));
    Odrv4 I__15490 (
            .O(N__66447),
            .I(\c0.n22748 ));
    CascadeMux I__15489 (
            .O(N__66444),
            .I(\c0.n14_adj_4623_cascade_ ));
    InMux I__15488 (
            .O(N__66441),
            .I(N__66438));
    LocalMux I__15487 (
            .O(N__66438),
            .I(\c0.n15_adj_4624 ));
    InMux I__15486 (
            .O(N__66435),
            .I(N__66432));
    LocalMux I__15485 (
            .O(N__66432),
            .I(N__66427));
    InMux I__15484 (
            .O(N__66431),
            .I(N__66422));
    InMux I__15483 (
            .O(N__66430),
            .I(N__66419));
    Span4Mux_h I__15482 (
            .O(N__66427),
            .I(N__66416));
    InMux I__15481 (
            .O(N__66426),
            .I(N__66411));
    InMux I__15480 (
            .O(N__66425),
            .I(N__66411));
    LocalMux I__15479 (
            .O(N__66422),
            .I(N__66408));
    LocalMux I__15478 (
            .O(N__66419),
            .I(N__66403));
    Span4Mux_h I__15477 (
            .O(N__66416),
            .I(N__66403));
    LocalMux I__15476 (
            .O(N__66411),
            .I(data_in_frame_21_1));
    Odrv4 I__15475 (
            .O(N__66408),
            .I(data_in_frame_21_1));
    Odrv4 I__15474 (
            .O(N__66403),
            .I(data_in_frame_21_1));
    CascadeMux I__15473 (
            .O(N__66396),
            .I(\c0.n13963_cascade_ ));
    InMux I__15472 (
            .O(N__66393),
            .I(N__66389));
    InMux I__15471 (
            .O(N__66392),
            .I(N__66386));
    LocalMux I__15470 (
            .O(N__66389),
            .I(N__66381));
    LocalMux I__15469 (
            .O(N__66386),
            .I(N__66381));
    Span4Mux_v I__15468 (
            .O(N__66381),
            .I(N__66378));
    Odrv4 I__15467 (
            .O(N__66378),
            .I(\c0.n22508 ));
    InMux I__15466 (
            .O(N__66375),
            .I(N__66372));
    LocalMux I__15465 (
            .O(N__66372),
            .I(\c0.n40_adj_4342 ));
    InMux I__15464 (
            .O(N__66369),
            .I(N__66366));
    LocalMux I__15463 (
            .O(N__66366),
            .I(N__66361));
    InMux I__15462 (
            .O(N__66365),
            .I(N__66356));
    InMux I__15461 (
            .O(N__66364),
            .I(N__66356));
    Span12Mux_h I__15460 (
            .O(N__66361),
            .I(N__66352));
    LocalMux I__15459 (
            .O(N__66356),
            .I(N__66349));
    InMux I__15458 (
            .O(N__66355),
            .I(N__66346));
    Odrv12 I__15457 (
            .O(N__66352),
            .I(\c0.n13604 ));
    Odrv4 I__15456 (
            .O(N__66349),
            .I(\c0.n13604 ));
    LocalMux I__15455 (
            .O(N__66346),
            .I(\c0.n13604 ));
    CascadeMux I__15454 (
            .O(N__66339),
            .I(\c0.n7_adj_4251_cascade_ ));
    InMux I__15453 (
            .O(N__66336),
            .I(N__66330));
    InMux I__15452 (
            .O(N__66335),
            .I(N__66327));
    InMux I__15451 (
            .O(N__66334),
            .I(N__66322));
    InMux I__15450 (
            .O(N__66333),
            .I(N__66322));
    LocalMux I__15449 (
            .O(N__66330),
            .I(\c0.n23224 ));
    LocalMux I__15448 (
            .O(N__66327),
            .I(\c0.n23224 ));
    LocalMux I__15447 (
            .O(N__66322),
            .I(\c0.n23224 ));
    InMux I__15446 (
            .O(N__66315),
            .I(N__66312));
    LocalMux I__15445 (
            .O(N__66312),
            .I(\c0.n7_adj_4251 ));
    InMux I__15444 (
            .O(N__66309),
            .I(N__66306));
    LocalMux I__15443 (
            .O(N__66306),
            .I(N__66303));
    Span4Mux_h I__15442 (
            .O(N__66303),
            .I(N__66299));
    InMux I__15441 (
            .O(N__66302),
            .I(N__66296));
    Span4Mux_h I__15440 (
            .O(N__66299),
            .I(N__66293));
    LocalMux I__15439 (
            .O(N__66296),
            .I(data_in_frame_22_7));
    Odrv4 I__15438 (
            .O(N__66293),
            .I(data_in_frame_22_7));
    InMux I__15437 (
            .O(N__66288),
            .I(N__66285));
    LocalMux I__15436 (
            .O(N__66285),
            .I(N__66282));
    Span4Mux_v I__15435 (
            .O(N__66282),
            .I(N__66279));
    Sp12to4 I__15434 (
            .O(N__66279),
            .I(N__66276));
    Odrv12 I__15433 (
            .O(N__66276),
            .I(\c0.n22825 ));
    CascadeMux I__15432 (
            .O(N__66273),
            .I(N__66268));
    InMux I__15431 (
            .O(N__66272),
            .I(N__66265));
    InMux I__15430 (
            .O(N__66271),
            .I(N__66262));
    InMux I__15429 (
            .O(N__66268),
            .I(N__66259));
    LocalMux I__15428 (
            .O(N__66265),
            .I(N__66256));
    LocalMux I__15427 (
            .O(N__66262),
            .I(N__66253));
    LocalMux I__15426 (
            .O(N__66259),
            .I(\c0.data_in_frame_15_4 ));
    Odrv12 I__15425 (
            .O(N__66256),
            .I(\c0.data_in_frame_15_4 ));
    Odrv4 I__15424 (
            .O(N__66253),
            .I(\c0.data_in_frame_15_4 ));
    InMux I__15423 (
            .O(N__66246),
            .I(N__66243));
    LocalMux I__15422 (
            .O(N__66243),
            .I(N__66239));
    InMux I__15421 (
            .O(N__66242),
            .I(N__66236));
    Span4Mux_v I__15420 (
            .O(N__66239),
            .I(N__66233));
    LocalMux I__15419 (
            .O(N__66236),
            .I(\c0.data_in_frame_18_2 ));
    Odrv4 I__15418 (
            .O(N__66233),
            .I(\c0.data_in_frame_18_2 ));
    InMux I__15417 (
            .O(N__66228),
            .I(N__66224));
    InMux I__15416 (
            .O(N__66227),
            .I(N__66221));
    LocalMux I__15415 (
            .O(N__66224),
            .I(N__66217));
    LocalMux I__15414 (
            .O(N__66221),
            .I(N__66214));
    CascadeMux I__15413 (
            .O(N__66220),
            .I(N__66211));
    Span4Mux_v I__15412 (
            .O(N__66217),
            .I(N__66208));
    Span4Mux_v I__15411 (
            .O(N__66214),
            .I(N__66205));
    InMux I__15410 (
            .O(N__66211),
            .I(N__66202));
    Span4Mux_h I__15409 (
            .O(N__66208),
            .I(N__66199));
    Span4Mux_v I__15408 (
            .O(N__66205),
            .I(N__66196));
    LocalMux I__15407 (
            .O(N__66202),
            .I(\c0.data_in_frame_18_4 ));
    Odrv4 I__15406 (
            .O(N__66199),
            .I(\c0.data_in_frame_18_4 ));
    Odrv4 I__15405 (
            .O(N__66196),
            .I(\c0.data_in_frame_18_4 ));
    InMux I__15404 (
            .O(N__66189),
            .I(N__66186));
    LocalMux I__15403 (
            .O(N__66186),
            .I(\c0.n12_adj_4455 ));
    CascadeMux I__15402 (
            .O(N__66183),
            .I(N__66180));
    InMux I__15401 (
            .O(N__66180),
            .I(N__66177));
    LocalMux I__15400 (
            .O(N__66177),
            .I(N__66174));
    Span12Mux_h I__15399 (
            .O(N__66174),
            .I(N__66170));
    InMux I__15398 (
            .O(N__66173),
            .I(N__66167));
    Odrv12 I__15397 (
            .O(N__66170),
            .I(\c0.n22463 ));
    LocalMux I__15396 (
            .O(N__66167),
            .I(\c0.n22463 ));
    InMux I__15395 (
            .O(N__66162),
            .I(N__66157));
    InMux I__15394 (
            .O(N__66161),
            .I(N__66154));
    InMux I__15393 (
            .O(N__66160),
            .I(N__66151));
    LocalMux I__15392 (
            .O(N__66157),
            .I(N__66146));
    LocalMux I__15391 (
            .O(N__66154),
            .I(N__66146));
    LocalMux I__15390 (
            .O(N__66151),
            .I(N__66143));
    Span4Mux_v I__15389 (
            .O(N__66146),
            .I(N__66138));
    Span4Mux_v I__15388 (
            .O(N__66143),
            .I(N__66138));
    Odrv4 I__15387 (
            .O(N__66138),
            .I(\c0.n24540 ));
    InMux I__15386 (
            .O(N__66135),
            .I(N__66130));
    InMux I__15385 (
            .O(N__66134),
            .I(N__66125));
    InMux I__15384 (
            .O(N__66133),
            .I(N__66125));
    LocalMux I__15383 (
            .O(N__66130),
            .I(N__66122));
    LocalMux I__15382 (
            .O(N__66125),
            .I(\c0.n23507 ));
    Odrv4 I__15381 (
            .O(N__66122),
            .I(\c0.n23507 ));
    CascadeMux I__15380 (
            .O(N__66117),
            .I(N__66113));
    InMux I__15379 (
            .O(N__66116),
            .I(N__66110));
    InMux I__15378 (
            .O(N__66113),
            .I(N__66107));
    LocalMux I__15377 (
            .O(N__66110),
            .I(N__66102));
    LocalMux I__15376 (
            .O(N__66107),
            .I(N__66102));
    Odrv4 I__15375 (
            .O(N__66102),
            .I(data_in_frame_21_0));
    InMux I__15374 (
            .O(N__66099),
            .I(N__66093));
    CascadeMux I__15373 (
            .O(N__66098),
            .I(N__66090));
    InMux I__15372 (
            .O(N__66097),
            .I(N__66087));
    InMux I__15371 (
            .O(N__66096),
            .I(N__66084));
    LocalMux I__15370 (
            .O(N__66093),
            .I(N__66081));
    InMux I__15369 (
            .O(N__66090),
            .I(N__66078));
    LocalMux I__15368 (
            .O(N__66087),
            .I(N__66073));
    LocalMux I__15367 (
            .O(N__66084),
            .I(N__66073));
    Span4Mux_h I__15366 (
            .O(N__66081),
            .I(N__66070));
    LocalMux I__15365 (
            .O(N__66078),
            .I(N__66063));
    Span4Mux_v I__15364 (
            .O(N__66073),
            .I(N__66063));
    Span4Mux_h I__15363 (
            .O(N__66070),
            .I(N__66063));
    Odrv4 I__15362 (
            .O(N__66063),
            .I(\c0.data_in_frame_17_0 ));
    InMux I__15361 (
            .O(N__66060),
            .I(N__66057));
    LocalMux I__15360 (
            .O(N__66057),
            .I(N__66054));
    Span4Mux_h I__15359 (
            .O(N__66054),
            .I(N__66049));
    InMux I__15358 (
            .O(N__66053),
            .I(N__66044));
    InMux I__15357 (
            .O(N__66052),
            .I(N__66044));
    Span4Mux_h I__15356 (
            .O(N__66049),
            .I(N__66041));
    LocalMux I__15355 (
            .O(N__66044),
            .I(N__66038));
    Odrv4 I__15354 (
            .O(N__66041),
            .I(\c0.n23313 ));
    Odrv4 I__15353 (
            .O(N__66038),
            .I(\c0.n23313 ));
    InMux I__15352 (
            .O(N__66033),
            .I(N__66027));
    InMux I__15351 (
            .O(N__66032),
            .I(N__66027));
    LocalMux I__15350 (
            .O(N__66027),
            .I(N__66024));
    Span4Mux_v I__15349 (
            .O(N__66024),
            .I(N__66021));
    Odrv4 I__15348 (
            .O(N__66021),
            .I(\c0.n26_adj_4578 ));
    InMux I__15347 (
            .O(N__66018),
            .I(N__66011));
    InMux I__15346 (
            .O(N__66017),
            .I(N__66011));
    CascadeMux I__15345 (
            .O(N__66016),
            .I(N__66007));
    LocalMux I__15344 (
            .O(N__66011),
            .I(N__66003));
    InMux I__15343 (
            .O(N__66010),
            .I(N__66000));
    InMux I__15342 (
            .O(N__66007),
            .I(N__65995));
    InMux I__15341 (
            .O(N__66006),
            .I(N__65995));
    Odrv4 I__15340 (
            .O(N__66003),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__15339 (
            .O(N__66000),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__15338 (
            .O(N__65995),
            .I(\c0.data_in_frame_13_5 ));
    InMux I__15337 (
            .O(N__65988),
            .I(N__65984));
    CascadeMux I__15336 (
            .O(N__65987),
            .I(N__65981));
    LocalMux I__15335 (
            .O(N__65984),
            .I(N__65977));
    InMux I__15334 (
            .O(N__65981),
            .I(N__65972));
    InMux I__15333 (
            .O(N__65980),
            .I(N__65972));
    Span4Mux_v I__15332 (
            .O(N__65977),
            .I(N__65969));
    LocalMux I__15331 (
            .O(N__65972),
            .I(\c0.data_in_frame_17_7 ));
    Odrv4 I__15330 (
            .O(N__65969),
            .I(\c0.data_in_frame_17_7 ));
    InMux I__15329 (
            .O(N__65964),
            .I(N__65961));
    LocalMux I__15328 (
            .O(N__65961),
            .I(N__65956));
    CascadeMux I__15327 (
            .O(N__65960),
            .I(N__65953));
    InMux I__15326 (
            .O(N__65959),
            .I(N__65950));
    Span4Mux_h I__15325 (
            .O(N__65956),
            .I(N__65947));
    InMux I__15324 (
            .O(N__65953),
            .I(N__65944));
    LocalMux I__15323 (
            .O(N__65950),
            .I(N__65941));
    Span4Mux_h I__15322 (
            .O(N__65947),
            .I(N__65938));
    LocalMux I__15321 (
            .O(N__65944),
            .I(\c0.data_in_frame_16_2 ));
    Odrv12 I__15320 (
            .O(N__65941),
            .I(\c0.data_in_frame_16_2 ));
    Odrv4 I__15319 (
            .O(N__65938),
            .I(\c0.data_in_frame_16_2 ));
    InMux I__15318 (
            .O(N__65931),
            .I(N__65928));
    LocalMux I__15317 (
            .O(N__65928),
            .I(N__65924));
    InMux I__15316 (
            .O(N__65927),
            .I(N__65921));
    Span4Mux_v I__15315 (
            .O(N__65924),
            .I(N__65918));
    LocalMux I__15314 (
            .O(N__65921),
            .I(N__65915));
    Span4Mux_h I__15313 (
            .O(N__65918),
            .I(N__65910));
    Span4Mux_v I__15312 (
            .O(N__65915),
            .I(N__65910));
    Span4Mux_v I__15311 (
            .O(N__65910),
            .I(N__65907));
    Odrv4 I__15310 (
            .O(N__65907),
            .I(\c0.n24527 ));
    InMux I__15309 (
            .O(N__65904),
            .I(N__65899));
    InMux I__15308 (
            .O(N__65903),
            .I(N__65896));
    CascadeMux I__15307 (
            .O(N__65902),
            .I(N__65893));
    LocalMux I__15306 (
            .O(N__65899),
            .I(N__65888));
    LocalMux I__15305 (
            .O(N__65896),
            .I(N__65888));
    InMux I__15304 (
            .O(N__65893),
            .I(N__65885));
    Span4Mux_h I__15303 (
            .O(N__65888),
            .I(N__65881));
    LocalMux I__15302 (
            .O(N__65885),
            .I(N__65878));
    InMux I__15301 (
            .O(N__65884),
            .I(N__65875));
    Span4Mux_h I__15300 (
            .O(N__65881),
            .I(N__65872));
    Span4Mux_h I__15299 (
            .O(N__65878),
            .I(N__65869));
    LocalMux I__15298 (
            .O(N__65875),
            .I(data_in_frame_21_3));
    Odrv4 I__15297 (
            .O(N__65872),
            .I(data_in_frame_21_3));
    Odrv4 I__15296 (
            .O(N__65869),
            .I(data_in_frame_21_3));
    InMux I__15295 (
            .O(N__65862),
            .I(N__65858));
    InMux I__15294 (
            .O(N__65861),
            .I(N__65855));
    LocalMux I__15293 (
            .O(N__65858),
            .I(N__65850));
    LocalMux I__15292 (
            .O(N__65855),
            .I(N__65847));
    InMux I__15291 (
            .O(N__65854),
            .I(N__65841));
    InMux I__15290 (
            .O(N__65853),
            .I(N__65841));
    Span4Mux_v I__15289 (
            .O(N__65850),
            .I(N__65836));
    Span4Mux_h I__15288 (
            .O(N__65847),
            .I(N__65836));
    InMux I__15287 (
            .O(N__65846),
            .I(N__65832));
    LocalMux I__15286 (
            .O(N__65841),
            .I(N__65829));
    Span4Mux_h I__15285 (
            .O(N__65836),
            .I(N__65826));
    InMux I__15284 (
            .O(N__65835),
            .I(N__65823));
    LocalMux I__15283 (
            .O(N__65832),
            .I(\c0.n21344 ));
    Odrv4 I__15282 (
            .O(N__65829),
            .I(\c0.n21344 ));
    Odrv4 I__15281 (
            .O(N__65826),
            .I(\c0.n21344 ));
    LocalMux I__15280 (
            .O(N__65823),
            .I(\c0.n21344 ));
    InMux I__15279 (
            .O(N__65814),
            .I(N__65811));
    LocalMux I__15278 (
            .O(N__65811),
            .I(N__65808));
    Odrv4 I__15277 (
            .O(N__65808),
            .I(\c0.n42_adj_4589 ));
    InMux I__15276 (
            .O(N__65805),
            .I(N__65802));
    LocalMux I__15275 (
            .O(N__65802),
            .I(N__65799));
    Span4Mux_v I__15274 (
            .O(N__65799),
            .I(N__65795));
    InMux I__15273 (
            .O(N__65798),
            .I(N__65792));
    Odrv4 I__15272 (
            .O(N__65795),
            .I(\c0.n22_adj_4243 ));
    LocalMux I__15271 (
            .O(N__65792),
            .I(\c0.n22_adj_4243 ));
    InMux I__15270 (
            .O(N__65787),
            .I(N__65783));
    InMux I__15269 (
            .O(N__65786),
            .I(N__65780));
    LocalMux I__15268 (
            .O(N__65783),
            .I(N__65776));
    LocalMux I__15267 (
            .O(N__65780),
            .I(N__65773));
    CascadeMux I__15266 (
            .O(N__65779),
            .I(N__65769));
    Span4Mux_v I__15265 (
            .O(N__65776),
            .I(N__65766));
    Span4Mux_h I__15264 (
            .O(N__65773),
            .I(N__65763));
    InMux I__15263 (
            .O(N__65772),
            .I(N__65760));
    InMux I__15262 (
            .O(N__65769),
            .I(N__65757));
    Odrv4 I__15261 (
            .O(N__65766),
            .I(\c0.n13738 ));
    Odrv4 I__15260 (
            .O(N__65763),
            .I(\c0.n13738 ));
    LocalMux I__15259 (
            .O(N__65760),
            .I(\c0.n13738 ));
    LocalMux I__15258 (
            .O(N__65757),
            .I(\c0.n13738 ));
    CascadeMux I__15257 (
            .O(N__65748),
            .I(N__65744));
    CascadeMux I__15256 (
            .O(N__65747),
            .I(N__65741));
    InMux I__15255 (
            .O(N__65744),
            .I(N__65738));
    InMux I__15254 (
            .O(N__65741),
            .I(N__65735));
    LocalMux I__15253 (
            .O(N__65738),
            .I(N__65732));
    LocalMux I__15252 (
            .O(N__65735),
            .I(N__65729));
    Span4Mux_h I__15251 (
            .O(N__65732),
            .I(N__65726));
    Odrv12 I__15250 (
            .O(N__65729),
            .I(\c0.n10_adj_4230 ));
    Odrv4 I__15249 (
            .O(N__65726),
            .I(\c0.n10_adj_4230 ));
    InMux I__15248 (
            .O(N__65721),
            .I(N__65718));
    LocalMux I__15247 (
            .O(N__65718),
            .I(N__65714));
    InMux I__15246 (
            .O(N__65717),
            .I(N__65711));
    Odrv4 I__15245 (
            .O(N__65714),
            .I(\c0.n5_adj_4310 ));
    LocalMux I__15244 (
            .O(N__65711),
            .I(\c0.n5_adj_4310 ));
    InMux I__15243 (
            .O(N__65706),
            .I(N__65698));
    InMux I__15242 (
            .O(N__65705),
            .I(N__65698));
    InMux I__15241 (
            .O(N__65704),
            .I(N__65691));
    InMux I__15240 (
            .O(N__65703),
            .I(N__65691));
    LocalMux I__15239 (
            .O(N__65698),
            .I(N__65688));
    CascadeMux I__15238 (
            .O(N__65697),
            .I(N__65685));
    CascadeMux I__15237 (
            .O(N__65696),
            .I(N__65682));
    LocalMux I__15236 (
            .O(N__65691),
            .I(N__65679));
    Span4Mux_v I__15235 (
            .O(N__65688),
            .I(N__65675));
    InMux I__15234 (
            .O(N__65685),
            .I(N__65670));
    InMux I__15233 (
            .O(N__65682),
            .I(N__65670));
    Span4Mux_v I__15232 (
            .O(N__65679),
            .I(N__65667));
    InMux I__15231 (
            .O(N__65678),
            .I(N__65664));
    Odrv4 I__15230 (
            .O(N__65675),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__15229 (
            .O(N__65670),
            .I(\c0.data_in_frame_4_5 ));
    Odrv4 I__15228 (
            .O(N__65667),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__15227 (
            .O(N__65664),
            .I(\c0.data_in_frame_4_5 ));
    CascadeMux I__15226 (
            .O(N__65655),
            .I(N__65651));
    InMux I__15225 (
            .O(N__65654),
            .I(N__65646));
    InMux I__15224 (
            .O(N__65651),
            .I(N__65646));
    LocalMux I__15223 (
            .O(N__65646),
            .I(N__65643));
    Odrv12 I__15222 (
            .O(N__65643),
            .I(\c0.n23283 ));
    InMux I__15221 (
            .O(N__65640),
            .I(N__65634));
    InMux I__15220 (
            .O(N__65639),
            .I(N__65627));
    InMux I__15219 (
            .O(N__65638),
            .I(N__65624));
    InMux I__15218 (
            .O(N__65637),
            .I(N__65621));
    LocalMux I__15217 (
            .O(N__65634),
            .I(N__65618));
    InMux I__15216 (
            .O(N__65633),
            .I(N__65613));
    InMux I__15215 (
            .O(N__65632),
            .I(N__65613));
    InMux I__15214 (
            .O(N__65631),
            .I(N__65608));
    InMux I__15213 (
            .O(N__65630),
            .I(N__65608));
    LocalMux I__15212 (
            .O(N__65627),
            .I(\c0.data_in_frame_8_7 ));
    LocalMux I__15211 (
            .O(N__65624),
            .I(\c0.data_in_frame_8_7 ));
    LocalMux I__15210 (
            .O(N__65621),
            .I(\c0.data_in_frame_8_7 ));
    Odrv4 I__15209 (
            .O(N__65618),
            .I(\c0.data_in_frame_8_7 ));
    LocalMux I__15208 (
            .O(N__65613),
            .I(\c0.data_in_frame_8_7 ));
    LocalMux I__15207 (
            .O(N__65608),
            .I(\c0.data_in_frame_8_7 ));
    InMux I__15206 (
            .O(N__65595),
            .I(N__65592));
    LocalMux I__15205 (
            .O(N__65592),
            .I(N__65588));
    InMux I__15204 (
            .O(N__65591),
            .I(N__65585));
    Odrv12 I__15203 (
            .O(N__65588),
            .I(\c0.n20_adj_4260 ));
    LocalMux I__15202 (
            .O(N__65585),
            .I(\c0.n20_adj_4260 ));
    CascadeMux I__15201 (
            .O(N__65580),
            .I(N__65577));
    InMux I__15200 (
            .O(N__65577),
            .I(N__65573));
    InMux I__15199 (
            .O(N__65576),
            .I(N__65570));
    LocalMux I__15198 (
            .O(N__65573),
            .I(N__65567));
    LocalMux I__15197 (
            .O(N__65570),
            .I(N__65564));
    Span4Mux_h I__15196 (
            .O(N__65567),
            .I(N__65561));
    Span4Mux_v I__15195 (
            .O(N__65564),
            .I(N__65558));
    Odrv4 I__15194 (
            .O(N__65561),
            .I(\c0.n22803 ));
    Odrv4 I__15193 (
            .O(N__65558),
            .I(\c0.n22803 ));
    InMux I__15192 (
            .O(N__65553),
            .I(N__65550));
    LocalMux I__15191 (
            .O(N__65550),
            .I(N__65546));
    InMux I__15190 (
            .O(N__65549),
            .I(N__65543));
    Odrv4 I__15189 (
            .O(N__65546),
            .I(\c0.n4_adj_4261 ));
    LocalMux I__15188 (
            .O(N__65543),
            .I(\c0.n4_adj_4261 ));
    InMux I__15187 (
            .O(N__65538),
            .I(N__65535));
    LocalMux I__15186 (
            .O(N__65535),
            .I(N__65532));
    Span12Mux_h I__15185 (
            .O(N__65532),
            .I(N__65529));
    Odrv12 I__15184 (
            .O(N__65529),
            .I(\c0.n31_adj_4743 ));
    InMux I__15183 (
            .O(N__65526),
            .I(N__65522));
    InMux I__15182 (
            .O(N__65525),
            .I(N__65519));
    LocalMux I__15181 (
            .O(N__65522),
            .I(N__65516));
    LocalMux I__15180 (
            .O(N__65519),
            .I(\c0.n5813 ));
    Odrv4 I__15179 (
            .O(N__65516),
            .I(\c0.n5813 ));
    CascadeMux I__15178 (
            .O(N__65511),
            .I(N__65507));
    CascadeMux I__15177 (
            .O(N__65510),
            .I(N__65504));
    InMux I__15176 (
            .O(N__65507),
            .I(N__65501));
    InMux I__15175 (
            .O(N__65504),
            .I(N__65498));
    LocalMux I__15174 (
            .O(N__65501),
            .I(\c0.n22602 ));
    LocalMux I__15173 (
            .O(N__65498),
            .I(\c0.n22602 ));
    InMux I__15172 (
            .O(N__65493),
            .I(N__65489));
    InMux I__15171 (
            .O(N__65492),
            .I(N__65486));
    LocalMux I__15170 (
            .O(N__65489),
            .I(N__65481));
    LocalMux I__15169 (
            .O(N__65486),
            .I(N__65481));
    Span4Mux_v I__15168 (
            .O(N__65481),
            .I(N__65478));
    Odrv4 I__15167 (
            .O(N__65478),
            .I(\c0.n11 ));
    InMux I__15166 (
            .O(N__65475),
            .I(N__65472));
    LocalMux I__15165 (
            .O(N__65472),
            .I(N__65469));
    Odrv12 I__15164 (
            .O(N__65469),
            .I(\c0.n17_adj_4219 ));
    CascadeMux I__15163 (
            .O(N__65466),
            .I(\c0.n16_adj_4218_cascade_ ));
    CascadeMux I__15162 (
            .O(N__65463),
            .I(\c0.n13767_cascade_ ));
    InMux I__15161 (
            .O(N__65460),
            .I(N__65457));
    LocalMux I__15160 (
            .O(N__65457),
            .I(N__65454));
    Span4Mux_v I__15159 (
            .O(N__65454),
            .I(N__65450));
    InMux I__15158 (
            .O(N__65453),
            .I(N__65447));
    Span4Mux_h I__15157 (
            .O(N__65450),
            .I(N__65444));
    LocalMux I__15156 (
            .O(N__65447),
            .I(N__65441));
    Odrv4 I__15155 (
            .O(N__65444),
            .I(\c0.n5965 ));
    Odrv4 I__15154 (
            .O(N__65441),
            .I(\c0.n5965 ));
    InMux I__15153 (
            .O(N__65436),
            .I(N__65430));
    InMux I__15152 (
            .O(N__65435),
            .I(N__65430));
    LocalMux I__15151 (
            .O(N__65430),
            .I(\c0.n6_adj_4454 ));
    InMux I__15150 (
            .O(N__65427),
            .I(N__65423));
    CascadeMux I__15149 (
            .O(N__65426),
            .I(N__65420));
    LocalMux I__15148 (
            .O(N__65423),
            .I(N__65416));
    InMux I__15147 (
            .O(N__65420),
            .I(N__65413));
    InMux I__15146 (
            .O(N__65419),
            .I(N__65410));
    Span4Mux_v I__15145 (
            .O(N__65416),
            .I(N__65407));
    LocalMux I__15144 (
            .O(N__65413),
            .I(N__65398));
    LocalMux I__15143 (
            .O(N__65410),
            .I(N__65398));
    Sp12to4 I__15142 (
            .O(N__65407),
            .I(N__65398));
    InMux I__15141 (
            .O(N__65406),
            .I(N__65395));
    InMux I__15140 (
            .O(N__65405),
            .I(N__65392));
    Odrv12 I__15139 (
            .O(N__65398),
            .I(\c0.data_in_frame_15_3 ));
    LocalMux I__15138 (
            .O(N__65395),
            .I(\c0.data_in_frame_15_3 ));
    LocalMux I__15137 (
            .O(N__65392),
            .I(\c0.data_in_frame_15_3 ));
    InMux I__15136 (
            .O(N__65385),
            .I(N__65382));
    LocalMux I__15135 (
            .O(N__65382),
            .I(N__65379));
    Span4Mux_v I__15134 (
            .O(N__65379),
            .I(N__65376));
    Span4Mux_v I__15133 (
            .O(N__65376),
            .I(N__65373));
    Odrv4 I__15132 (
            .O(N__65373),
            .I(\c0.n23_adj_4665 ));
    InMux I__15131 (
            .O(N__65370),
            .I(N__65365));
    CascadeMux I__15130 (
            .O(N__65369),
            .I(N__65362));
    CascadeMux I__15129 (
            .O(N__65368),
            .I(N__65359));
    LocalMux I__15128 (
            .O(N__65365),
            .I(N__65356));
    InMux I__15127 (
            .O(N__65362),
            .I(N__65353));
    InMux I__15126 (
            .O(N__65359),
            .I(N__65350));
    Span4Mux_h I__15125 (
            .O(N__65356),
            .I(N__65347));
    LocalMux I__15124 (
            .O(N__65353),
            .I(N__65344));
    LocalMux I__15123 (
            .O(N__65350),
            .I(\c0.data_in_frame_15_2 ));
    Odrv4 I__15122 (
            .O(N__65347),
            .I(\c0.data_in_frame_15_2 ));
    Odrv4 I__15121 (
            .O(N__65344),
            .I(\c0.data_in_frame_15_2 ));
    CascadeMux I__15120 (
            .O(N__65337),
            .I(N__65332));
    InMux I__15119 (
            .O(N__65336),
            .I(N__65328));
    InMux I__15118 (
            .O(N__65335),
            .I(N__65324));
    InMux I__15117 (
            .O(N__65332),
            .I(N__65319));
    InMux I__15116 (
            .O(N__65331),
            .I(N__65319));
    LocalMux I__15115 (
            .O(N__65328),
            .I(N__65316));
    InMux I__15114 (
            .O(N__65327),
            .I(N__65313));
    LocalMux I__15113 (
            .O(N__65324),
            .I(\c0.data_in_frame_8_5 ));
    LocalMux I__15112 (
            .O(N__65319),
            .I(\c0.data_in_frame_8_5 ));
    Odrv4 I__15111 (
            .O(N__65316),
            .I(\c0.data_in_frame_8_5 ));
    LocalMux I__15110 (
            .O(N__65313),
            .I(\c0.data_in_frame_8_5 ));
    CascadeMux I__15109 (
            .O(N__65304),
            .I(N__65301));
    InMux I__15108 (
            .O(N__65301),
            .I(N__65298));
    LocalMux I__15107 (
            .O(N__65298),
            .I(N__65292));
    InMux I__15106 (
            .O(N__65297),
            .I(N__65287));
    InMux I__15105 (
            .O(N__65296),
            .I(N__65287));
    CascadeMux I__15104 (
            .O(N__65295),
            .I(N__65283));
    Span4Mux_v I__15103 (
            .O(N__65292),
            .I(N__65278));
    LocalMux I__15102 (
            .O(N__65287),
            .I(N__65278));
    CascadeMux I__15101 (
            .O(N__65286),
            .I(N__65275));
    InMux I__15100 (
            .O(N__65283),
            .I(N__65272));
    Span4Mux_h I__15099 (
            .O(N__65278),
            .I(N__65269));
    InMux I__15098 (
            .O(N__65275),
            .I(N__65266));
    LocalMux I__15097 (
            .O(N__65272),
            .I(N__65263));
    Span4Mux_h I__15096 (
            .O(N__65269),
            .I(N__65260));
    LocalMux I__15095 (
            .O(N__65266),
            .I(\c0.data_in_frame_11_1 ));
    Odrv12 I__15094 (
            .O(N__65263),
            .I(\c0.data_in_frame_11_1 ));
    Odrv4 I__15093 (
            .O(N__65260),
            .I(\c0.data_in_frame_11_1 ));
    InMux I__15092 (
            .O(N__65253),
            .I(N__65250));
    LocalMux I__15091 (
            .O(N__65250),
            .I(\c0.n22176 ));
    CascadeMux I__15090 (
            .O(N__65247),
            .I(\c0.n28_adj_4637_cascade_ ));
    InMux I__15089 (
            .O(N__65244),
            .I(N__65241));
    LocalMux I__15088 (
            .O(N__65241),
            .I(\c0.n24_adj_4636 ));
    InMux I__15087 (
            .O(N__65238),
            .I(N__65235));
    LocalMux I__15086 (
            .O(N__65235),
            .I(\c0.n7_adj_4634 ));
    InMux I__15085 (
            .O(N__65232),
            .I(N__65229));
    LocalMux I__15084 (
            .O(N__65229),
            .I(\c0.n16_adj_4635 ));
    InMux I__15083 (
            .O(N__65226),
            .I(N__65223));
    LocalMux I__15082 (
            .O(N__65223),
            .I(N__65217));
    InMux I__15081 (
            .O(N__65222),
            .I(N__65214));
    InMux I__15080 (
            .O(N__65221),
            .I(N__65209));
    InMux I__15079 (
            .O(N__65220),
            .I(N__65209));
    Odrv4 I__15078 (
            .O(N__65217),
            .I(\c0.n23406 ));
    LocalMux I__15077 (
            .O(N__65214),
            .I(\c0.n23406 ));
    LocalMux I__15076 (
            .O(N__65209),
            .I(\c0.n23406 ));
    InMux I__15075 (
            .O(N__65202),
            .I(N__65197));
    InMux I__15074 (
            .O(N__65201),
            .I(N__65194));
    InMux I__15073 (
            .O(N__65200),
            .I(N__65190));
    LocalMux I__15072 (
            .O(N__65197),
            .I(N__65185));
    LocalMux I__15071 (
            .O(N__65194),
            .I(N__65185));
    InMux I__15070 (
            .O(N__65193),
            .I(N__65181));
    LocalMux I__15069 (
            .O(N__65190),
            .I(N__65178));
    Span4Mux_h I__15068 (
            .O(N__65185),
            .I(N__65175));
    InMux I__15067 (
            .O(N__65184),
            .I(N__65172));
    LocalMux I__15066 (
            .O(N__65181),
            .I(data_in_frame_6_4));
    Odrv12 I__15065 (
            .O(N__65178),
            .I(data_in_frame_6_4));
    Odrv4 I__15064 (
            .O(N__65175),
            .I(data_in_frame_6_4));
    LocalMux I__15063 (
            .O(N__65172),
            .I(data_in_frame_6_4));
    CascadeMux I__15062 (
            .O(N__65163),
            .I(\c0.n14_adj_4609_cascade_ ));
    InMux I__15061 (
            .O(N__65160),
            .I(N__65157));
    LocalMux I__15060 (
            .O(N__65157),
            .I(\c0.n10_adj_4617 ));
    InMux I__15059 (
            .O(N__65154),
            .I(N__65151));
    LocalMux I__15058 (
            .O(N__65151),
            .I(N__65147));
    InMux I__15057 (
            .O(N__65150),
            .I(N__65144));
    Span4Mux_v I__15056 (
            .O(N__65147),
            .I(N__65140));
    LocalMux I__15055 (
            .O(N__65144),
            .I(N__65137));
    InMux I__15054 (
            .O(N__65143),
            .I(N__65134));
    Odrv4 I__15053 (
            .O(N__65140),
            .I(\c0.n17 ));
    Odrv12 I__15052 (
            .O(N__65137),
            .I(\c0.n17 ));
    LocalMux I__15051 (
            .O(N__65134),
            .I(\c0.n17 ));
    InMux I__15050 (
            .O(N__65127),
            .I(N__65121));
    InMux I__15049 (
            .O(N__65126),
            .I(N__65121));
    LocalMux I__15048 (
            .O(N__65121),
            .I(N__65118));
    Odrv12 I__15047 (
            .O(N__65118),
            .I(\c0.n8_adj_4216 ));
    CascadeMux I__15046 (
            .O(N__65115),
            .I(\c0.n12_cascade_ ));
    InMux I__15045 (
            .O(N__65112),
            .I(N__65105));
    InMux I__15044 (
            .O(N__65111),
            .I(N__65102));
    InMux I__15043 (
            .O(N__65110),
            .I(N__65097));
    InMux I__15042 (
            .O(N__65109),
            .I(N__65097));
    InMux I__15041 (
            .O(N__65108),
            .I(N__65093));
    LocalMux I__15040 (
            .O(N__65105),
            .I(N__65088));
    LocalMux I__15039 (
            .O(N__65102),
            .I(N__65088));
    LocalMux I__15038 (
            .O(N__65097),
            .I(N__65085));
    InMux I__15037 (
            .O(N__65096),
            .I(N__65082));
    LocalMux I__15036 (
            .O(N__65093),
            .I(N__65079));
    Span4Mux_v I__15035 (
            .O(N__65088),
            .I(N__65074));
    Span4Mux_h I__15034 (
            .O(N__65085),
            .I(N__65074));
    LocalMux I__15033 (
            .O(N__65082),
            .I(N__65070));
    Span12Mux_h I__15032 (
            .O(N__65079),
            .I(N__65065));
    Span4Mux_h I__15031 (
            .O(N__65074),
            .I(N__65062));
    InMux I__15030 (
            .O(N__65073),
            .I(N__65059));
    Span4Mux_v I__15029 (
            .O(N__65070),
            .I(N__65056));
    InMux I__15028 (
            .O(N__65069),
            .I(N__65051));
    InMux I__15027 (
            .O(N__65068),
            .I(N__65051));
    Odrv12 I__15026 (
            .O(N__65065),
            .I(\c0.data_in_frame_4_2 ));
    Odrv4 I__15025 (
            .O(N__65062),
            .I(\c0.data_in_frame_4_2 ));
    LocalMux I__15024 (
            .O(N__65059),
            .I(\c0.data_in_frame_4_2 ));
    Odrv4 I__15023 (
            .O(N__65056),
            .I(\c0.data_in_frame_4_2 ));
    LocalMux I__15022 (
            .O(N__65051),
            .I(\c0.data_in_frame_4_2 ));
    CascadeMux I__15021 (
            .O(N__65040),
            .I(N__65036));
    CascadeMux I__15020 (
            .O(N__65039),
            .I(N__65032));
    InMux I__15019 (
            .O(N__65036),
            .I(N__65029));
    CascadeMux I__15018 (
            .O(N__65035),
            .I(N__65026));
    InMux I__15017 (
            .O(N__65032),
            .I(N__65023));
    LocalMux I__15016 (
            .O(N__65029),
            .I(N__65020));
    InMux I__15015 (
            .O(N__65026),
            .I(N__65017));
    LocalMux I__15014 (
            .O(N__65023),
            .I(\c0.data_in_frame_12_2 ));
    Odrv4 I__15013 (
            .O(N__65020),
            .I(\c0.data_in_frame_12_2 ));
    LocalMux I__15012 (
            .O(N__65017),
            .I(\c0.data_in_frame_12_2 ));
    InMux I__15011 (
            .O(N__65010),
            .I(N__65006));
    InMux I__15010 (
            .O(N__65009),
            .I(N__65003));
    LocalMux I__15009 (
            .O(N__65006),
            .I(N__65000));
    LocalMux I__15008 (
            .O(N__65003),
            .I(N__64997));
    Span4Mux_h I__15007 (
            .O(N__65000),
            .I(N__64994));
    Odrv4 I__15006 (
            .O(N__64997),
            .I(\c0.n13809 ));
    Odrv4 I__15005 (
            .O(N__64994),
            .I(\c0.n13809 ));
    CascadeMux I__15004 (
            .O(N__64989),
            .I(N__64983));
    InMux I__15003 (
            .O(N__64988),
            .I(N__64980));
    CascadeMux I__15002 (
            .O(N__64987),
            .I(N__64977));
    InMux I__15001 (
            .O(N__64986),
            .I(N__64974));
    InMux I__15000 (
            .O(N__64983),
            .I(N__64971));
    LocalMux I__14999 (
            .O(N__64980),
            .I(N__64968));
    InMux I__14998 (
            .O(N__64977),
            .I(N__64962));
    LocalMux I__14997 (
            .O(N__64974),
            .I(N__64959));
    LocalMux I__14996 (
            .O(N__64971),
            .I(N__64956));
    Span4Mux_v I__14995 (
            .O(N__64968),
            .I(N__64953));
    InMux I__14994 (
            .O(N__64967),
            .I(N__64950));
    CascadeMux I__14993 (
            .O(N__64966),
            .I(N__64947));
    InMux I__14992 (
            .O(N__64965),
            .I(N__64944));
    LocalMux I__14991 (
            .O(N__64962),
            .I(N__64939));
    Span4Mux_v I__14990 (
            .O(N__64959),
            .I(N__64939));
    Span4Mux_v I__14989 (
            .O(N__64956),
            .I(N__64936));
    Span4Mux_h I__14988 (
            .O(N__64953),
            .I(N__64931));
    LocalMux I__14987 (
            .O(N__64950),
            .I(N__64931));
    InMux I__14986 (
            .O(N__64947),
            .I(N__64928));
    LocalMux I__14985 (
            .O(N__64944),
            .I(N__64923));
    Span4Mux_h I__14984 (
            .O(N__64939),
            .I(N__64923));
    Odrv4 I__14983 (
            .O(N__64936),
            .I(\c0.data_in_frame_11_5 ));
    Odrv4 I__14982 (
            .O(N__64931),
            .I(\c0.data_in_frame_11_5 ));
    LocalMux I__14981 (
            .O(N__64928),
            .I(\c0.data_in_frame_11_5 ));
    Odrv4 I__14980 (
            .O(N__64923),
            .I(\c0.data_in_frame_11_5 ));
    InMux I__14979 (
            .O(N__64914),
            .I(N__64911));
    LocalMux I__14978 (
            .O(N__64911),
            .I(N__64908));
    Span4Mux_v I__14977 (
            .O(N__64908),
            .I(N__64905));
    Odrv4 I__14976 (
            .O(N__64905),
            .I(\c0.n22751 ));
    CascadeMux I__14975 (
            .O(N__64902),
            .I(N__64898));
    CascadeMux I__14974 (
            .O(N__64901),
            .I(N__64894));
    InMux I__14973 (
            .O(N__64898),
            .I(N__64891));
    InMux I__14972 (
            .O(N__64897),
            .I(N__64888));
    InMux I__14971 (
            .O(N__64894),
            .I(N__64885));
    LocalMux I__14970 (
            .O(N__64891),
            .I(N__64880));
    LocalMux I__14969 (
            .O(N__64888),
            .I(N__64877));
    LocalMux I__14968 (
            .O(N__64885),
            .I(N__64874));
    InMux I__14967 (
            .O(N__64884),
            .I(N__64868));
    InMux I__14966 (
            .O(N__64883),
            .I(N__64868));
    Span4Mux_v I__14965 (
            .O(N__64880),
            .I(N__64863));
    Span4Mux_h I__14964 (
            .O(N__64877),
            .I(N__64863));
    Span4Mux_h I__14963 (
            .O(N__64874),
            .I(N__64860));
    InMux I__14962 (
            .O(N__64873),
            .I(N__64857));
    LocalMux I__14961 (
            .O(N__64868),
            .I(N__64854));
    Span4Mux_h I__14960 (
            .O(N__64863),
            .I(N__64851));
    Span4Mux_h I__14959 (
            .O(N__64860),
            .I(N__64848));
    LocalMux I__14958 (
            .O(N__64857),
            .I(data_in_frame_6_7));
    Odrv12 I__14957 (
            .O(N__64854),
            .I(data_in_frame_6_7));
    Odrv4 I__14956 (
            .O(N__64851),
            .I(data_in_frame_6_7));
    Odrv4 I__14955 (
            .O(N__64848),
            .I(data_in_frame_6_7));
    InMux I__14954 (
            .O(N__64839),
            .I(N__64835));
    CascadeMux I__14953 (
            .O(N__64838),
            .I(N__64831));
    LocalMux I__14952 (
            .O(N__64835),
            .I(N__64828));
    InMux I__14951 (
            .O(N__64834),
            .I(N__64824));
    InMux I__14950 (
            .O(N__64831),
            .I(N__64821));
    Span4Mux_h I__14949 (
            .O(N__64828),
            .I(N__64814));
    InMux I__14948 (
            .O(N__64827),
            .I(N__64811));
    LocalMux I__14947 (
            .O(N__64824),
            .I(N__64808));
    LocalMux I__14946 (
            .O(N__64821),
            .I(N__64805));
    InMux I__14945 (
            .O(N__64820),
            .I(N__64796));
    InMux I__14944 (
            .O(N__64819),
            .I(N__64796));
    InMux I__14943 (
            .O(N__64818),
            .I(N__64796));
    InMux I__14942 (
            .O(N__64817),
            .I(N__64796));
    Span4Mux_h I__14941 (
            .O(N__64814),
            .I(N__64793));
    LocalMux I__14940 (
            .O(N__64811),
            .I(N__64788));
    Span12Mux_v I__14939 (
            .O(N__64808),
            .I(N__64788));
    Odrv12 I__14938 (
            .O(N__64805),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__14937 (
            .O(N__64796),
            .I(\c0.data_in_frame_4_7 ));
    Odrv4 I__14936 (
            .O(N__64793),
            .I(\c0.data_in_frame_4_7 ));
    Odrv12 I__14935 (
            .O(N__64788),
            .I(\c0.data_in_frame_4_7 ));
    InMux I__14934 (
            .O(N__64779),
            .I(N__64774));
    InMux I__14933 (
            .O(N__64778),
            .I(N__64769));
    InMux I__14932 (
            .O(N__64777),
            .I(N__64765));
    LocalMux I__14931 (
            .O(N__64774),
            .I(N__64761));
    InMux I__14930 (
            .O(N__64773),
            .I(N__64756));
    InMux I__14929 (
            .O(N__64772),
            .I(N__64756));
    LocalMux I__14928 (
            .O(N__64769),
            .I(N__64752));
    InMux I__14927 (
            .O(N__64768),
            .I(N__64749));
    LocalMux I__14926 (
            .O(N__64765),
            .I(N__64746));
    InMux I__14925 (
            .O(N__64764),
            .I(N__64743));
    Span4Mux_v I__14924 (
            .O(N__64761),
            .I(N__64738));
    LocalMux I__14923 (
            .O(N__64756),
            .I(N__64738));
    CascadeMux I__14922 (
            .O(N__64755),
            .I(N__64734));
    Span4Mux_h I__14921 (
            .O(N__64752),
            .I(N__64728));
    LocalMux I__14920 (
            .O(N__64749),
            .I(N__64728));
    Span4Mux_h I__14919 (
            .O(N__64746),
            .I(N__64725));
    LocalMux I__14918 (
            .O(N__64743),
            .I(N__64719));
    Span4Mux_h I__14917 (
            .O(N__64738),
            .I(N__64719));
    InMux I__14916 (
            .O(N__64737),
            .I(N__64716));
    InMux I__14915 (
            .O(N__64734),
            .I(N__64713));
    InMux I__14914 (
            .O(N__64733),
            .I(N__64710));
    Span4Mux_h I__14913 (
            .O(N__64728),
            .I(N__64705));
    Span4Mux_h I__14912 (
            .O(N__64725),
            .I(N__64705));
    InMux I__14911 (
            .O(N__64724),
            .I(N__64702));
    Sp12to4 I__14910 (
            .O(N__64719),
            .I(N__64697));
    LocalMux I__14909 (
            .O(N__64716),
            .I(N__64697));
    LocalMux I__14908 (
            .O(N__64713),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__14907 (
            .O(N__64710),
            .I(\c0.data_in_frame_2_7 ));
    Odrv4 I__14906 (
            .O(N__64705),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__14905 (
            .O(N__64702),
            .I(\c0.data_in_frame_2_7 ));
    Odrv12 I__14904 (
            .O(N__64697),
            .I(\c0.data_in_frame_2_7 ));
    CascadeMux I__14903 (
            .O(N__64686),
            .I(N__64683));
    InMux I__14902 (
            .O(N__64683),
            .I(N__64680));
    LocalMux I__14901 (
            .O(N__64680),
            .I(\c0.n49 ));
    InMux I__14900 (
            .O(N__64677),
            .I(N__64674));
    LocalMux I__14899 (
            .O(N__64674),
            .I(N__64670));
    InMux I__14898 (
            .O(N__64673),
            .I(N__64667));
    Odrv12 I__14897 (
            .O(N__64670),
            .I(\c0.n23528 ));
    LocalMux I__14896 (
            .O(N__64667),
            .I(\c0.n23528 ));
    InMux I__14895 (
            .O(N__64662),
            .I(N__64659));
    LocalMux I__14894 (
            .O(N__64659),
            .I(N__64656));
    Span4Mux_v I__14893 (
            .O(N__64656),
            .I(N__64652));
    InMux I__14892 (
            .O(N__64655),
            .I(N__64649));
    Span4Mux_h I__14891 (
            .O(N__64652),
            .I(N__64644));
    LocalMux I__14890 (
            .O(N__64649),
            .I(N__64644));
    Span4Mux_v I__14889 (
            .O(N__64644),
            .I(N__64641));
    Odrv4 I__14888 (
            .O(N__64641),
            .I(\c0.n7_adj_4229 ));
    InMux I__14887 (
            .O(N__64638),
            .I(N__64635));
    LocalMux I__14886 (
            .O(N__64635),
            .I(N__64630));
    InMux I__14885 (
            .O(N__64634),
            .I(N__64625));
    InMux I__14884 (
            .O(N__64633),
            .I(N__64625));
    Span12Mux_v I__14883 (
            .O(N__64630),
            .I(N__64622));
    LocalMux I__14882 (
            .O(N__64625),
            .I(N__64619));
    Odrv12 I__14881 (
            .O(N__64622),
            .I(\c0.data_out_frame_0__7__N_2743 ));
    Odrv4 I__14880 (
            .O(N__64619),
            .I(\c0.data_out_frame_0__7__N_2743 ));
    InMux I__14879 (
            .O(N__64614),
            .I(N__64610));
    InMux I__14878 (
            .O(N__64613),
            .I(N__64607));
    LocalMux I__14877 (
            .O(N__64610),
            .I(N__64602));
    LocalMux I__14876 (
            .O(N__64607),
            .I(N__64599));
    InMux I__14875 (
            .O(N__64606),
            .I(N__64596));
    InMux I__14874 (
            .O(N__64605),
            .I(N__64593));
    Span4Mux_v I__14873 (
            .O(N__64602),
            .I(N__64590));
    Span4Mux_v I__14872 (
            .O(N__64599),
            .I(N__64585));
    LocalMux I__14871 (
            .O(N__64596),
            .I(N__64585));
    LocalMux I__14870 (
            .O(N__64593),
            .I(N__64582));
    Span4Mux_h I__14869 (
            .O(N__64590),
            .I(N__64578));
    Span4Mux_v I__14868 (
            .O(N__64585),
            .I(N__64573));
    Span4Mux_v I__14867 (
            .O(N__64582),
            .I(N__64573));
    InMux I__14866 (
            .O(N__64581),
            .I(N__64570));
    Odrv4 I__14865 (
            .O(N__64578),
            .I(\c0.n13523 ));
    Odrv4 I__14864 (
            .O(N__64573),
            .I(\c0.n13523 ));
    LocalMux I__14863 (
            .O(N__64570),
            .I(\c0.n13523 ));
    InMux I__14862 (
            .O(N__64563),
            .I(N__64557));
    InMux I__14861 (
            .O(N__64562),
            .I(N__64557));
    LocalMux I__14860 (
            .O(N__64557),
            .I(\c0.n47 ));
    CascadeMux I__14859 (
            .O(N__64554),
            .I(N__64551));
    InMux I__14858 (
            .O(N__64551),
            .I(N__64548));
    LocalMux I__14857 (
            .O(N__64548),
            .I(\c0.n10_adj_4664 ));
    InMux I__14856 (
            .O(N__64545),
            .I(N__64541));
    CascadeMux I__14855 (
            .O(N__64544),
            .I(N__64538));
    LocalMux I__14854 (
            .O(N__64541),
            .I(N__64535));
    InMux I__14853 (
            .O(N__64538),
            .I(N__64532));
    Span4Mux_v I__14852 (
            .O(N__64535),
            .I(N__64524));
    LocalMux I__14851 (
            .O(N__64532),
            .I(N__64524));
    InMux I__14850 (
            .O(N__64531),
            .I(N__64521));
    InMux I__14849 (
            .O(N__64530),
            .I(N__64516));
    InMux I__14848 (
            .O(N__64529),
            .I(N__64516));
    Span4Mux_v I__14847 (
            .O(N__64524),
            .I(N__64513));
    LocalMux I__14846 (
            .O(N__64521),
            .I(\c0.data_in_frame_9_2 ));
    LocalMux I__14845 (
            .O(N__64516),
            .I(\c0.data_in_frame_9_2 ));
    Odrv4 I__14844 (
            .O(N__64513),
            .I(\c0.data_in_frame_9_2 ));
    InMux I__14843 (
            .O(N__64506),
            .I(N__64503));
    LocalMux I__14842 (
            .O(N__64503),
            .I(N__64498));
    CascadeMux I__14841 (
            .O(N__64502),
            .I(N__64495));
    InMux I__14840 (
            .O(N__64501),
            .I(N__64492));
    Span4Mux_v I__14839 (
            .O(N__64498),
            .I(N__64487));
    InMux I__14838 (
            .O(N__64495),
            .I(N__64484));
    LocalMux I__14837 (
            .O(N__64492),
            .I(N__64481));
    InMux I__14836 (
            .O(N__64491),
            .I(N__64478));
    InMux I__14835 (
            .O(N__64490),
            .I(N__64475));
    Span4Mux_h I__14834 (
            .O(N__64487),
            .I(N__64472));
    LocalMux I__14833 (
            .O(N__64484),
            .I(N__64465));
    Span4Mux_v I__14832 (
            .O(N__64481),
            .I(N__64465));
    LocalMux I__14831 (
            .O(N__64478),
            .I(N__64465));
    LocalMux I__14830 (
            .O(N__64475),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__14829 (
            .O(N__64472),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__14828 (
            .O(N__64465),
            .I(\c0.data_in_frame_7_0 ));
    CascadeMux I__14827 (
            .O(N__64458),
            .I(N__64454));
    InMux I__14826 (
            .O(N__64457),
            .I(N__64451));
    InMux I__14825 (
            .O(N__64454),
            .I(N__64447));
    LocalMux I__14824 (
            .O(N__64451),
            .I(N__64444));
    CascadeMux I__14823 (
            .O(N__64450),
            .I(N__64441));
    LocalMux I__14822 (
            .O(N__64447),
            .I(N__64437));
    Span4Mux_h I__14821 (
            .O(N__64444),
            .I(N__64434));
    InMux I__14820 (
            .O(N__64441),
            .I(N__64431));
    InMux I__14819 (
            .O(N__64440),
            .I(N__64428));
    Span4Mux_v I__14818 (
            .O(N__64437),
            .I(N__64423));
    Span4Mux_h I__14817 (
            .O(N__64434),
            .I(N__64423));
    LocalMux I__14816 (
            .O(N__64431),
            .I(\c0.data_in_frame_7_5 ));
    LocalMux I__14815 (
            .O(N__64428),
            .I(\c0.data_in_frame_7_5 ));
    Odrv4 I__14814 (
            .O(N__64423),
            .I(\c0.data_in_frame_7_5 ));
    CascadeMux I__14813 (
            .O(N__64416),
            .I(\c0.n22417_cascade_ ));
    InMux I__14812 (
            .O(N__64413),
            .I(N__64410));
    LocalMux I__14811 (
            .O(N__64410),
            .I(N__64406));
    InMux I__14810 (
            .O(N__64409),
            .I(N__64403));
    Span4Mux_h I__14809 (
            .O(N__64406),
            .I(N__64400));
    LocalMux I__14808 (
            .O(N__64403),
            .I(N__64397));
    Span4Mux_h I__14807 (
            .O(N__64400),
            .I(N__64394));
    Odrv4 I__14806 (
            .O(N__64397),
            .I(\c0.n4_adj_4333 ));
    Odrv4 I__14805 (
            .O(N__64394),
            .I(\c0.n4_adj_4333 ));
    InMux I__14804 (
            .O(N__64389),
            .I(N__64386));
    LocalMux I__14803 (
            .O(N__64386),
            .I(N__64383));
    Span4Mux_h I__14802 (
            .O(N__64383),
            .I(N__64380));
    Odrv4 I__14801 (
            .O(N__64380),
            .I(\c0.n86 ));
    InMux I__14800 (
            .O(N__64377),
            .I(N__64374));
    LocalMux I__14799 (
            .O(N__64374),
            .I(N__64370));
    InMux I__14798 (
            .O(N__64373),
            .I(N__64367));
    Span4Mux_h I__14797 (
            .O(N__64370),
            .I(N__64364));
    LocalMux I__14796 (
            .O(N__64367),
            .I(N__64361));
    Span4Mux_h I__14795 (
            .O(N__64364),
            .I(N__64355));
    Span4Mux_v I__14794 (
            .O(N__64361),
            .I(N__64355));
    InMux I__14793 (
            .O(N__64360),
            .I(N__64352));
    Odrv4 I__14792 (
            .O(N__64355),
            .I(\c0.n13085 ));
    LocalMux I__14791 (
            .O(N__64352),
            .I(\c0.n13085 ));
    InMux I__14790 (
            .O(N__64347),
            .I(N__64342));
    InMux I__14789 (
            .O(N__64346),
            .I(N__64337));
    InMux I__14788 (
            .O(N__64345),
            .I(N__64334));
    LocalMux I__14787 (
            .O(N__64342),
            .I(N__64331));
    InMux I__14786 (
            .O(N__64341),
            .I(N__64328));
    InMux I__14785 (
            .O(N__64340),
            .I(N__64325));
    LocalMux I__14784 (
            .O(N__64337),
            .I(N__64322));
    LocalMux I__14783 (
            .O(N__64334),
            .I(N__64317));
    Span4Mux_h I__14782 (
            .O(N__64331),
            .I(N__64317));
    LocalMux I__14781 (
            .O(N__64328),
            .I(N__64314));
    LocalMux I__14780 (
            .O(N__64325),
            .I(N__64311));
    Span4Mux_v I__14779 (
            .O(N__64322),
            .I(N__64306));
    Span4Mux_v I__14778 (
            .O(N__64317),
            .I(N__64306));
    Span4Mux_h I__14777 (
            .O(N__64314),
            .I(N__64303));
    Span4Mux_v I__14776 (
            .O(N__64311),
            .I(N__64300));
    Odrv4 I__14775 (
            .O(N__64306),
            .I(\c0.n7_adj_4282 ));
    Odrv4 I__14774 (
            .O(N__64303),
            .I(\c0.n7_adj_4282 ));
    Odrv4 I__14773 (
            .O(N__64300),
            .I(\c0.n7_adj_4282 ));
    InMux I__14772 (
            .O(N__64293),
            .I(N__64290));
    LocalMux I__14771 (
            .O(N__64290),
            .I(\c0.n50 ));
    CascadeMux I__14770 (
            .O(N__64287),
            .I(n22121_cascade_));
    CascadeMux I__14769 (
            .O(N__64284),
            .I(N__64280));
    InMux I__14768 (
            .O(N__64283),
            .I(N__64275));
    InMux I__14767 (
            .O(N__64280),
            .I(N__64275));
    LocalMux I__14766 (
            .O(N__64275),
            .I(data_in_frame_6_6));
    InMux I__14765 (
            .O(N__64272),
            .I(N__64269));
    LocalMux I__14764 (
            .O(N__64269),
            .I(N__64266));
    Span4Mux_h I__14763 (
            .O(N__64266),
            .I(N__64263));
    Span4Mux_v I__14762 (
            .O(N__64263),
            .I(N__64256));
    InMux I__14761 (
            .O(N__64262),
            .I(N__64251));
    InMux I__14760 (
            .O(N__64261),
            .I(N__64251));
    InMux I__14759 (
            .O(N__64260),
            .I(N__64246));
    InMux I__14758 (
            .O(N__64259),
            .I(N__64246));
    Odrv4 I__14757 (
            .O(N__64256),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__14756 (
            .O(N__64251),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__14755 (
            .O(N__64246),
            .I(\c0.data_in_frame_2_2 ));
    CascadeMux I__14754 (
            .O(N__64239),
            .I(N__64236));
    InMux I__14753 (
            .O(N__64236),
            .I(N__64233));
    LocalMux I__14752 (
            .O(N__64233),
            .I(N__64230));
    Span4Mux_v I__14751 (
            .O(N__64230),
            .I(N__64226));
    CascadeMux I__14750 (
            .O(N__64229),
            .I(N__64223));
    Span4Mux_h I__14749 (
            .O(N__64226),
            .I(N__64220));
    InMux I__14748 (
            .O(N__64223),
            .I(N__64217));
    Odrv4 I__14747 (
            .O(N__64220),
            .I(\c0.n4_adj_4211 ));
    LocalMux I__14746 (
            .O(N__64217),
            .I(\c0.n4_adj_4211 ));
    InMux I__14745 (
            .O(N__64212),
            .I(N__64206));
    InMux I__14744 (
            .O(N__64211),
            .I(N__64206));
    LocalMux I__14743 (
            .O(N__64206),
            .I(\c0.n22647 ));
    CascadeMux I__14742 (
            .O(N__64203),
            .I(\c0.n13904_cascade_ ));
    InMux I__14741 (
            .O(N__64200),
            .I(N__64197));
    LocalMux I__14740 (
            .O(N__64197),
            .I(\c0.n21_adj_4327 ));
    CascadeMux I__14739 (
            .O(N__64194),
            .I(\c0.n19_adj_4324_cascade_ ));
    InMux I__14738 (
            .O(N__64191),
            .I(N__64188));
    LocalMux I__14737 (
            .O(N__64188),
            .I(N__64185));
    Span4Mux_h I__14736 (
            .O(N__64185),
            .I(N__64182));
    Odrv4 I__14735 (
            .O(N__64182),
            .I(\c0.n22417 ));
    CascadeMux I__14734 (
            .O(N__64179),
            .I(N__64174));
    InMux I__14733 (
            .O(N__64178),
            .I(N__64169));
    InMux I__14732 (
            .O(N__64177),
            .I(N__64169));
    InMux I__14731 (
            .O(N__64174),
            .I(N__64165));
    LocalMux I__14730 (
            .O(N__64169),
            .I(N__64162));
    CascadeMux I__14729 (
            .O(N__64168),
            .I(N__64159));
    LocalMux I__14728 (
            .O(N__64165),
            .I(N__64153));
    Span4Mux_v I__14727 (
            .O(N__64162),
            .I(N__64153));
    InMux I__14726 (
            .O(N__64159),
            .I(N__64148));
    InMux I__14725 (
            .O(N__64158),
            .I(N__64148));
    Odrv4 I__14724 (
            .O(N__64153),
            .I(\c0.data_in_frame_24_1 ));
    LocalMux I__14723 (
            .O(N__64148),
            .I(\c0.data_in_frame_24_1 ));
    InMux I__14722 (
            .O(N__64143),
            .I(N__64140));
    LocalMux I__14721 (
            .O(N__64140),
            .I(N__64135));
    CascadeMux I__14720 (
            .O(N__64139),
            .I(N__64130));
    InMux I__14719 (
            .O(N__64138),
            .I(N__64127));
    Span4Mux_v I__14718 (
            .O(N__64135),
            .I(N__64124));
    InMux I__14717 (
            .O(N__64134),
            .I(N__64121));
    InMux I__14716 (
            .O(N__64133),
            .I(N__64118));
    InMux I__14715 (
            .O(N__64130),
            .I(N__64115));
    LocalMux I__14714 (
            .O(N__64127),
            .I(N__64112));
    Sp12to4 I__14713 (
            .O(N__64124),
            .I(N__64107));
    LocalMux I__14712 (
            .O(N__64121),
            .I(N__64107));
    LocalMux I__14711 (
            .O(N__64118),
            .I(N__64104));
    LocalMux I__14710 (
            .O(N__64115),
            .I(N__64099));
    Span4Mux_h I__14709 (
            .O(N__64112),
            .I(N__64099));
    Span12Mux_h I__14708 (
            .O(N__64107),
            .I(N__64096));
    Odrv12 I__14707 (
            .O(N__64104),
            .I(\c0.data_in_frame_27_1 ));
    Odrv4 I__14706 (
            .O(N__64099),
            .I(\c0.data_in_frame_27_1 ));
    Odrv12 I__14705 (
            .O(N__64096),
            .I(\c0.data_in_frame_27_1 ));
    InMux I__14704 (
            .O(N__64089),
            .I(N__64086));
    LocalMux I__14703 (
            .O(N__64086),
            .I(N__64082));
    InMux I__14702 (
            .O(N__64085),
            .I(N__64079));
    Span4Mux_h I__14701 (
            .O(N__64082),
            .I(N__64076));
    LocalMux I__14700 (
            .O(N__64079),
            .I(N__64073));
    Odrv4 I__14699 (
            .O(N__64076),
            .I(\c0.n39_adj_4515 ));
    Odrv4 I__14698 (
            .O(N__64073),
            .I(\c0.n39_adj_4515 ));
    InMux I__14697 (
            .O(N__64068),
            .I(N__64065));
    LocalMux I__14696 (
            .O(N__64065),
            .I(N__64062));
    Odrv4 I__14695 (
            .O(N__64062),
            .I(\c0.n10_adj_4675 ));
    CascadeMux I__14694 (
            .O(N__64059),
            .I(N__64056));
    InMux I__14693 (
            .O(N__64056),
            .I(N__64053));
    LocalMux I__14692 (
            .O(N__64053),
            .I(N__64050));
    Span4Mux_v I__14691 (
            .O(N__64050),
            .I(N__64045));
    InMux I__14690 (
            .O(N__64049),
            .I(N__64042));
    CascadeMux I__14689 (
            .O(N__64048),
            .I(N__64039));
    Span4Mux_v I__14688 (
            .O(N__64045),
            .I(N__64034));
    LocalMux I__14687 (
            .O(N__64042),
            .I(N__64034));
    InMux I__14686 (
            .O(N__64039),
            .I(N__64030));
    Span4Mux_h I__14685 (
            .O(N__64034),
            .I(N__64027));
    InMux I__14684 (
            .O(N__64033),
            .I(N__64024));
    LocalMux I__14683 (
            .O(N__64030),
            .I(\c0.data_in_frame_11_0 ));
    Odrv4 I__14682 (
            .O(N__64027),
            .I(\c0.data_in_frame_11_0 ));
    LocalMux I__14681 (
            .O(N__64024),
            .I(\c0.data_in_frame_11_0 ));
    InMux I__14680 (
            .O(N__64017),
            .I(N__64014));
    LocalMux I__14679 (
            .O(N__64014),
            .I(N__64009));
    CascadeMux I__14678 (
            .O(N__64013),
            .I(N__64003));
    InMux I__14677 (
            .O(N__64012),
            .I(N__64000));
    Span4Mux_h I__14676 (
            .O(N__64009),
            .I(N__63997));
    InMux I__14675 (
            .O(N__64008),
            .I(N__63994));
    InMux I__14674 (
            .O(N__64007),
            .I(N__63989));
    InMux I__14673 (
            .O(N__64006),
            .I(N__63989));
    InMux I__14672 (
            .O(N__64003),
            .I(N__63986));
    LocalMux I__14671 (
            .O(N__64000),
            .I(N__63983));
    Odrv4 I__14670 (
            .O(N__63997),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__14669 (
            .O(N__63994),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__14668 (
            .O(N__63989),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__14667 (
            .O(N__63986),
            .I(\c0.data_in_frame_4_6 ));
    Odrv4 I__14666 (
            .O(N__63983),
            .I(\c0.data_in_frame_4_6 ));
    InMux I__14665 (
            .O(N__63972),
            .I(N__63969));
    LocalMux I__14664 (
            .O(N__63969),
            .I(N__63966));
    Span4Mux_h I__14663 (
            .O(N__63966),
            .I(N__63962));
    InMux I__14662 (
            .O(N__63965),
            .I(N__63958));
    Span4Mux_h I__14661 (
            .O(N__63962),
            .I(N__63955));
    InMux I__14660 (
            .O(N__63961),
            .I(N__63952));
    LocalMux I__14659 (
            .O(N__63958),
            .I(\c0.data_in_frame_23_7 ));
    Odrv4 I__14658 (
            .O(N__63955),
            .I(\c0.data_in_frame_23_7 ));
    LocalMux I__14657 (
            .O(N__63952),
            .I(\c0.data_in_frame_23_7 ));
    CascadeMux I__14656 (
            .O(N__63945),
            .I(\c0.n7_adj_4364_cascade_ ));
    InMux I__14655 (
            .O(N__63942),
            .I(N__63939));
    LocalMux I__14654 (
            .O(N__63939),
            .I(N__63936));
    Span4Mux_h I__14653 (
            .O(N__63936),
            .I(N__63933));
    Span4Mux_h I__14652 (
            .O(N__63933),
            .I(N__63929));
    InMux I__14651 (
            .O(N__63932),
            .I(N__63926));
    Odrv4 I__14650 (
            .O(N__63929),
            .I(\c0.n21426 ));
    LocalMux I__14649 (
            .O(N__63926),
            .I(\c0.n21426 ));
    CascadeMux I__14648 (
            .O(N__63921),
            .I(\c0.n23031_cascade_ ));
    InMux I__14647 (
            .O(N__63918),
            .I(N__63914));
    CascadeMux I__14646 (
            .O(N__63917),
            .I(N__63911));
    LocalMux I__14645 (
            .O(N__63914),
            .I(N__63908));
    InMux I__14644 (
            .O(N__63911),
            .I(N__63903));
    Span4Mux_v I__14643 (
            .O(N__63908),
            .I(N__63900));
    InMux I__14642 (
            .O(N__63907),
            .I(N__63895));
    InMux I__14641 (
            .O(N__63906),
            .I(N__63895));
    LocalMux I__14640 (
            .O(N__63903),
            .I(\c0.data_in_frame_25_7 ));
    Odrv4 I__14639 (
            .O(N__63900),
            .I(\c0.data_in_frame_25_7 ));
    LocalMux I__14638 (
            .O(N__63895),
            .I(\c0.data_in_frame_25_7 ));
    CascadeMux I__14637 (
            .O(N__63888),
            .I(N__63885));
    InMux I__14636 (
            .O(N__63885),
            .I(N__63882));
    LocalMux I__14635 (
            .O(N__63882),
            .I(N__63879));
    Span4Mux_h I__14634 (
            .O(N__63879),
            .I(N__63874));
    CascadeMux I__14633 (
            .O(N__63878),
            .I(N__63871));
    CascadeMux I__14632 (
            .O(N__63877),
            .I(N__63868));
    Span4Mux_h I__14631 (
            .O(N__63874),
            .I(N__63865));
    InMux I__14630 (
            .O(N__63871),
            .I(N__63860));
    InMux I__14629 (
            .O(N__63868),
            .I(N__63860));
    Odrv4 I__14628 (
            .O(N__63865),
            .I(\c0.data_in_frame_26_5 ));
    LocalMux I__14627 (
            .O(N__63860),
            .I(\c0.data_in_frame_26_5 ));
    InMux I__14626 (
            .O(N__63855),
            .I(N__63852));
    LocalMux I__14625 (
            .O(N__63852),
            .I(\c0.n24482 ));
    InMux I__14624 (
            .O(N__63849),
            .I(N__63843));
    InMux I__14623 (
            .O(N__63848),
            .I(N__63838));
    InMux I__14622 (
            .O(N__63847),
            .I(N__63838));
    InMux I__14621 (
            .O(N__63846),
            .I(N__63835));
    LocalMux I__14620 (
            .O(N__63843),
            .I(\c0.n23031 ));
    LocalMux I__14619 (
            .O(N__63838),
            .I(\c0.n23031 ));
    LocalMux I__14618 (
            .O(N__63835),
            .I(\c0.n23031 ));
    CascadeMux I__14617 (
            .O(N__63828),
            .I(N__63825));
    InMux I__14616 (
            .O(N__63825),
            .I(N__63821));
    InMux I__14615 (
            .O(N__63824),
            .I(N__63818));
    LocalMux I__14614 (
            .O(N__63821),
            .I(\c0.data_in_frame_28_2 ));
    LocalMux I__14613 (
            .O(N__63818),
            .I(\c0.data_in_frame_28_2 ));
    CascadeMux I__14612 (
            .O(N__63813),
            .I(\c0.n36_adj_4460_cascade_ ));
    InMux I__14611 (
            .O(N__63810),
            .I(N__63807));
    LocalMux I__14610 (
            .O(N__63807),
            .I(\c0.n41_adj_4511 ));
    InMux I__14609 (
            .O(N__63804),
            .I(N__63798));
    InMux I__14608 (
            .O(N__63803),
            .I(N__63798));
    LocalMux I__14607 (
            .O(N__63798),
            .I(N__63795));
    Odrv4 I__14606 (
            .O(N__63795),
            .I(\c0.n6_adj_4459 ));
    InMux I__14605 (
            .O(N__63792),
            .I(N__63783));
    InMux I__14604 (
            .O(N__63791),
            .I(N__63779));
    InMux I__14603 (
            .O(N__63790),
            .I(N__63776));
    InMux I__14602 (
            .O(N__63789),
            .I(N__63771));
    InMux I__14601 (
            .O(N__63788),
            .I(N__63771));
    InMux I__14600 (
            .O(N__63787),
            .I(N__63768));
    InMux I__14599 (
            .O(N__63786),
            .I(N__63765));
    LocalMux I__14598 (
            .O(N__63783),
            .I(N__63762));
    InMux I__14597 (
            .O(N__63782),
            .I(N__63759));
    LocalMux I__14596 (
            .O(N__63779),
            .I(N__63750));
    LocalMux I__14595 (
            .O(N__63776),
            .I(N__63750));
    LocalMux I__14594 (
            .O(N__63771),
            .I(N__63750));
    LocalMux I__14593 (
            .O(N__63768),
            .I(N__63750));
    LocalMux I__14592 (
            .O(N__63765),
            .I(\c0.n22426 ));
    Odrv4 I__14591 (
            .O(N__63762),
            .I(\c0.n22426 ));
    LocalMux I__14590 (
            .O(N__63759),
            .I(\c0.n22426 ));
    Odrv4 I__14589 (
            .O(N__63750),
            .I(\c0.n22426 ));
    CascadeMux I__14588 (
            .O(N__63741),
            .I(N__63736));
    CascadeMux I__14587 (
            .O(N__63740),
            .I(N__63732));
    CascadeMux I__14586 (
            .O(N__63739),
            .I(N__63728));
    InMux I__14585 (
            .O(N__63736),
            .I(N__63724));
    InMux I__14584 (
            .O(N__63735),
            .I(N__63719));
    InMux I__14583 (
            .O(N__63732),
            .I(N__63719));
    CascadeMux I__14582 (
            .O(N__63731),
            .I(N__63716));
    InMux I__14581 (
            .O(N__63728),
            .I(N__63713));
    InMux I__14580 (
            .O(N__63727),
            .I(N__63710));
    LocalMux I__14579 (
            .O(N__63724),
            .I(N__63705));
    LocalMux I__14578 (
            .O(N__63719),
            .I(N__63705));
    InMux I__14577 (
            .O(N__63716),
            .I(N__63702));
    LocalMux I__14576 (
            .O(N__63713),
            .I(N__63697));
    LocalMux I__14575 (
            .O(N__63710),
            .I(N__63697));
    Span4Mux_h I__14574 (
            .O(N__63705),
            .I(N__63694));
    LocalMux I__14573 (
            .O(N__63702),
            .I(\c0.data_in_frame_26_1 ));
    Odrv4 I__14572 (
            .O(N__63697),
            .I(\c0.data_in_frame_26_1 ));
    Odrv4 I__14571 (
            .O(N__63694),
            .I(\c0.data_in_frame_26_1 ));
    CascadeMux I__14570 (
            .O(N__63687),
            .I(N__63681));
    InMux I__14569 (
            .O(N__63686),
            .I(N__63677));
    InMux I__14568 (
            .O(N__63685),
            .I(N__63672));
    InMux I__14567 (
            .O(N__63684),
            .I(N__63672));
    InMux I__14566 (
            .O(N__63681),
            .I(N__63669));
    InMux I__14565 (
            .O(N__63680),
            .I(N__63666));
    LocalMux I__14564 (
            .O(N__63677),
            .I(\c0.n22340 ));
    LocalMux I__14563 (
            .O(N__63672),
            .I(\c0.n22340 ));
    LocalMux I__14562 (
            .O(N__63669),
            .I(\c0.n22340 ));
    LocalMux I__14561 (
            .O(N__63666),
            .I(\c0.n22340 ));
    CascadeMux I__14560 (
            .O(N__63657),
            .I(\c0.n5_adj_4472_cascade_ ));
    InMux I__14559 (
            .O(N__63654),
            .I(N__63650));
    InMux I__14558 (
            .O(N__63653),
            .I(N__63647));
    LocalMux I__14557 (
            .O(N__63650),
            .I(\c0.n21010 ));
    LocalMux I__14556 (
            .O(N__63647),
            .I(\c0.n21010 ));
    InMux I__14555 (
            .O(N__63642),
            .I(N__63639));
    LocalMux I__14554 (
            .O(N__63639),
            .I(\c0.n24_adj_4496 ));
    InMux I__14553 (
            .O(N__63636),
            .I(N__63631));
    InMux I__14552 (
            .O(N__63635),
            .I(N__63626));
    InMux I__14551 (
            .O(N__63634),
            .I(N__63626));
    LocalMux I__14550 (
            .O(N__63631),
            .I(\c0.n34_adj_4361 ));
    LocalMux I__14549 (
            .O(N__63626),
            .I(\c0.n34_adj_4361 ));
    CascadeMux I__14548 (
            .O(N__63621),
            .I(\c0.n57_cascade_ ));
    InMux I__14547 (
            .O(N__63618),
            .I(N__63615));
    LocalMux I__14546 (
            .O(N__63615),
            .I(\c0.n48_adj_4365 ));
    CascadeMux I__14545 (
            .O(N__63612),
            .I(\c0.n21426_cascade_ ));
    InMux I__14544 (
            .O(N__63609),
            .I(N__63606));
    LocalMux I__14543 (
            .O(N__63606),
            .I(N__63603));
    Span4Mux_h I__14542 (
            .O(N__63603),
            .I(N__63600));
    Span4Mux_h I__14541 (
            .O(N__63600),
            .I(N__63595));
    InMux I__14540 (
            .O(N__63599),
            .I(N__63592));
    InMux I__14539 (
            .O(N__63598),
            .I(N__63589));
    Odrv4 I__14538 (
            .O(N__63595),
            .I(\c0.n23032 ));
    LocalMux I__14537 (
            .O(N__63592),
            .I(\c0.n23032 ));
    LocalMux I__14536 (
            .O(N__63589),
            .I(\c0.n23032 ));
    CascadeMux I__14535 (
            .O(N__63582),
            .I(\c0.n23032_cascade_ ));
    InMux I__14534 (
            .O(N__63579),
            .I(N__63576));
    LocalMux I__14533 (
            .O(N__63576),
            .I(N__63573));
    Odrv4 I__14532 (
            .O(N__63573),
            .I(\c0.n25456 ));
    CascadeMux I__14531 (
            .O(N__63570),
            .I(\c0.n23209_cascade_ ));
    InMux I__14530 (
            .O(N__63567),
            .I(N__63564));
    LocalMux I__14529 (
            .O(N__63564),
            .I(\c0.n56_adj_4479 ));
    InMux I__14528 (
            .O(N__63561),
            .I(N__63557));
    InMux I__14527 (
            .O(N__63560),
            .I(N__63554));
    LocalMux I__14526 (
            .O(N__63557),
            .I(N__63551));
    LocalMux I__14525 (
            .O(N__63554),
            .I(N__63548));
    Odrv12 I__14524 (
            .O(N__63551),
            .I(\c0.n21299 ));
    Odrv12 I__14523 (
            .O(N__63548),
            .I(\c0.n21299 ));
    InMux I__14522 (
            .O(N__63543),
            .I(N__63539));
    InMux I__14521 (
            .O(N__63542),
            .I(N__63536));
    LocalMux I__14520 (
            .O(N__63539),
            .I(N__63533));
    LocalMux I__14519 (
            .O(N__63536),
            .I(N__63530));
    Span4Mux_h I__14518 (
            .O(N__63533),
            .I(N__63527));
    Span4Mux_v I__14517 (
            .O(N__63530),
            .I(N__63524));
    Span4Mux_v I__14516 (
            .O(N__63527),
            .I(N__63517));
    Span4Mux_h I__14515 (
            .O(N__63524),
            .I(N__63517));
    InMux I__14514 (
            .O(N__63523),
            .I(N__63512));
    InMux I__14513 (
            .O(N__63522),
            .I(N__63512));
    Odrv4 I__14512 (
            .O(N__63517),
            .I(data_in_frame_22_6));
    LocalMux I__14511 (
            .O(N__63512),
            .I(data_in_frame_22_6));
    InMux I__14510 (
            .O(N__63507),
            .I(N__63503));
    InMux I__14509 (
            .O(N__63506),
            .I(N__63500));
    LocalMux I__14508 (
            .O(N__63503),
            .I(N__63496));
    LocalMux I__14507 (
            .O(N__63500),
            .I(N__63493));
    InMux I__14506 (
            .O(N__63499),
            .I(N__63490));
    Span4Mux_h I__14505 (
            .O(N__63496),
            .I(N__63487));
    Span4Mux_h I__14504 (
            .O(N__63493),
            .I(N__63484));
    LocalMux I__14503 (
            .O(N__63490),
            .I(N__63479));
    Span4Mux_h I__14502 (
            .O(N__63487),
            .I(N__63479));
    Odrv4 I__14501 (
            .O(N__63484),
            .I(data_in_frame_22_0));
    Odrv4 I__14500 (
            .O(N__63479),
            .I(data_in_frame_22_0));
    CascadeMux I__14499 (
            .O(N__63474),
            .I(\c0.n12559_cascade_ ));
    InMux I__14498 (
            .O(N__63471),
            .I(N__63468));
    LocalMux I__14497 (
            .O(N__63468),
            .I(N__63465));
    Span12Mux_v I__14496 (
            .O(N__63465),
            .I(N__63461));
    InMux I__14495 (
            .O(N__63464),
            .I(N__63458));
    Odrv12 I__14494 (
            .O(N__63461),
            .I(\c0.n22375 ));
    LocalMux I__14493 (
            .O(N__63458),
            .I(\c0.n22375 ));
    InMux I__14492 (
            .O(N__63453),
            .I(N__63450));
    LocalMux I__14491 (
            .O(N__63450),
            .I(N__63447));
    Span4Mux_h I__14490 (
            .O(N__63447),
            .I(N__63444));
    Odrv4 I__14489 (
            .O(N__63444),
            .I(\c0.n24451 ));
    CascadeMux I__14488 (
            .O(N__63441),
            .I(N__63437));
    InMux I__14487 (
            .O(N__63440),
            .I(N__63434));
    InMux I__14486 (
            .O(N__63437),
            .I(N__63431));
    LocalMux I__14485 (
            .O(N__63434),
            .I(N__63427));
    LocalMux I__14484 (
            .O(N__63431),
            .I(N__63424));
    InMux I__14483 (
            .O(N__63430),
            .I(N__63421));
    Span4Mux_h I__14482 (
            .O(N__63427),
            .I(N__63418));
    Span4Mux_h I__14481 (
            .O(N__63424),
            .I(N__63413));
    LocalMux I__14480 (
            .O(N__63421),
            .I(N__63413));
    Span4Mux_h I__14479 (
            .O(N__63418),
            .I(N__63409));
    Span4Mux_v I__14478 (
            .O(N__63413),
            .I(N__63406));
    CascadeMux I__14477 (
            .O(N__63412),
            .I(N__63403));
    Sp12to4 I__14476 (
            .O(N__63409),
            .I(N__63400));
    Span4Mux_h I__14475 (
            .O(N__63406),
            .I(N__63397));
    InMux I__14474 (
            .O(N__63403),
            .I(N__63394));
    Span12Mux_v I__14473 (
            .O(N__63400),
            .I(N__63391));
    Span4Mux_v I__14472 (
            .O(N__63397),
            .I(N__63388));
    LocalMux I__14471 (
            .O(N__63394),
            .I(\c0.data_in_frame_19_1 ));
    Odrv12 I__14470 (
            .O(N__63391),
            .I(\c0.data_in_frame_19_1 ));
    Odrv4 I__14469 (
            .O(N__63388),
            .I(\c0.data_in_frame_19_1 ));
    InMux I__14468 (
            .O(N__63381),
            .I(N__63375));
    InMux I__14467 (
            .O(N__63380),
            .I(N__63372));
    InMux I__14466 (
            .O(N__63379),
            .I(N__63367));
    InMux I__14465 (
            .O(N__63378),
            .I(N__63367));
    LocalMux I__14464 (
            .O(N__63375),
            .I(N__63364));
    LocalMux I__14463 (
            .O(N__63372),
            .I(N__63359));
    LocalMux I__14462 (
            .O(N__63367),
            .I(N__63359));
    Span4Mux_v I__14461 (
            .O(N__63364),
            .I(N__63356));
    Span4Mux_v I__14460 (
            .O(N__63359),
            .I(N__63353));
    Odrv4 I__14459 (
            .O(N__63356),
            .I(\c0.n6215 ));
    Odrv4 I__14458 (
            .O(N__63353),
            .I(\c0.n6215 ));
    CascadeMux I__14457 (
            .O(N__63348),
            .I(N__63342));
    InMux I__14456 (
            .O(N__63347),
            .I(N__63339));
    InMux I__14455 (
            .O(N__63346),
            .I(N__63332));
    InMux I__14454 (
            .O(N__63345),
            .I(N__63332));
    InMux I__14453 (
            .O(N__63342),
            .I(N__63332));
    LocalMux I__14452 (
            .O(N__63339),
            .I(N__63329));
    LocalMux I__14451 (
            .O(N__63332),
            .I(N__63325));
    Span4Mux_h I__14450 (
            .O(N__63329),
            .I(N__63322));
    InMux I__14449 (
            .O(N__63328),
            .I(N__63319));
    Sp12to4 I__14448 (
            .O(N__63325),
            .I(N__63316));
    Span4Mux_h I__14447 (
            .O(N__63322),
            .I(N__63313));
    LocalMux I__14446 (
            .O(N__63319),
            .I(\c0.data_in_frame_19_2 ));
    Odrv12 I__14445 (
            .O(N__63316),
            .I(\c0.data_in_frame_19_2 ));
    Odrv4 I__14444 (
            .O(N__63313),
            .I(\c0.data_in_frame_19_2 ));
    InMux I__14443 (
            .O(N__63306),
            .I(N__63303));
    LocalMux I__14442 (
            .O(N__63303),
            .I(N__63300));
    Span4Mux_h I__14441 (
            .O(N__63300),
            .I(N__63296));
    InMux I__14440 (
            .O(N__63299),
            .I(N__63292));
    Span4Mux_h I__14439 (
            .O(N__63296),
            .I(N__63289));
    InMux I__14438 (
            .O(N__63295),
            .I(N__63286));
    LocalMux I__14437 (
            .O(N__63292),
            .I(\c0.n21275 ));
    Odrv4 I__14436 (
            .O(N__63289),
            .I(\c0.n21275 ));
    LocalMux I__14435 (
            .O(N__63286),
            .I(\c0.n21275 ));
    CascadeMux I__14434 (
            .O(N__63279),
            .I(\c0.n21275_cascade_ ));
    InMux I__14433 (
            .O(N__63276),
            .I(N__63273));
    LocalMux I__14432 (
            .O(N__63273),
            .I(N__63270));
    Span4Mux_v I__14431 (
            .O(N__63270),
            .I(N__63267));
    Odrv4 I__14430 (
            .O(N__63267),
            .I(\c0.n14_adj_4440 ));
    InMux I__14429 (
            .O(N__63264),
            .I(N__63260));
    InMux I__14428 (
            .O(N__63263),
            .I(N__63257));
    LocalMux I__14427 (
            .O(N__63260),
            .I(N__63254));
    LocalMux I__14426 (
            .O(N__63257),
            .I(N__63251));
    Span4Mux_h I__14425 (
            .O(N__63254),
            .I(N__63246));
    Span4Mux_v I__14424 (
            .O(N__63251),
            .I(N__63246));
    Odrv4 I__14423 (
            .O(N__63246),
            .I(\c0.n63_adj_4516 ));
    InMux I__14422 (
            .O(N__63243),
            .I(N__63237));
    InMux I__14421 (
            .O(N__63242),
            .I(N__63234));
    InMux I__14420 (
            .O(N__63241),
            .I(N__63231));
    InMux I__14419 (
            .O(N__63240),
            .I(N__63227));
    LocalMux I__14418 (
            .O(N__63237),
            .I(N__63223));
    LocalMux I__14417 (
            .O(N__63234),
            .I(N__63218));
    LocalMux I__14416 (
            .O(N__63231),
            .I(N__63218));
    InMux I__14415 (
            .O(N__63230),
            .I(N__63215));
    LocalMux I__14414 (
            .O(N__63227),
            .I(N__63212));
    InMux I__14413 (
            .O(N__63226),
            .I(N__63208));
    Span4Mux_v I__14412 (
            .O(N__63223),
            .I(N__63203));
    Span4Mux_v I__14411 (
            .O(N__63218),
            .I(N__63203));
    LocalMux I__14410 (
            .O(N__63215),
            .I(N__63198));
    Span4Mux_v I__14409 (
            .O(N__63212),
            .I(N__63198));
    InMux I__14408 (
            .O(N__63211),
            .I(N__63195));
    LocalMux I__14407 (
            .O(N__63208),
            .I(N__63192));
    Span4Mux_h I__14406 (
            .O(N__63203),
            .I(N__63185));
    Span4Mux_h I__14405 (
            .O(N__63198),
            .I(N__63185));
    LocalMux I__14404 (
            .O(N__63195),
            .I(N__63185));
    Span4Mux_h I__14403 (
            .O(N__63192),
            .I(N__63182));
    Span4Mux_v I__14402 (
            .O(N__63185),
            .I(N__63179));
    Odrv4 I__14401 (
            .O(N__63182),
            .I(\c0.n14189 ));
    Odrv4 I__14400 (
            .O(N__63179),
            .I(\c0.n14189 ));
    CascadeMux I__14399 (
            .O(N__63174),
            .I(N__63171));
    InMux I__14398 (
            .O(N__63171),
            .I(N__63167));
    InMux I__14397 (
            .O(N__63170),
            .I(N__63164));
    LocalMux I__14396 (
            .O(N__63167),
            .I(\c0.n46 ));
    LocalMux I__14395 (
            .O(N__63164),
            .I(\c0.n46 ));
    CascadeMux I__14394 (
            .O(N__63159),
            .I(\c0.n46_cascade_ ));
    CascadeMux I__14393 (
            .O(N__63156),
            .I(N__63153));
    InMux I__14392 (
            .O(N__63153),
            .I(N__63149));
    InMux I__14391 (
            .O(N__63152),
            .I(N__63145));
    LocalMux I__14390 (
            .O(N__63149),
            .I(N__63142));
    InMux I__14389 (
            .O(N__63148),
            .I(N__63138));
    LocalMux I__14388 (
            .O(N__63145),
            .I(N__63135));
    Span4Mux_h I__14387 (
            .O(N__63142),
            .I(N__63132));
    InMux I__14386 (
            .O(N__63141),
            .I(N__63129));
    LocalMux I__14385 (
            .O(N__63138),
            .I(\c0.data_in_frame_12_7 ));
    Odrv4 I__14384 (
            .O(N__63135),
            .I(\c0.data_in_frame_12_7 ));
    Odrv4 I__14383 (
            .O(N__63132),
            .I(\c0.data_in_frame_12_7 ));
    LocalMux I__14382 (
            .O(N__63129),
            .I(\c0.data_in_frame_12_7 ));
    InMux I__14381 (
            .O(N__63120),
            .I(N__63117));
    LocalMux I__14380 (
            .O(N__63117),
            .I(\c0.n25_adj_4579 ));
    CascadeMux I__14379 (
            .O(N__63114),
            .I(\c0.n25_adj_4579_cascade_ ));
    CascadeMux I__14378 (
            .O(N__63111),
            .I(\c0.n23433_cascade_ ));
    InMux I__14377 (
            .O(N__63108),
            .I(N__63102));
    InMux I__14376 (
            .O(N__63107),
            .I(N__63102));
    LocalMux I__14375 (
            .O(N__63102),
            .I(N__63099));
    Odrv12 I__14374 (
            .O(N__63099),
            .I(\c0.n18_adj_4580 ));
    InMux I__14373 (
            .O(N__63096),
            .I(N__63093));
    LocalMux I__14372 (
            .O(N__63093),
            .I(\c0.n24_adj_4655 ));
    InMux I__14371 (
            .O(N__63090),
            .I(N__63086));
    CascadeMux I__14370 (
            .O(N__63089),
            .I(N__63083));
    LocalMux I__14369 (
            .O(N__63086),
            .I(N__63080));
    InMux I__14368 (
            .O(N__63083),
            .I(N__63077));
    Span4Mux_h I__14367 (
            .O(N__63080),
            .I(N__63074));
    LocalMux I__14366 (
            .O(N__63077),
            .I(\c0.n41_adj_4592 ));
    Odrv4 I__14365 (
            .O(N__63074),
            .I(\c0.n41_adj_4592 ));
    InMux I__14364 (
            .O(N__63069),
            .I(N__63066));
    LocalMux I__14363 (
            .O(N__63066),
            .I(\c0.n43_adj_4661 ));
    CascadeMux I__14362 (
            .O(N__63063),
            .I(N__63060));
    InMux I__14361 (
            .O(N__63060),
            .I(N__63057));
    LocalMux I__14360 (
            .O(N__63057),
            .I(N__63054));
    Odrv4 I__14359 (
            .O(N__63054),
            .I(\c0.n44_adj_4588 ));
    InMux I__14358 (
            .O(N__63051),
            .I(N__63048));
    LocalMux I__14357 (
            .O(N__63048),
            .I(N__63045));
    Span4Mux_h I__14356 (
            .O(N__63045),
            .I(N__63042));
    Odrv4 I__14355 (
            .O(N__63042),
            .I(\c0.n39_adj_4341 ));
    InMux I__14354 (
            .O(N__63039),
            .I(N__63036));
    LocalMux I__14353 (
            .O(N__63036),
            .I(N__63033));
    Span4Mux_v I__14352 (
            .O(N__63033),
            .I(N__63029));
    InMux I__14351 (
            .O(N__63032),
            .I(N__63026));
    Odrv4 I__14350 (
            .O(N__63029),
            .I(\c0.n22205 ));
    LocalMux I__14349 (
            .O(N__63026),
            .I(\c0.n22205 ));
    CascadeMux I__14348 (
            .O(N__63021),
            .I(\c0.n50_adj_4340_cascade_ ));
    InMux I__14347 (
            .O(N__63018),
            .I(N__63015));
    LocalMux I__14346 (
            .O(N__63015),
            .I(N__63012));
    Span4Mux_v I__14345 (
            .O(N__63012),
            .I(N__63008));
    InMux I__14344 (
            .O(N__63011),
            .I(N__63005));
    Span4Mux_h I__14343 (
            .O(N__63008),
            .I(N__63002));
    LocalMux I__14342 (
            .O(N__63005),
            .I(N__62999));
    Odrv4 I__14341 (
            .O(N__63002),
            .I(\c0.n5_adj_4486 ));
    Odrv4 I__14340 (
            .O(N__62999),
            .I(\c0.n5_adj_4486 ));
    InMux I__14339 (
            .O(N__62994),
            .I(N__62991));
    LocalMux I__14338 (
            .O(N__62991),
            .I(N__62988));
    Odrv4 I__14337 (
            .O(N__62988),
            .I(\c0.n20467 ));
    CascadeMux I__14336 (
            .O(N__62985),
            .I(\c0.n20467_cascade_ ));
    CascadeMux I__14335 (
            .O(N__62982),
            .I(N__62977));
    InMux I__14334 (
            .O(N__62981),
            .I(N__62974));
    CascadeMux I__14333 (
            .O(N__62980),
            .I(N__62971));
    InMux I__14332 (
            .O(N__62977),
            .I(N__62968));
    LocalMux I__14331 (
            .O(N__62974),
            .I(N__62965));
    InMux I__14330 (
            .O(N__62971),
            .I(N__62962));
    LocalMux I__14329 (
            .O(N__62968),
            .I(N__62959));
    Span4Mux_h I__14328 (
            .O(N__62965),
            .I(N__62956));
    LocalMux I__14327 (
            .O(N__62962),
            .I(N__62953));
    Span4Mux_v I__14326 (
            .O(N__62959),
            .I(N__62948));
    Span4Mux_v I__14325 (
            .O(N__62956),
            .I(N__62948));
    Odrv4 I__14324 (
            .O(N__62953),
            .I(\c0.n6404 ));
    Odrv4 I__14323 (
            .O(N__62948),
            .I(\c0.n6404 ));
    CascadeMux I__14322 (
            .O(N__62943),
            .I(\c0.n17_adj_4354_cascade_ ));
    InMux I__14321 (
            .O(N__62940),
            .I(N__62934));
    InMux I__14320 (
            .O(N__62939),
            .I(N__62934));
    LocalMux I__14319 (
            .O(N__62934),
            .I(\c0.n10_adj_4630 ));
    InMux I__14318 (
            .O(N__62931),
            .I(N__62928));
    LocalMux I__14317 (
            .O(N__62928),
            .I(N__62924));
    CascadeMux I__14316 (
            .O(N__62927),
            .I(N__62921));
    Span4Mux_h I__14315 (
            .O(N__62924),
            .I(N__62916));
    InMux I__14314 (
            .O(N__62921),
            .I(N__62911));
    InMux I__14313 (
            .O(N__62920),
            .I(N__62911));
    InMux I__14312 (
            .O(N__62919),
            .I(N__62908));
    Span4Mux_v I__14311 (
            .O(N__62916),
            .I(N__62905));
    LocalMux I__14310 (
            .O(N__62911),
            .I(N__62900));
    LocalMux I__14309 (
            .O(N__62908),
            .I(N__62900));
    Odrv4 I__14308 (
            .O(N__62905),
            .I(\c0.n23523 ));
    Odrv12 I__14307 (
            .O(N__62900),
            .I(\c0.n23523 ));
    InMux I__14306 (
            .O(N__62895),
            .I(N__62891));
    InMux I__14305 (
            .O(N__62894),
            .I(N__62888));
    LocalMux I__14304 (
            .O(N__62891),
            .I(N__62881));
    LocalMux I__14303 (
            .O(N__62888),
            .I(N__62881));
    InMux I__14302 (
            .O(N__62887),
            .I(N__62876));
    InMux I__14301 (
            .O(N__62886),
            .I(N__62876));
    Span4Mux_v I__14300 (
            .O(N__62881),
            .I(N__62872));
    LocalMux I__14299 (
            .O(N__62876),
            .I(N__62869));
    InMux I__14298 (
            .O(N__62875),
            .I(N__62866));
    Odrv4 I__14297 (
            .O(N__62872),
            .I(\c0.n6_adj_4209 ));
    Odrv12 I__14296 (
            .O(N__62869),
            .I(\c0.n6_adj_4209 ));
    LocalMux I__14295 (
            .O(N__62866),
            .I(\c0.n6_adj_4209 ));
    CascadeMux I__14294 (
            .O(N__62859),
            .I(N__62855));
    InMux I__14293 (
            .O(N__62858),
            .I(N__62849));
    InMux I__14292 (
            .O(N__62855),
            .I(N__62849));
    InMux I__14291 (
            .O(N__62854),
            .I(N__62844));
    LocalMux I__14290 (
            .O(N__62849),
            .I(N__62841));
    InMux I__14289 (
            .O(N__62848),
            .I(N__62838));
    CascadeMux I__14288 (
            .O(N__62847),
            .I(N__62835));
    LocalMux I__14287 (
            .O(N__62844),
            .I(N__62832));
    Span4Mux_v I__14286 (
            .O(N__62841),
            .I(N__62829));
    LocalMux I__14285 (
            .O(N__62838),
            .I(N__62826));
    InMux I__14284 (
            .O(N__62835),
            .I(N__62823));
    Span12Mux_v I__14283 (
            .O(N__62832),
            .I(N__62820));
    Span4Mux_v I__14282 (
            .O(N__62829),
            .I(N__62815));
    Span4Mux_h I__14281 (
            .O(N__62826),
            .I(N__62815));
    LocalMux I__14280 (
            .O(N__62823),
            .I(\c0.data_in_frame_13_7 ));
    Odrv12 I__14279 (
            .O(N__62820),
            .I(\c0.data_in_frame_13_7 ));
    Odrv4 I__14278 (
            .O(N__62815),
            .I(\c0.data_in_frame_13_7 ));
    InMux I__14277 (
            .O(N__62808),
            .I(N__62803));
    CascadeMux I__14276 (
            .O(N__62807),
            .I(N__62800));
    CascadeMux I__14275 (
            .O(N__62806),
            .I(N__62796));
    LocalMux I__14274 (
            .O(N__62803),
            .I(N__62792));
    InMux I__14273 (
            .O(N__62800),
            .I(N__62787));
    InMux I__14272 (
            .O(N__62799),
            .I(N__62787));
    InMux I__14271 (
            .O(N__62796),
            .I(N__62784));
    InMux I__14270 (
            .O(N__62795),
            .I(N__62781));
    Span4Mux_h I__14269 (
            .O(N__62792),
            .I(N__62774));
    LocalMux I__14268 (
            .O(N__62787),
            .I(N__62774));
    LocalMux I__14267 (
            .O(N__62784),
            .I(N__62774));
    LocalMux I__14266 (
            .O(N__62781),
            .I(\c0.data_in_frame_12_6 ));
    Odrv4 I__14265 (
            .O(N__62774),
            .I(\c0.data_in_frame_12_6 ));
    InMux I__14264 (
            .O(N__62769),
            .I(N__62759));
    InMux I__14263 (
            .O(N__62768),
            .I(N__62759));
    InMux I__14262 (
            .O(N__62767),
            .I(N__62759));
    InMux I__14261 (
            .O(N__62766),
            .I(N__62753));
    LocalMux I__14260 (
            .O(N__62759),
            .I(N__62750));
    InMux I__14259 (
            .O(N__62758),
            .I(N__62743));
    InMux I__14258 (
            .O(N__62757),
            .I(N__62743));
    InMux I__14257 (
            .O(N__62756),
            .I(N__62743));
    LocalMux I__14256 (
            .O(N__62753),
            .I(N__62735));
    Span4Mux_v I__14255 (
            .O(N__62750),
            .I(N__62735));
    LocalMux I__14254 (
            .O(N__62743),
            .I(N__62735));
    InMux I__14253 (
            .O(N__62742),
            .I(N__62732));
    Odrv4 I__14252 (
            .O(N__62735),
            .I(\c0.n22782 ));
    LocalMux I__14251 (
            .O(N__62732),
            .I(\c0.n22782 ));
    InMux I__14250 (
            .O(N__62727),
            .I(N__62724));
    LocalMux I__14249 (
            .O(N__62724),
            .I(\c0.n12_adj_4246 ));
    InMux I__14248 (
            .O(N__62721),
            .I(N__62715));
    InMux I__14247 (
            .O(N__62720),
            .I(N__62715));
    LocalMux I__14246 (
            .O(N__62715),
            .I(\c0.n23453 ));
    InMux I__14245 (
            .O(N__62712),
            .I(N__62705));
    InMux I__14244 (
            .O(N__62711),
            .I(N__62705));
    InMux I__14243 (
            .O(N__62710),
            .I(N__62702));
    LocalMux I__14242 (
            .O(N__62705),
            .I(N__62699));
    LocalMux I__14241 (
            .O(N__62702),
            .I(N__62696));
    Span4Mux_h I__14240 (
            .O(N__62699),
            .I(N__62693));
    Odrv4 I__14239 (
            .O(N__62696),
            .I(\c0.n22540 ));
    Odrv4 I__14238 (
            .O(N__62693),
            .I(\c0.n22540 ));
    InMux I__14237 (
            .O(N__62688),
            .I(N__62683));
    InMux I__14236 (
            .O(N__62687),
            .I(N__62677));
    InMux I__14235 (
            .O(N__62686),
            .I(N__62677));
    LocalMux I__14234 (
            .O(N__62683),
            .I(N__62674));
    InMux I__14233 (
            .O(N__62682),
            .I(N__62671));
    LocalMux I__14232 (
            .O(N__62677),
            .I(N__62668));
    Span4Mux_v I__14231 (
            .O(N__62674),
            .I(N__62663));
    LocalMux I__14230 (
            .O(N__62671),
            .I(N__62658));
    Span4Mux_h I__14229 (
            .O(N__62668),
            .I(N__62658));
    InMux I__14228 (
            .O(N__62667),
            .I(N__62655));
    InMux I__14227 (
            .O(N__62666),
            .I(N__62652));
    Odrv4 I__14226 (
            .O(N__62663),
            .I(\c0.n24333 ));
    Odrv4 I__14225 (
            .O(N__62658),
            .I(\c0.n24333 ));
    LocalMux I__14224 (
            .O(N__62655),
            .I(\c0.n24333 ));
    LocalMux I__14223 (
            .O(N__62652),
            .I(\c0.n24333 ));
    CascadeMux I__14222 (
            .O(N__62643),
            .I(N__62640));
    InMux I__14221 (
            .O(N__62640),
            .I(N__62635));
    InMux I__14220 (
            .O(N__62639),
            .I(N__62632));
    InMux I__14219 (
            .O(N__62638),
            .I(N__62629));
    LocalMux I__14218 (
            .O(N__62635),
            .I(N__62624));
    LocalMux I__14217 (
            .O(N__62632),
            .I(N__62624));
    LocalMux I__14216 (
            .O(N__62629),
            .I(N__62621));
    Odrv4 I__14215 (
            .O(N__62624),
            .I(\c0.n22822 ));
    Odrv4 I__14214 (
            .O(N__62621),
            .I(\c0.n22822 ));
    CascadeMux I__14213 (
            .O(N__62616),
            .I(N__62610));
    CascadeMux I__14212 (
            .O(N__62615),
            .I(N__62607));
    InMux I__14211 (
            .O(N__62614),
            .I(N__62604));
    InMux I__14210 (
            .O(N__62613),
            .I(N__62598));
    InMux I__14209 (
            .O(N__62610),
            .I(N__62598));
    InMux I__14208 (
            .O(N__62607),
            .I(N__62595));
    LocalMux I__14207 (
            .O(N__62604),
            .I(N__62592));
    CascadeMux I__14206 (
            .O(N__62603),
            .I(N__62588));
    LocalMux I__14205 (
            .O(N__62598),
            .I(N__62585));
    LocalMux I__14204 (
            .O(N__62595),
            .I(N__62582));
    Span4Mux_v I__14203 (
            .O(N__62592),
            .I(N__62579));
    InMux I__14202 (
            .O(N__62591),
            .I(N__62574));
    InMux I__14201 (
            .O(N__62588),
            .I(N__62574));
    Span4Mux_v I__14200 (
            .O(N__62585),
            .I(N__62571));
    Span4Mux_v I__14199 (
            .O(N__62582),
            .I(N__62566));
    Span4Mux_h I__14198 (
            .O(N__62579),
            .I(N__62566));
    LocalMux I__14197 (
            .O(N__62574),
            .I(data_in_frame_14_7));
    Odrv4 I__14196 (
            .O(N__62571),
            .I(data_in_frame_14_7));
    Odrv4 I__14195 (
            .O(N__62566),
            .I(data_in_frame_14_7));
    CascadeMux I__14194 (
            .O(N__62559),
            .I(\c0.n12_adj_4246_cascade_ ));
    CascadeMux I__14193 (
            .O(N__62556),
            .I(\c0.n23691_cascade_ ));
    InMux I__14192 (
            .O(N__62553),
            .I(N__62550));
    LocalMux I__14191 (
            .O(N__62550),
            .I(N__62546));
    InMux I__14190 (
            .O(N__62549),
            .I(N__62543));
    Span4Mux_v I__14189 (
            .O(N__62546),
            .I(N__62538));
    LocalMux I__14188 (
            .O(N__62543),
            .I(N__62538));
    Span4Mux_h I__14187 (
            .O(N__62538),
            .I(N__62535));
    Odrv4 I__14186 (
            .O(N__62535),
            .I(\c0.n20543 ));
    InMux I__14185 (
            .O(N__62532),
            .I(N__62529));
    LocalMux I__14184 (
            .O(N__62529),
            .I(N__62523));
    InMux I__14183 (
            .O(N__62528),
            .I(N__62518));
    InMux I__14182 (
            .O(N__62527),
            .I(N__62518));
    CascadeMux I__14181 (
            .O(N__62526),
            .I(N__62515));
    Span4Mux_h I__14180 (
            .O(N__62523),
            .I(N__62512));
    LocalMux I__14179 (
            .O(N__62518),
            .I(N__62509));
    InMux I__14178 (
            .O(N__62515),
            .I(N__62506));
    Span4Mux_h I__14177 (
            .O(N__62512),
            .I(N__62503));
    Span4Mux_v I__14176 (
            .O(N__62509),
            .I(N__62500));
    LocalMux I__14175 (
            .O(N__62506),
            .I(\c0.data_in_frame_16_5 ));
    Odrv4 I__14174 (
            .O(N__62503),
            .I(\c0.data_in_frame_16_5 ));
    Odrv4 I__14173 (
            .O(N__62500),
            .I(\c0.data_in_frame_16_5 ));
    InMux I__14172 (
            .O(N__62493),
            .I(N__62490));
    LocalMux I__14171 (
            .O(N__62490),
            .I(\c0.n10_adj_4602 ));
    InMux I__14170 (
            .O(N__62487),
            .I(N__62484));
    LocalMux I__14169 (
            .O(N__62484),
            .I(N__62480));
    InMux I__14168 (
            .O(N__62483),
            .I(N__62477));
    Span4Mux_h I__14167 (
            .O(N__62480),
            .I(N__62471));
    LocalMux I__14166 (
            .O(N__62477),
            .I(N__62471));
    InMux I__14165 (
            .O(N__62476),
            .I(N__62468));
    Odrv4 I__14164 (
            .O(N__62471),
            .I(\c0.n22644 ));
    LocalMux I__14163 (
            .O(N__62468),
            .I(\c0.n22644 ));
    InMux I__14162 (
            .O(N__62463),
            .I(N__62460));
    LocalMux I__14161 (
            .O(N__62460),
            .I(N__62455));
    CascadeMux I__14160 (
            .O(N__62459),
            .I(N__62452));
    InMux I__14159 (
            .O(N__62458),
            .I(N__62449));
    Span4Mux_h I__14158 (
            .O(N__62455),
            .I(N__62446));
    InMux I__14157 (
            .O(N__62452),
            .I(N__62442));
    LocalMux I__14156 (
            .O(N__62449),
            .I(N__62439));
    Span4Mux_h I__14155 (
            .O(N__62446),
            .I(N__62436));
    InMux I__14154 (
            .O(N__62445),
            .I(N__62433));
    LocalMux I__14153 (
            .O(N__62442),
            .I(\c0.data_in_frame_15_1 ));
    Odrv4 I__14152 (
            .O(N__62439),
            .I(\c0.data_in_frame_15_1 ));
    Odrv4 I__14151 (
            .O(N__62436),
            .I(\c0.data_in_frame_15_1 ));
    LocalMux I__14150 (
            .O(N__62433),
            .I(\c0.data_in_frame_15_1 ));
    InMux I__14149 (
            .O(N__62424),
            .I(N__62420));
    InMux I__14148 (
            .O(N__62423),
            .I(N__62417));
    LocalMux I__14147 (
            .O(N__62420),
            .I(\c0.n14165 ));
    LocalMux I__14146 (
            .O(N__62417),
            .I(\c0.n14165 ));
    CascadeMux I__14145 (
            .O(N__62412),
            .I(N__62408));
    InMux I__14144 (
            .O(N__62411),
            .I(N__62404));
    InMux I__14143 (
            .O(N__62408),
            .I(N__62401));
    InMux I__14142 (
            .O(N__62407),
            .I(N__62398));
    LocalMux I__14141 (
            .O(N__62404),
            .I(N__62389));
    LocalMux I__14140 (
            .O(N__62401),
            .I(N__62389));
    LocalMux I__14139 (
            .O(N__62398),
            .I(N__62389));
    InMux I__14138 (
            .O(N__62397),
            .I(N__62386));
    InMux I__14137 (
            .O(N__62396),
            .I(N__62383));
    Span4Mux_v I__14136 (
            .O(N__62389),
            .I(N__62380));
    LocalMux I__14135 (
            .O(N__62386),
            .I(N__62376));
    LocalMux I__14134 (
            .O(N__62383),
            .I(N__62371));
    Span4Mux_h I__14133 (
            .O(N__62380),
            .I(N__62371));
    InMux I__14132 (
            .O(N__62379),
            .I(N__62368));
    Odrv4 I__14131 (
            .O(N__62376),
            .I(data_in_frame_14_5));
    Odrv4 I__14130 (
            .O(N__62371),
            .I(data_in_frame_14_5));
    LocalMux I__14129 (
            .O(N__62368),
            .I(data_in_frame_14_5));
    CascadeMux I__14128 (
            .O(N__62361),
            .I(N__62357));
    InMux I__14127 (
            .O(N__62360),
            .I(N__62350));
    InMux I__14126 (
            .O(N__62357),
            .I(N__62345));
    InMux I__14125 (
            .O(N__62356),
            .I(N__62345));
    InMux I__14124 (
            .O(N__62355),
            .I(N__62338));
    InMux I__14123 (
            .O(N__62354),
            .I(N__62338));
    InMux I__14122 (
            .O(N__62353),
            .I(N__62338));
    LocalMux I__14121 (
            .O(N__62350),
            .I(\c0.n24444 ));
    LocalMux I__14120 (
            .O(N__62345),
            .I(\c0.n24444 ));
    LocalMux I__14119 (
            .O(N__62338),
            .I(\c0.n24444 ));
    CascadeMux I__14118 (
            .O(N__62331),
            .I(N__62328));
    InMux I__14117 (
            .O(N__62328),
            .I(N__62325));
    LocalMux I__14116 (
            .O(N__62325),
            .I(N__62322));
    Odrv4 I__14115 (
            .O(N__62322),
            .I(\c0.n7_adj_4581 ));
    InMux I__14114 (
            .O(N__62319),
            .I(N__62313));
    InMux I__14113 (
            .O(N__62318),
            .I(N__62310));
    InMux I__14112 (
            .O(N__62317),
            .I(N__62306));
    InMux I__14111 (
            .O(N__62316),
            .I(N__62303));
    LocalMux I__14110 (
            .O(N__62313),
            .I(N__62300));
    LocalMux I__14109 (
            .O(N__62310),
            .I(N__62297));
    InMux I__14108 (
            .O(N__62309),
            .I(N__62291));
    LocalMux I__14107 (
            .O(N__62306),
            .I(N__62286));
    LocalMux I__14106 (
            .O(N__62303),
            .I(N__62286));
    Span4Mux_h I__14105 (
            .O(N__62300),
            .I(N__62281));
    Span4Mux_v I__14104 (
            .O(N__62297),
            .I(N__62281));
    InMux I__14103 (
            .O(N__62296),
            .I(N__62278));
    InMux I__14102 (
            .O(N__62295),
            .I(N__62275));
    InMux I__14101 (
            .O(N__62294),
            .I(N__62272));
    LocalMux I__14100 (
            .O(N__62291),
            .I(N__62268));
    Span4Mux_v I__14099 (
            .O(N__62286),
            .I(N__62265));
    Span4Mux_v I__14098 (
            .O(N__62281),
            .I(N__62262));
    LocalMux I__14097 (
            .O(N__62278),
            .I(N__62259));
    LocalMux I__14096 (
            .O(N__62275),
            .I(N__62254));
    LocalMux I__14095 (
            .O(N__62272),
            .I(N__62254));
    InMux I__14094 (
            .O(N__62271),
            .I(N__62250));
    Span4Mux_h I__14093 (
            .O(N__62268),
            .I(N__62245));
    Span4Mux_v I__14092 (
            .O(N__62265),
            .I(N__62245));
    Span4Mux_v I__14091 (
            .O(N__62262),
            .I(N__62241));
    Span4Mux_h I__14090 (
            .O(N__62259),
            .I(N__62236));
    Span4Mux_h I__14089 (
            .O(N__62254),
            .I(N__62236));
    InMux I__14088 (
            .O(N__62253),
            .I(N__62233));
    LocalMux I__14087 (
            .O(N__62250),
            .I(N__62228));
    Span4Mux_h I__14086 (
            .O(N__62245),
            .I(N__62228));
    InMux I__14085 (
            .O(N__62244),
            .I(N__62225));
    Span4Mux_v I__14084 (
            .O(N__62241),
            .I(N__62222));
    Span4Mux_v I__14083 (
            .O(N__62236),
            .I(N__62219));
    LocalMux I__14082 (
            .O(N__62233),
            .I(N__62216));
    Span4Mux_v I__14081 (
            .O(N__62228),
            .I(N__62213));
    LocalMux I__14080 (
            .O(N__62225),
            .I(N__62210));
    Span4Mux_v I__14079 (
            .O(N__62222),
            .I(N__62207));
    Span4Mux_v I__14078 (
            .O(N__62219),
            .I(N__62204));
    Span12Mux_v I__14077 (
            .O(N__62216),
            .I(N__62201));
    Span4Mux_v I__14076 (
            .O(N__62213),
            .I(N__62198));
    Span12Mux_h I__14075 (
            .O(N__62210),
            .I(N__62194));
    Span4Mux_h I__14074 (
            .O(N__62207),
            .I(N__62191));
    Span4Mux_v I__14073 (
            .O(N__62204),
            .I(N__62188));
    Span12Mux_v I__14072 (
            .O(N__62201),
            .I(N__62185));
    Span4Mux_v I__14071 (
            .O(N__62198),
            .I(N__62182));
    InMux I__14070 (
            .O(N__62197),
            .I(N__62179));
    Odrv12 I__14069 (
            .O(N__62194),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__14068 (
            .O(N__62191),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__14067 (
            .O(N__62188),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv12 I__14066 (
            .O(N__62185),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__14065 (
            .O(N__62182),
            .I(\c0.FRAME_MATCHER_i_3 ));
    LocalMux I__14064 (
            .O(N__62179),
            .I(\c0.FRAME_MATCHER_i_3 ));
    SRMux I__14063 (
            .O(N__62166),
            .I(N__62163));
    LocalMux I__14062 (
            .O(N__62163),
            .I(N__62160));
    Span12Mux_s5_v I__14061 (
            .O(N__62160),
            .I(N__62157));
    Span12Mux_v I__14060 (
            .O(N__62157),
            .I(N__62154));
    Odrv12 I__14059 (
            .O(N__62154),
            .I(\c0.n3_adj_4430 ));
    InMux I__14058 (
            .O(N__62151),
            .I(N__62148));
    LocalMux I__14057 (
            .O(N__62148),
            .I(N__62145));
    Odrv12 I__14056 (
            .O(N__62145),
            .I(\c0.n124 ));
    InMux I__14055 (
            .O(N__62142),
            .I(N__62136));
    InMux I__14054 (
            .O(N__62141),
            .I(N__62136));
    LocalMux I__14053 (
            .O(N__62136),
            .I(\c0.n10_adj_4247 ));
    InMux I__14052 (
            .O(N__62133),
            .I(N__62127));
    InMux I__14051 (
            .O(N__62132),
            .I(N__62127));
    LocalMux I__14050 (
            .O(N__62127),
            .I(\c0.n22547 ));
    InMux I__14049 (
            .O(N__62124),
            .I(N__62120));
    InMux I__14048 (
            .O(N__62123),
            .I(N__62116));
    LocalMux I__14047 (
            .O(N__62120),
            .I(N__62113));
    InMux I__14046 (
            .O(N__62119),
            .I(N__62110));
    LocalMux I__14045 (
            .O(N__62116),
            .I(N__62107));
    Span4Mux_v I__14044 (
            .O(N__62113),
            .I(N__62102));
    LocalMux I__14043 (
            .O(N__62110),
            .I(N__62102));
    Span4Mux_v I__14042 (
            .O(N__62107),
            .I(N__62099));
    Span4Mux_v I__14041 (
            .O(N__62102),
            .I(N__62096));
    Odrv4 I__14040 (
            .O(N__62099),
            .I(\c0.n13998 ));
    Odrv4 I__14039 (
            .O(N__62096),
            .I(\c0.n13998 ));
    InMux I__14038 (
            .O(N__62091),
            .I(N__62088));
    LocalMux I__14037 (
            .O(N__62088),
            .I(N__62085));
    Span4Mux_v I__14036 (
            .O(N__62085),
            .I(N__62081));
    InMux I__14035 (
            .O(N__62084),
            .I(N__62078));
    Span4Mux_v I__14034 (
            .O(N__62081),
            .I(N__62075));
    LocalMux I__14033 (
            .O(N__62078),
            .I(N__62072));
    Span4Mux_h I__14032 (
            .O(N__62075),
            .I(N__62064));
    Span4Mux_v I__14031 (
            .O(N__62072),
            .I(N__62064));
    InMux I__14030 (
            .O(N__62071),
            .I(N__62057));
    InMux I__14029 (
            .O(N__62070),
            .I(N__62057));
    InMux I__14028 (
            .O(N__62069),
            .I(N__62057));
    Odrv4 I__14027 (
            .O(N__62064),
            .I(\c0.n23156 ));
    LocalMux I__14026 (
            .O(N__62057),
            .I(\c0.n23156 ));
    InMux I__14025 (
            .O(N__62052),
            .I(N__62049));
    LocalMux I__14024 (
            .O(N__62049),
            .I(N__62046));
    Span4Mux_v I__14023 (
            .O(N__62046),
            .I(N__62043));
    Span4Mux_h I__14022 (
            .O(N__62043),
            .I(N__62040));
    Odrv4 I__14021 (
            .O(N__62040),
            .I(\c0.n65 ));
    InMux I__14020 (
            .O(N__62037),
            .I(N__62034));
    LocalMux I__14019 (
            .O(N__62034),
            .I(N__62030));
    InMux I__14018 (
            .O(N__62033),
            .I(N__62027));
    Odrv12 I__14017 (
            .O(N__62030),
            .I(\c0.n60 ));
    LocalMux I__14016 (
            .O(N__62027),
            .I(\c0.n60 ));
    CascadeMux I__14015 (
            .O(N__62022),
            .I(\c0.n59_cascade_ ));
    InMux I__14014 (
            .O(N__62019),
            .I(N__62016));
    LocalMux I__14013 (
            .O(N__62016),
            .I(\c0.n70 ));
    CascadeMux I__14012 (
            .O(N__62013),
            .I(\c0.n24444_cascade_ ));
    InMux I__14011 (
            .O(N__62010),
            .I(N__62006));
    InMux I__14010 (
            .O(N__62009),
            .I(N__62003));
    LocalMux I__14009 (
            .O(N__62006),
            .I(N__62000));
    LocalMux I__14008 (
            .O(N__62003),
            .I(\c0.n21282 ));
    Odrv4 I__14007 (
            .O(N__62000),
            .I(\c0.n21282 ));
    InMux I__14006 (
            .O(N__61995),
            .I(N__61992));
    LocalMux I__14005 (
            .O(N__61992),
            .I(N__61988));
    CascadeMux I__14004 (
            .O(N__61991),
            .I(N__61984));
    Span4Mux_h I__14003 (
            .O(N__61988),
            .I(N__61981));
    CascadeMux I__14002 (
            .O(N__61987),
            .I(N__61978));
    InMux I__14001 (
            .O(N__61984),
            .I(N__61975));
    Span4Mux_v I__14000 (
            .O(N__61981),
            .I(N__61972));
    InMux I__13999 (
            .O(N__61978),
            .I(N__61969));
    LocalMux I__13998 (
            .O(N__61975),
            .I(\c0.data_in_frame_15_7 ));
    Odrv4 I__13997 (
            .O(N__61972),
            .I(\c0.data_in_frame_15_7 ));
    LocalMux I__13996 (
            .O(N__61969),
            .I(\c0.data_in_frame_15_7 ));
    CascadeMux I__13995 (
            .O(N__61962),
            .I(N__61959));
    InMux I__13994 (
            .O(N__61959),
            .I(N__61956));
    LocalMux I__13993 (
            .O(N__61956),
            .I(N__61953));
    Span4Mux_h I__13992 (
            .O(N__61953),
            .I(N__61950));
    Span4Mux_h I__13991 (
            .O(N__61950),
            .I(N__61946));
    InMux I__13990 (
            .O(N__61949),
            .I(N__61943));
    Odrv4 I__13989 (
            .O(N__61946),
            .I(\c0.n22514 ));
    LocalMux I__13988 (
            .O(N__61943),
            .I(\c0.n22514 ));
    CascadeMux I__13987 (
            .O(N__61938),
            .I(\c0.n23224_cascade_ ));
    InMux I__13986 (
            .O(N__61935),
            .I(N__61931));
    InMux I__13985 (
            .O(N__61934),
            .I(N__61928));
    LocalMux I__13984 (
            .O(N__61931),
            .I(N__61921));
    LocalMux I__13983 (
            .O(N__61928),
            .I(N__61921));
    InMux I__13982 (
            .O(N__61927),
            .I(N__61916));
    InMux I__13981 (
            .O(N__61926),
            .I(N__61916));
    Span4Mux_v I__13980 (
            .O(N__61921),
            .I(N__61913));
    LocalMux I__13979 (
            .O(N__61916),
            .I(N__61910));
    Span4Mux_h I__13978 (
            .O(N__61913),
            .I(N__61905));
    Span4Mux_v I__13977 (
            .O(N__61910),
            .I(N__61905));
    Odrv4 I__13976 (
            .O(N__61905),
            .I(\c0.n21409 ));
    InMux I__13975 (
            .O(N__61902),
            .I(N__61898));
    InMux I__13974 (
            .O(N__61901),
            .I(N__61894));
    LocalMux I__13973 (
            .O(N__61898),
            .I(N__61891));
    CascadeMux I__13972 (
            .O(N__61897),
            .I(N__61887));
    LocalMux I__13971 (
            .O(N__61894),
            .I(N__61884));
    Span4Mux_v I__13970 (
            .O(N__61891),
            .I(N__61881));
    InMux I__13969 (
            .O(N__61890),
            .I(N__61878));
    InMux I__13968 (
            .O(N__61887),
            .I(N__61875));
    Span4Mux_h I__13967 (
            .O(N__61884),
            .I(N__61872));
    Sp12to4 I__13966 (
            .O(N__61881),
            .I(N__61867));
    LocalMux I__13965 (
            .O(N__61878),
            .I(N__61867));
    LocalMux I__13964 (
            .O(N__61875),
            .I(\c0.data_in_frame_18_6 ));
    Odrv4 I__13963 (
            .O(N__61872),
            .I(\c0.data_in_frame_18_6 ));
    Odrv12 I__13962 (
            .O(N__61867),
            .I(\c0.data_in_frame_18_6 ));
    InMux I__13961 (
            .O(N__61860),
            .I(N__61856));
    InMux I__13960 (
            .O(N__61859),
            .I(N__61853));
    LocalMux I__13959 (
            .O(N__61856),
            .I(N__61846));
    LocalMux I__13958 (
            .O(N__61853),
            .I(N__61846));
    InMux I__13957 (
            .O(N__61852),
            .I(N__61841));
    InMux I__13956 (
            .O(N__61851),
            .I(N__61841));
    Span4Mux_h I__13955 (
            .O(N__61846),
            .I(N__61838));
    LocalMux I__13954 (
            .O(N__61841),
            .I(\c0.n13128 ));
    Odrv4 I__13953 (
            .O(N__61838),
            .I(\c0.n13128 ));
    CascadeMux I__13952 (
            .O(N__61833),
            .I(N__61830));
    InMux I__13951 (
            .O(N__61830),
            .I(N__61827));
    LocalMux I__13950 (
            .O(N__61827),
            .I(N__61824));
    Span4Mux_v I__13949 (
            .O(N__61824),
            .I(N__61821));
    Span4Mux_v I__13948 (
            .O(N__61821),
            .I(N__61818));
    Odrv4 I__13947 (
            .O(N__61818),
            .I(\c0.n7_adj_4603 ));
    InMux I__13946 (
            .O(N__61815),
            .I(N__61812));
    LocalMux I__13945 (
            .O(N__61812),
            .I(N__61808));
    InMux I__13944 (
            .O(N__61811),
            .I(N__61805));
    Odrv4 I__13943 (
            .O(N__61808),
            .I(\c0.n22589 ));
    LocalMux I__13942 (
            .O(N__61805),
            .I(\c0.n22589 ));
    CascadeMux I__13941 (
            .O(N__61800),
            .I(\c0.n13738_cascade_ ));
    InMux I__13940 (
            .O(N__61797),
            .I(N__61793));
    InMux I__13939 (
            .O(N__61796),
            .I(N__61789));
    LocalMux I__13938 (
            .O(N__61793),
            .I(N__61786));
    InMux I__13937 (
            .O(N__61792),
            .I(N__61783));
    LocalMux I__13936 (
            .O(N__61789),
            .I(N__61774));
    Span4Mux_v I__13935 (
            .O(N__61786),
            .I(N__61774));
    LocalMux I__13934 (
            .O(N__61783),
            .I(N__61774));
    InMux I__13933 (
            .O(N__61782),
            .I(N__61771));
    CascadeMux I__13932 (
            .O(N__61781),
            .I(N__61768));
    Span4Mux_v I__13931 (
            .O(N__61774),
            .I(N__61762));
    LocalMux I__13930 (
            .O(N__61771),
            .I(N__61762));
    InMux I__13929 (
            .O(N__61768),
            .I(N__61759));
    InMux I__13928 (
            .O(N__61767),
            .I(N__61756));
    Span4Mux_v I__13927 (
            .O(N__61762),
            .I(N__61753));
    LocalMux I__13926 (
            .O(N__61759),
            .I(\c0.data_in_frame_10_6 ));
    LocalMux I__13925 (
            .O(N__61756),
            .I(\c0.data_in_frame_10_6 ));
    Odrv4 I__13924 (
            .O(N__61753),
            .I(\c0.data_in_frame_10_6 ));
    InMux I__13923 (
            .O(N__61746),
            .I(N__61742));
    CascadeMux I__13922 (
            .O(N__61745),
            .I(N__61735));
    LocalMux I__13921 (
            .O(N__61742),
            .I(N__61732));
    InMux I__13920 (
            .O(N__61741),
            .I(N__61725));
    InMux I__13919 (
            .O(N__61740),
            .I(N__61725));
    InMux I__13918 (
            .O(N__61739),
            .I(N__61725));
    InMux I__13917 (
            .O(N__61738),
            .I(N__61720));
    InMux I__13916 (
            .O(N__61735),
            .I(N__61720));
    Span4Mux_v I__13915 (
            .O(N__61732),
            .I(N__61716));
    LocalMux I__13914 (
            .O(N__61725),
            .I(N__61711));
    LocalMux I__13913 (
            .O(N__61720),
            .I(N__61711));
    InMux I__13912 (
            .O(N__61719),
            .I(N__61708));
    Sp12to4 I__13911 (
            .O(N__61716),
            .I(N__61703));
    Span12Mux_v I__13910 (
            .O(N__61711),
            .I(N__61703));
    LocalMux I__13909 (
            .O(N__61708),
            .I(\c0.data_in_frame_10_7 ));
    Odrv12 I__13908 (
            .O(N__61703),
            .I(\c0.data_in_frame_10_7 ));
    InMux I__13907 (
            .O(N__61698),
            .I(N__61695));
    LocalMux I__13906 (
            .O(N__61695),
            .I(N__61692));
    Span4Mux_h I__13905 (
            .O(N__61692),
            .I(N__61688));
    InMux I__13904 (
            .O(N__61691),
            .I(N__61685));
    Odrv4 I__13903 (
            .O(N__61688),
            .I(\c0.n13734 ));
    LocalMux I__13902 (
            .O(N__61685),
            .I(\c0.n13734 ));
    CascadeMux I__13901 (
            .O(N__61680),
            .I(\c0.n39_adj_4708_cascade_ ));
    InMux I__13900 (
            .O(N__61677),
            .I(N__61674));
    LocalMux I__13899 (
            .O(N__61674),
            .I(N__61671));
    Span4Mux_h I__13898 (
            .O(N__61671),
            .I(N__61668));
    Span4Mux_v I__13897 (
            .O(N__61668),
            .I(N__61665));
    Odrv4 I__13896 (
            .O(N__61665),
            .I(\c0.n63 ));
    CascadeMux I__13895 (
            .O(N__61662),
            .I(\c0.n64_cascade_ ));
    CascadeMux I__13894 (
            .O(N__61659),
            .I(N__61655));
    InMux I__13893 (
            .O(N__61658),
            .I(N__61652));
    InMux I__13892 (
            .O(N__61655),
            .I(N__61649));
    LocalMux I__13891 (
            .O(N__61652),
            .I(N__61645));
    LocalMux I__13890 (
            .O(N__61649),
            .I(N__61642));
    InMux I__13889 (
            .O(N__61648),
            .I(N__61639));
    Span4Mux_h I__13888 (
            .O(N__61645),
            .I(N__61634));
    Span4Mux_h I__13887 (
            .O(N__61642),
            .I(N__61634));
    LocalMux I__13886 (
            .O(N__61639),
            .I(\c0.n13721 ));
    Odrv4 I__13885 (
            .O(N__61634),
            .I(\c0.n13721 ));
    InMux I__13884 (
            .O(N__61629),
            .I(N__61626));
    LocalMux I__13883 (
            .O(N__61626),
            .I(\c0.n55_adj_4709 ));
    CascadeMux I__13882 (
            .O(N__61623),
            .I(N__61620));
    InMux I__13881 (
            .O(N__61620),
            .I(N__61617));
    LocalMux I__13880 (
            .O(N__61617),
            .I(N__61613));
    InMux I__13879 (
            .O(N__61616),
            .I(N__61610));
    Span4Mux_v I__13878 (
            .O(N__61613),
            .I(N__61607));
    LocalMux I__13877 (
            .O(N__61610),
            .I(N__61604));
    Span4Mux_h I__13876 (
            .O(N__61607),
            .I(N__61601));
    Odrv4 I__13875 (
            .O(N__61604),
            .I(\c0.n13186 ));
    Odrv4 I__13874 (
            .O(N__61601),
            .I(\c0.n13186 ));
    CascadeMux I__13873 (
            .O(N__61596),
            .I(N__61593));
    InMux I__13872 (
            .O(N__61593),
            .I(N__61590));
    LocalMux I__13871 (
            .O(N__61590),
            .I(N__61586));
    InMux I__13870 (
            .O(N__61589),
            .I(N__61583));
    Span4Mux_v I__13869 (
            .O(N__61586),
            .I(N__61579));
    LocalMux I__13868 (
            .O(N__61583),
            .I(N__61576));
    InMux I__13867 (
            .O(N__61582),
            .I(N__61573));
    Span4Mux_h I__13866 (
            .O(N__61579),
            .I(N__61570));
    Span12Mux_h I__13865 (
            .O(N__61576),
            .I(N__61567));
    LocalMux I__13864 (
            .O(N__61573),
            .I(\c0.data_in_frame_10_5 ));
    Odrv4 I__13863 (
            .O(N__61570),
            .I(\c0.data_in_frame_10_5 ));
    Odrv12 I__13862 (
            .O(N__61567),
            .I(\c0.data_in_frame_10_5 ));
    CascadeMux I__13861 (
            .O(N__61560),
            .I(\c0.n96_cascade_ ));
    InMux I__13860 (
            .O(N__61557),
            .I(N__61554));
    LocalMux I__13859 (
            .O(N__61554),
            .I(N__61549));
    InMux I__13858 (
            .O(N__61553),
            .I(N__61545));
    InMux I__13857 (
            .O(N__61552),
            .I(N__61542));
    Span4Mux_h I__13856 (
            .O(N__61549),
            .I(N__61538));
    CascadeMux I__13855 (
            .O(N__61548),
            .I(N__61535));
    LocalMux I__13854 (
            .O(N__61545),
            .I(N__61530));
    LocalMux I__13853 (
            .O(N__61542),
            .I(N__61530));
    CascadeMux I__13852 (
            .O(N__61541),
            .I(N__61527));
    Span4Mux_h I__13851 (
            .O(N__61538),
            .I(N__61524));
    InMux I__13850 (
            .O(N__61535),
            .I(N__61521));
    Span4Mux_v I__13849 (
            .O(N__61530),
            .I(N__61518));
    InMux I__13848 (
            .O(N__61527),
            .I(N__61515));
    Span4Mux_v I__13847 (
            .O(N__61524),
            .I(N__61512));
    LocalMux I__13846 (
            .O(N__61521),
            .I(\c0.data_in_frame_8_0 ));
    Odrv4 I__13845 (
            .O(N__61518),
            .I(\c0.data_in_frame_8_0 ));
    LocalMux I__13844 (
            .O(N__61515),
            .I(\c0.data_in_frame_8_0 ));
    Odrv4 I__13843 (
            .O(N__61512),
            .I(\c0.data_in_frame_8_0 ));
    CascadeMux I__13842 (
            .O(N__61503),
            .I(N__61500));
    InMux I__13841 (
            .O(N__61500),
            .I(N__61497));
    LocalMux I__13840 (
            .O(N__61497),
            .I(N__61494));
    Span4Mux_v I__13839 (
            .O(N__61494),
            .I(N__61491));
    Odrv4 I__13838 (
            .O(N__61491),
            .I(\c0.n104 ));
    InMux I__13837 (
            .O(N__61488),
            .I(N__61482));
    InMux I__13836 (
            .O(N__61487),
            .I(N__61482));
    LocalMux I__13835 (
            .O(N__61482),
            .I(\c0.n7_adj_4253 ));
    CascadeMux I__13834 (
            .O(N__61479),
            .I(N__61476));
    InMux I__13833 (
            .O(N__61476),
            .I(N__61470));
    InMux I__13832 (
            .O(N__61475),
            .I(N__61470));
    LocalMux I__13831 (
            .O(N__61470),
            .I(\c0.n5_adj_4252 ));
    InMux I__13830 (
            .O(N__61467),
            .I(N__61463));
    InMux I__13829 (
            .O(N__61466),
            .I(N__61460));
    LocalMux I__13828 (
            .O(N__61463),
            .I(N__61457));
    LocalMux I__13827 (
            .O(N__61460),
            .I(N__61454));
    Span4Mux_h I__13826 (
            .O(N__61457),
            .I(N__61451));
    Span4Mux_v I__13825 (
            .O(N__61454),
            .I(N__61448));
    Span4Mux_h I__13824 (
            .O(N__61451),
            .I(N__61443));
    Span4Mux_h I__13823 (
            .O(N__61448),
            .I(N__61443));
    Odrv4 I__13822 (
            .O(N__61443),
            .I(\c0.n5_adj_4443 ));
    CascadeMux I__13821 (
            .O(N__61440),
            .I(\c0.n13734_cascade_ ));
    InMux I__13820 (
            .O(N__61437),
            .I(N__61434));
    LocalMux I__13819 (
            .O(N__61434),
            .I(N__61430));
    InMux I__13818 (
            .O(N__61433),
            .I(N__61426));
    Span4Mux_v I__13817 (
            .O(N__61430),
            .I(N__61421));
    InMux I__13816 (
            .O(N__61429),
            .I(N__61418));
    LocalMux I__13815 (
            .O(N__61426),
            .I(N__61415));
    InMux I__13814 (
            .O(N__61425),
            .I(N__61412));
    InMux I__13813 (
            .O(N__61424),
            .I(N__61409));
    Sp12to4 I__13812 (
            .O(N__61421),
            .I(N__61404));
    LocalMux I__13811 (
            .O(N__61418),
            .I(N__61404));
    Span4Mux_v I__13810 (
            .O(N__61415),
            .I(N__61399));
    LocalMux I__13809 (
            .O(N__61412),
            .I(N__61399));
    LocalMux I__13808 (
            .O(N__61409),
            .I(\c0.n17734 ));
    Odrv12 I__13807 (
            .O(N__61404),
            .I(\c0.n17734 ));
    Odrv4 I__13806 (
            .O(N__61399),
            .I(\c0.n17734 ));
    InMux I__13805 (
            .O(N__61392),
            .I(N__61388));
    InMux I__13804 (
            .O(N__61391),
            .I(N__61385));
    LocalMux I__13803 (
            .O(N__61388),
            .I(N__61381));
    LocalMux I__13802 (
            .O(N__61385),
            .I(N__61377));
    InMux I__13801 (
            .O(N__61384),
            .I(N__61374));
    Span4Mux_v I__13800 (
            .O(N__61381),
            .I(N__61371));
    InMux I__13799 (
            .O(N__61380),
            .I(N__61368));
    Span4Mux_v I__13798 (
            .O(N__61377),
            .I(N__61363));
    LocalMux I__13797 (
            .O(N__61374),
            .I(N__61363));
    Sp12to4 I__13796 (
            .O(N__61371),
            .I(N__61360));
    LocalMux I__13795 (
            .O(N__61368),
            .I(N__61357));
    Sp12to4 I__13794 (
            .O(N__61363),
            .I(N__61352));
    Span12Mux_h I__13793 (
            .O(N__61360),
            .I(N__61352));
    Odrv4 I__13792 (
            .O(N__61357),
            .I(\c0.n12973 ));
    Odrv12 I__13791 (
            .O(N__61352),
            .I(\c0.n12973 ));
    CascadeMux I__13790 (
            .O(N__61347),
            .I(\c0.n30_adj_4705_cascade_ ));
    CascadeMux I__13789 (
            .O(N__61344),
            .I(\c0.n23523_cascade_ ));
    InMux I__13788 (
            .O(N__61341),
            .I(N__61338));
    LocalMux I__13787 (
            .O(N__61338),
            .I(\c0.n30 ));
    InMux I__13786 (
            .O(N__61335),
            .I(N__61330));
    InMux I__13785 (
            .O(N__61334),
            .I(N__61327));
    InMux I__13784 (
            .O(N__61333),
            .I(N__61324));
    LocalMux I__13783 (
            .O(N__61330),
            .I(N__61321));
    LocalMux I__13782 (
            .O(N__61327),
            .I(N__61316));
    LocalMux I__13781 (
            .O(N__61324),
            .I(N__61316));
    Span12Mux_h I__13780 (
            .O(N__61321),
            .I(N__61313));
    Span12Mux_h I__13779 (
            .O(N__61316),
            .I(N__61310));
    Odrv12 I__13778 (
            .O(N__61313),
            .I(\c0.n13075 ));
    Odrv12 I__13777 (
            .O(N__61310),
            .I(\c0.n13075 ));
    CascadeMux I__13776 (
            .O(N__61305),
            .I(\c0.n7_adj_4634_cascade_ ));
    InMux I__13775 (
            .O(N__61302),
            .I(N__61299));
    LocalMux I__13774 (
            .O(N__61299),
            .I(N__61295));
    CascadeMux I__13773 (
            .O(N__61298),
            .I(N__61289));
    Span4Mux_h I__13772 (
            .O(N__61295),
            .I(N__61285));
    InMux I__13771 (
            .O(N__61294),
            .I(N__61282));
    InMux I__13770 (
            .O(N__61293),
            .I(N__61277));
    InMux I__13769 (
            .O(N__61292),
            .I(N__61277));
    InMux I__13768 (
            .O(N__61289),
            .I(N__61272));
    InMux I__13767 (
            .O(N__61288),
            .I(N__61272));
    Odrv4 I__13766 (
            .O(N__61285),
            .I(\c0.n22230 ));
    LocalMux I__13765 (
            .O(N__61282),
            .I(\c0.n22230 ));
    LocalMux I__13764 (
            .O(N__61277),
            .I(\c0.n22230 ));
    LocalMux I__13763 (
            .O(N__61272),
            .I(\c0.n22230 ));
    InMux I__13762 (
            .O(N__61263),
            .I(N__61259));
    InMux I__13761 (
            .O(N__61262),
            .I(N__61256));
    LocalMux I__13760 (
            .O(N__61259),
            .I(N__61252));
    LocalMux I__13759 (
            .O(N__61256),
            .I(N__61249));
    InMux I__13758 (
            .O(N__61255),
            .I(N__61246));
    Span4Mux_v I__13757 (
            .O(N__61252),
            .I(N__61242));
    Span4Mux_v I__13756 (
            .O(N__61249),
            .I(N__61239));
    LocalMux I__13755 (
            .O(N__61246),
            .I(N__61236));
    InMux I__13754 (
            .O(N__61245),
            .I(N__61232));
    Span4Mux_v I__13753 (
            .O(N__61242),
            .I(N__61227));
    Span4Mux_v I__13752 (
            .O(N__61239),
            .I(N__61227));
    Span4Mux_h I__13751 (
            .O(N__61236),
            .I(N__61224));
    InMux I__13750 (
            .O(N__61235),
            .I(N__61221));
    LocalMux I__13749 (
            .O(N__61232),
            .I(\c0.data_in_frame_9_4 ));
    Odrv4 I__13748 (
            .O(N__61227),
            .I(\c0.data_in_frame_9_4 ));
    Odrv4 I__13747 (
            .O(N__61224),
            .I(\c0.data_in_frame_9_4 ));
    LocalMux I__13746 (
            .O(N__61221),
            .I(\c0.data_in_frame_9_4 ));
    CascadeMux I__13745 (
            .O(N__61212),
            .I(N__61209));
    InMux I__13744 (
            .O(N__61209),
            .I(N__61206));
    LocalMux I__13743 (
            .O(N__61206),
            .I(N__61203));
    Span4Mux_h I__13742 (
            .O(N__61203),
            .I(N__61200));
    Span4Mux_v I__13741 (
            .O(N__61200),
            .I(N__61197));
    Odrv4 I__13740 (
            .O(N__61197),
            .I(\c0.n150 ));
    InMux I__13739 (
            .O(N__61194),
            .I(N__61191));
    LocalMux I__13738 (
            .O(N__61191),
            .I(N__61188));
    Span4Mux_v I__13737 (
            .O(N__61188),
            .I(N__61185));
    Span4Mux_h I__13736 (
            .O(N__61185),
            .I(N__61182));
    Span4Mux_h I__13735 (
            .O(N__61182),
            .I(N__61179));
    Odrv4 I__13734 (
            .O(N__61179),
            .I(\c0.n13651 ));
    CascadeMux I__13733 (
            .O(N__61176),
            .I(N__61172));
    InMux I__13732 (
            .O(N__61175),
            .I(N__61169));
    InMux I__13731 (
            .O(N__61172),
            .I(N__61166));
    LocalMux I__13730 (
            .O(N__61169),
            .I(N__61163));
    LocalMux I__13729 (
            .O(N__61166),
            .I(N__61160));
    Span4Mux_v I__13728 (
            .O(N__61163),
            .I(N__61157));
    Odrv4 I__13727 (
            .O(N__61160),
            .I(\c0.n18_adj_4228 ));
    Odrv4 I__13726 (
            .O(N__61157),
            .I(\c0.n18_adj_4228 ));
    CascadeMux I__13725 (
            .O(N__61152),
            .I(\c0.n27_cascade_ ));
    InMux I__13724 (
            .O(N__61149),
            .I(N__61146));
    LocalMux I__13723 (
            .O(N__61146),
            .I(N__61143));
    Span4Mux_h I__13722 (
            .O(N__61143),
            .I(N__61139));
    InMux I__13721 (
            .O(N__61142),
            .I(N__61136));
    Span4Mux_h I__13720 (
            .O(N__61139),
            .I(N__61133));
    LocalMux I__13719 (
            .O(N__61136),
            .I(\c0.n19 ));
    Odrv4 I__13718 (
            .O(N__61133),
            .I(\c0.n19 ));
    CascadeMux I__13717 (
            .O(N__61128),
            .I(\c0.n23528_cascade_ ));
    CascadeMux I__13716 (
            .O(N__61125),
            .I(\c0.n34_adj_4278_cascade_ ));
    InMux I__13715 (
            .O(N__61122),
            .I(N__61119));
    LocalMux I__13714 (
            .O(N__61119),
            .I(N__61116));
    Odrv4 I__13713 (
            .O(N__61116),
            .I(\c0.n36 ));
    InMux I__13712 (
            .O(N__61113),
            .I(N__61104));
    InMux I__13711 (
            .O(N__61112),
            .I(N__61104));
    InMux I__13710 (
            .O(N__61111),
            .I(N__61104));
    LocalMux I__13709 (
            .O(N__61104),
            .I(\c0.n48_adj_4227 ));
    InMux I__13708 (
            .O(N__61101),
            .I(N__61098));
    LocalMux I__13707 (
            .O(N__61098),
            .I(N__61095));
    Span4Mux_v I__13706 (
            .O(N__61095),
            .I(N__61091));
    InMux I__13705 (
            .O(N__61094),
            .I(N__61088));
    Odrv4 I__13704 (
            .O(N__61091),
            .I(\c0.n18_adj_4314 ));
    LocalMux I__13703 (
            .O(N__61088),
            .I(\c0.n18_adj_4314 ));
    CascadeMux I__13702 (
            .O(N__61083),
            .I(N__61080));
    InMux I__13701 (
            .O(N__61080),
            .I(N__61077));
    LocalMux I__13700 (
            .O(N__61077),
            .I(N__61074));
    Span4Mux_h I__13699 (
            .O(N__61074),
            .I(N__61071));
    Odrv4 I__13698 (
            .O(N__61071),
            .I(\c0.n24_adj_4724 ));
    InMux I__13697 (
            .O(N__61068),
            .I(N__61065));
    LocalMux I__13696 (
            .O(N__61065),
            .I(N__61061));
    CascadeMux I__13695 (
            .O(N__61064),
            .I(N__61058));
    Span4Mux_v I__13694 (
            .O(N__61061),
            .I(N__61054));
    InMux I__13693 (
            .O(N__61058),
            .I(N__61051));
    InMux I__13692 (
            .O(N__61057),
            .I(N__61048));
    Span4Mux_v I__13691 (
            .O(N__61054),
            .I(N__61045));
    LocalMux I__13690 (
            .O(N__61051),
            .I(N__61040));
    LocalMux I__13689 (
            .O(N__61048),
            .I(N__61037));
    Span4Mux_v I__13688 (
            .O(N__61045),
            .I(N__61032));
    InMux I__13687 (
            .O(N__61044),
            .I(N__61025));
    InMux I__13686 (
            .O(N__61043),
            .I(N__61025));
    Span4Mux_v I__13685 (
            .O(N__61040),
            .I(N__61020));
    Span4Mux_v I__13684 (
            .O(N__61037),
            .I(N__61020));
    InMux I__13683 (
            .O(N__61036),
            .I(N__61017));
    InMux I__13682 (
            .O(N__61035),
            .I(N__61014));
    Span4Mux_h I__13681 (
            .O(N__61032),
            .I(N__61011));
    InMux I__13680 (
            .O(N__61031),
            .I(N__61008));
    InMux I__13679 (
            .O(N__61030),
            .I(N__61005));
    LocalMux I__13678 (
            .O(N__61025),
            .I(N__60998));
    Sp12to4 I__13677 (
            .O(N__61020),
            .I(N__60998));
    LocalMux I__13676 (
            .O(N__61017),
            .I(N__60998));
    LocalMux I__13675 (
            .O(N__61014),
            .I(data_in_frame_1_0));
    Odrv4 I__13674 (
            .O(N__61011),
            .I(data_in_frame_1_0));
    LocalMux I__13673 (
            .O(N__61008),
            .I(data_in_frame_1_0));
    LocalMux I__13672 (
            .O(N__61005),
            .I(data_in_frame_1_0));
    Odrv12 I__13671 (
            .O(N__60998),
            .I(data_in_frame_1_0));
    InMux I__13670 (
            .O(N__60987),
            .I(N__60984));
    LocalMux I__13669 (
            .O(N__60984),
            .I(\c0.n5_adj_4711 ));
    InMux I__13668 (
            .O(N__60981),
            .I(N__60978));
    LocalMux I__13667 (
            .O(N__60978),
            .I(N__60975));
    Span4Mux_v I__13666 (
            .O(N__60975),
            .I(N__60972));
    Odrv4 I__13665 (
            .O(N__60972),
            .I(\c0.n16_adj_4716 ));
    CascadeMux I__13664 (
            .O(N__60969),
            .I(\c0.n28_adj_4718_cascade_ ));
    InMux I__13663 (
            .O(N__60966),
            .I(N__60963));
    LocalMux I__13662 (
            .O(N__60963),
            .I(N__60960));
    Odrv4 I__13661 (
            .O(N__60960),
            .I(\c0.n24_adj_4717 ));
    InMux I__13660 (
            .O(N__60957),
            .I(N__60954));
    LocalMux I__13659 (
            .O(N__60954),
            .I(N__60949));
    CascadeMux I__13658 (
            .O(N__60953),
            .I(N__60946));
    CascadeMux I__13657 (
            .O(N__60952),
            .I(N__60943));
    Span4Mux_h I__13656 (
            .O(N__60949),
            .I(N__60939));
    InMux I__13655 (
            .O(N__60946),
            .I(N__60934));
    InMux I__13654 (
            .O(N__60943),
            .I(N__60934));
    InMux I__13653 (
            .O(N__60942),
            .I(N__60931));
    Odrv4 I__13652 (
            .O(N__60939),
            .I(\c0.n23_adj_4599 ));
    LocalMux I__13651 (
            .O(N__60934),
            .I(\c0.n23_adj_4599 ));
    LocalMux I__13650 (
            .O(N__60931),
            .I(\c0.n23_adj_4599 ));
    InMux I__13649 (
            .O(N__60924),
            .I(N__60921));
    LocalMux I__13648 (
            .O(N__60921),
            .I(N__60918));
    Odrv4 I__13647 (
            .O(N__60918),
            .I(\c0.n4_adj_4446 ));
    CascadeMux I__13646 (
            .O(N__60915),
            .I(\c0.n4_adj_4446_cascade_ ));
    InMux I__13645 (
            .O(N__60912),
            .I(N__60909));
    LocalMux I__13644 (
            .O(N__60909),
            .I(\c0.n26_adj_4714 ));
    InMux I__13643 (
            .O(N__60906),
            .I(N__60900));
    InMux I__13642 (
            .O(N__60905),
            .I(N__60900));
    LocalMux I__13641 (
            .O(N__60900),
            .I(N__60896));
    CascadeMux I__13640 (
            .O(N__60899),
            .I(N__60892));
    Span4Mux_v I__13639 (
            .O(N__60896),
            .I(N__60888));
    CascadeMux I__13638 (
            .O(N__60895),
            .I(N__60885));
    InMux I__13637 (
            .O(N__60892),
            .I(N__60877));
    InMux I__13636 (
            .O(N__60891),
            .I(N__60877));
    Span4Mux_h I__13635 (
            .O(N__60888),
            .I(N__60874));
    InMux I__13634 (
            .O(N__60885),
            .I(N__60867));
    InMux I__13633 (
            .O(N__60884),
            .I(N__60867));
    InMux I__13632 (
            .O(N__60883),
            .I(N__60867));
    InMux I__13631 (
            .O(N__60882),
            .I(N__60864));
    LocalMux I__13630 (
            .O(N__60877),
            .I(\c0.data_in_frame_4_0 ));
    Odrv4 I__13629 (
            .O(N__60874),
            .I(\c0.data_in_frame_4_0 ));
    LocalMux I__13628 (
            .O(N__60867),
            .I(\c0.data_in_frame_4_0 ));
    LocalMux I__13627 (
            .O(N__60864),
            .I(\c0.data_in_frame_4_0 ));
    InMux I__13626 (
            .O(N__60855),
            .I(N__60851));
    InMux I__13625 (
            .O(N__60854),
            .I(N__60847));
    LocalMux I__13624 (
            .O(N__60851),
            .I(N__60844));
    InMux I__13623 (
            .O(N__60850),
            .I(N__60841));
    LocalMux I__13622 (
            .O(N__60847),
            .I(N__60836));
    Span4Mux_v I__13621 (
            .O(N__60844),
            .I(N__60836));
    LocalMux I__13620 (
            .O(N__60841),
            .I(N__60829));
    Span4Mux_h I__13619 (
            .O(N__60836),
            .I(N__60829));
    InMux I__13618 (
            .O(N__60835),
            .I(N__60824));
    InMux I__13617 (
            .O(N__60834),
            .I(N__60824));
    Odrv4 I__13616 (
            .O(N__60829),
            .I(\c0.data_in_frame_3_6 ));
    LocalMux I__13615 (
            .O(N__60824),
            .I(\c0.data_in_frame_3_6 ));
    InMux I__13614 (
            .O(N__60819),
            .I(N__60814));
    InMux I__13613 (
            .O(N__60818),
            .I(N__60809));
    InMux I__13612 (
            .O(N__60817),
            .I(N__60809));
    LocalMux I__13611 (
            .O(N__60814),
            .I(N__60806));
    LocalMux I__13610 (
            .O(N__60809),
            .I(N__60803));
    Odrv4 I__13609 (
            .O(N__60806),
            .I(\c0.n23597 ));
    Odrv4 I__13608 (
            .O(N__60803),
            .I(\c0.n23597 ));
    CascadeMux I__13607 (
            .O(N__60798),
            .I(N__60793));
    CascadeMux I__13606 (
            .O(N__60797),
            .I(N__60789));
    CascadeMux I__13605 (
            .O(N__60796),
            .I(N__60786));
    InMux I__13604 (
            .O(N__60793),
            .I(N__60783));
    InMux I__13603 (
            .O(N__60792),
            .I(N__60780));
    InMux I__13602 (
            .O(N__60789),
            .I(N__60775));
    InMux I__13601 (
            .O(N__60786),
            .I(N__60775));
    LocalMux I__13600 (
            .O(N__60783),
            .I(N__60770));
    LocalMux I__13599 (
            .O(N__60780),
            .I(N__60765));
    LocalMux I__13598 (
            .O(N__60775),
            .I(N__60765));
    InMux I__13597 (
            .O(N__60774),
            .I(N__60760));
    InMux I__13596 (
            .O(N__60773),
            .I(N__60760));
    Odrv12 I__13595 (
            .O(N__60770),
            .I(\c0.data_in_frame_2_0 ));
    Odrv4 I__13594 (
            .O(N__60765),
            .I(\c0.data_in_frame_2_0 ));
    LocalMux I__13593 (
            .O(N__60760),
            .I(\c0.data_in_frame_2_0 ));
    CascadeMux I__13592 (
            .O(N__60753),
            .I(\c0.n37_cascade_ ));
    CascadeMux I__13591 (
            .O(N__60750),
            .I(\c0.n22647_cascade_ ));
    CascadeMux I__13590 (
            .O(N__60747),
            .I(N__60743));
    CascadeMux I__13589 (
            .O(N__60746),
            .I(N__60738));
    InMux I__13588 (
            .O(N__60743),
            .I(N__60734));
    InMux I__13587 (
            .O(N__60742),
            .I(N__60731));
    InMux I__13586 (
            .O(N__60741),
            .I(N__60728));
    InMux I__13585 (
            .O(N__60738),
            .I(N__60723));
    InMux I__13584 (
            .O(N__60737),
            .I(N__60723));
    LocalMux I__13583 (
            .O(N__60734),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__13582 (
            .O(N__60731),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__13581 (
            .O(N__60728),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__13580 (
            .O(N__60723),
            .I(\c0.data_in_frame_2_6 ));
    InMux I__13579 (
            .O(N__60714),
            .I(N__60711));
    LocalMux I__13578 (
            .O(N__60711),
            .I(N__60708));
    Span4Mux_h I__13577 (
            .O(N__60708),
            .I(N__60705));
    Span4Mux_h I__13576 (
            .O(N__60705),
            .I(N__60702));
    Odrv4 I__13575 (
            .O(N__60702),
            .I(\c0.n24747 ));
    InMux I__13574 (
            .O(N__60699),
            .I(N__60696));
    LocalMux I__13573 (
            .O(N__60696),
            .I(\c0.n10_adj_4722 ));
    CascadeMux I__13572 (
            .O(N__60693),
            .I(\c0.n14_adj_4616_cascade_ ));
    InMux I__13571 (
            .O(N__60690),
            .I(N__60687));
    LocalMux I__13570 (
            .O(N__60687),
            .I(N__60683));
    InMux I__13569 (
            .O(N__60686),
            .I(N__60680));
    Span4Mux_v I__13568 (
            .O(N__60683),
            .I(N__60677));
    LocalMux I__13567 (
            .O(N__60680),
            .I(N__60674));
    Span4Mux_h I__13566 (
            .O(N__60677),
            .I(N__60671));
    Odrv4 I__13565 (
            .O(N__60674),
            .I(\c0.n23666 ));
    Odrv4 I__13564 (
            .O(N__60671),
            .I(\c0.n23666 ));
    CascadeMux I__13563 (
            .O(N__60666),
            .I(N__60663));
    InMux I__13562 (
            .O(N__60663),
            .I(N__60660));
    LocalMux I__13561 (
            .O(N__60660),
            .I(N__60657));
    Odrv4 I__13560 (
            .O(N__60657),
            .I(\c0.n37 ));
    InMux I__13559 (
            .O(N__60654),
            .I(N__60651));
    LocalMux I__13558 (
            .O(N__60651),
            .I(\c0.n55 ));
    CascadeMux I__13557 (
            .O(N__60648),
            .I(N__60645));
    InMux I__13556 (
            .O(N__60645),
            .I(N__60641));
    InMux I__13555 (
            .O(N__60644),
            .I(N__60638));
    LocalMux I__13554 (
            .O(N__60641),
            .I(N__60628));
    LocalMux I__13553 (
            .O(N__60638),
            .I(N__60625));
    InMux I__13552 (
            .O(N__60637),
            .I(N__60620));
    InMux I__13551 (
            .O(N__60636),
            .I(N__60620));
    InMux I__13550 (
            .O(N__60635),
            .I(N__60617));
    InMux I__13549 (
            .O(N__60634),
            .I(N__60610));
    InMux I__13548 (
            .O(N__60633),
            .I(N__60610));
    InMux I__13547 (
            .O(N__60632),
            .I(N__60610));
    InMux I__13546 (
            .O(N__60631),
            .I(N__60607));
    Odrv4 I__13545 (
            .O(N__60628),
            .I(\c0.data_in_frame_0_6 ));
    Odrv4 I__13544 (
            .O(N__60625),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__13543 (
            .O(N__60620),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__13542 (
            .O(N__60617),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__13541 (
            .O(N__60610),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__13540 (
            .O(N__60607),
            .I(\c0.data_in_frame_0_6 ));
    InMux I__13539 (
            .O(N__60594),
            .I(N__60591));
    LocalMux I__13538 (
            .O(N__60591),
            .I(\c0.n24016 ));
    InMux I__13537 (
            .O(N__60588),
            .I(N__60585));
    LocalMux I__13536 (
            .O(N__60585),
            .I(N__60582));
    Span4Mux_h I__13535 (
            .O(N__60582),
            .I(N__60579));
    Span4Mux_h I__13534 (
            .O(N__60579),
            .I(N__60576));
    Odrv4 I__13533 (
            .O(N__60576),
            .I(\c0.n24749 ));
    InMux I__13532 (
            .O(N__60573),
            .I(N__60570));
    LocalMux I__13531 (
            .O(N__60570),
            .I(N__60567));
    Span4Mux_v I__13530 (
            .O(N__60567),
            .I(N__60563));
    InMux I__13529 (
            .O(N__60566),
            .I(N__60559));
    Span4Mux_h I__13528 (
            .O(N__60563),
            .I(N__60554));
    CascadeMux I__13527 (
            .O(N__60562),
            .I(N__60549));
    LocalMux I__13526 (
            .O(N__60559),
            .I(N__60542));
    InMux I__13525 (
            .O(N__60558),
            .I(N__60537));
    InMux I__13524 (
            .O(N__60557),
            .I(N__60537));
    Sp12to4 I__13523 (
            .O(N__60554),
            .I(N__60530));
    InMux I__13522 (
            .O(N__60553),
            .I(N__60527));
    InMux I__13521 (
            .O(N__60552),
            .I(N__60524));
    InMux I__13520 (
            .O(N__60549),
            .I(N__60521));
    InMux I__13519 (
            .O(N__60548),
            .I(N__60518));
    InMux I__13518 (
            .O(N__60547),
            .I(N__60515));
    CascadeMux I__13517 (
            .O(N__60546),
            .I(N__60512));
    CascadeMux I__13516 (
            .O(N__60545),
            .I(N__60508));
    Span4Mux_v I__13515 (
            .O(N__60542),
            .I(N__60504));
    LocalMux I__13514 (
            .O(N__60537),
            .I(N__60501));
    InMux I__13513 (
            .O(N__60536),
            .I(N__60494));
    InMux I__13512 (
            .O(N__60535),
            .I(N__60494));
    InMux I__13511 (
            .O(N__60534),
            .I(N__60494));
    CascadeMux I__13510 (
            .O(N__60533),
            .I(N__60491));
    Span12Mux_h I__13509 (
            .O(N__60530),
            .I(N__60481));
    LocalMux I__13508 (
            .O(N__60527),
            .I(N__60481));
    LocalMux I__13507 (
            .O(N__60524),
            .I(N__60481));
    LocalMux I__13506 (
            .O(N__60521),
            .I(N__60481));
    LocalMux I__13505 (
            .O(N__60518),
            .I(N__60478));
    LocalMux I__13504 (
            .O(N__60515),
            .I(N__60475));
    InMux I__13503 (
            .O(N__60512),
            .I(N__60470));
    InMux I__13502 (
            .O(N__60511),
            .I(N__60470));
    InMux I__13501 (
            .O(N__60508),
            .I(N__60465));
    InMux I__13500 (
            .O(N__60507),
            .I(N__60465));
    Span4Mux_h I__13499 (
            .O(N__60504),
            .I(N__60458));
    Span4Mux_h I__13498 (
            .O(N__60501),
            .I(N__60458));
    LocalMux I__13497 (
            .O(N__60494),
            .I(N__60458));
    InMux I__13496 (
            .O(N__60491),
            .I(N__60453));
    InMux I__13495 (
            .O(N__60490),
            .I(N__60453));
    Odrv12 I__13494 (
            .O(N__60481),
            .I(data_in_frame_1_4));
    Odrv4 I__13493 (
            .O(N__60478),
            .I(data_in_frame_1_4));
    Odrv4 I__13492 (
            .O(N__60475),
            .I(data_in_frame_1_4));
    LocalMux I__13491 (
            .O(N__60470),
            .I(data_in_frame_1_4));
    LocalMux I__13490 (
            .O(N__60465),
            .I(data_in_frame_1_4));
    Odrv4 I__13489 (
            .O(N__60458),
            .I(data_in_frame_1_4));
    LocalMux I__13488 (
            .O(N__60453),
            .I(data_in_frame_1_4));
    InMux I__13487 (
            .O(N__60438),
            .I(N__60435));
    LocalMux I__13486 (
            .O(N__60435),
            .I(N__60432));
    Span4Mux_v I__13485 (
            .O(N__60432),
            .I(N__60428));
    InMux I__13484 (
            .O(N__60431),
            .I(N__60424));
    Span4Mux_h I__13483 (
            .O(N__60428),
            .I(N__60421));
    CascadeMux I__13482 (
            .O(N__60427),
            .I(N__60418));
    LocalMux I__13481 (
            .O(N__60424),
            .I(N__60410));
    Span4Mux_v I__13480 (
            .O(N__60421),
            .I(N__60405));
    InMux I__13479 (
            .O(N__60418),
            .I(N__60394));
    InMux I__13478 (
            .O(N__60417),
            .I(N__60394));
    InMux I__13477 (
            .O(N__60416),
            .I(N__60394));
    InMux I__13476 (
            .O(N__60415),
            .I(N__60394));
    InMux I__13475 (
            .O(N__60414),
            .I(N__60394));
    InMux I__13474 (
            .O(N__60413),
            .I(N__60391));
    Span4Mux_h I__13473 (
            .O(N__60410),
            .I(N__60388));
    CascadeMux I__13472 (
            .O(N__60409),
            .I(N__60382));
    CascadeMux I__13471 (
            .O(N__60408),
            .I(N__60379));
    Span4Mux_v I__13470 (
            .O(N__60405),
            .I(N__60372));
    LocalMux I__13469 (
            .O(N__60394),
            .I(N__60372));
    LocalMux I__13468 (
            .O(N__60391),
            .I(N__60369));
    Span4Mux_h I__13467 (
            .O(N__60388),
            .I(N__60366));
    InMux I__13466 (
            .O(N__60387),
            .I(N__60363));
    InMux I__13465 (
            .O(N__60386),
            .I(N__60360));
    InMux I__13464 (
            .O(N__60385),
            .I(N__60357));
    InMux I__13463 (
            .O(N__60382),
            .I(N__60354));
    InMux I__13462 (
            .O(N__60379),
            .I(N__60347));
    InMux I__13461 (
            .O(N__60378),
            .I(N__60347));
    InMux I__13460 (
            .O(N__60377),
            .I(N__60347));
    Span4Mux_v I__13459 (
            .O(N__60372),
            .I(N__60342));
    Span4Mux_v I__13458 (
            .O(N__60369),
            .I(N__60342));
    Odrv4 I__13457 (
            .O(N__60366),
            .I(data_in_frame_1_5));
    LocalMux I__13456 (
            .O(N__60363),
            .I(data_in_frame_1_5));
    LocalMux I__13455 (
            .O(N__60360),
            .I(data_in_frame_1_5));
    LocalMux I__13454 (
            .O(N__60357),
            .I(data_in_frame_1_5));
    LocalMux I__13453 (
            .O(N__60354),
            .I(data_in_frame_1_5));
    LocalMux I__13452 (
            .O(N__60347),
            .I(data_in_frame_1_5));
    Odrv4 I__13451 (
            .O(N__60342),
            .I(data_in_frame_1_5));
    InMux I__13450 (
            .O(N__60327),
            .I(N__60324));
    LocalMux I__13449 (
            .O(N__60324),
            .I(N__60321));
    Span4Mux_h I__13448 (
            .O(N__60321),
            .I(N__60318));
    Span4Mux_h I__13447 (
            .O(N__60318),
            .I(N__60315));
    Odrv4 I__13446 (
            .O(N__60315),
            .I(\c0.n37_adj_4738 ));
    CascadeMux I__13445 (
            .O(N__60312),
            .I(N__60309));
    InMux I__13444 (
            .O(N__60309),
            .I(N__60306));
    LocalMux I__13443 (
            .O(N__60306),
            .I(N__60298));
    InMux I__13442 (
            .O(N__60305),
            .I(N__60292));
    InMux I__13441 (
            .O(N__60304),
            .I(N__60289));
    InMux I__13440 (
            .O(N__60303),
            .I(N__60284));
    InMux I__13439 (
            .O(N__60302),
            .I(N__60284));
    InMux I__13438 (
            .O(N__60301),
            .I(N__60280));
    Span4Mux_v I__13437 (
            .O(N__60298),
            .I(N__60277));
    InMux I__13436 (
            .O(N__60297),
            .I(N__60274));
    InMux I__13435 (
            .O(N__60296),
            .I(N__60269));
    InMux I__13434 (
            .O(N__60295),
            .I(N__60269));
    LocalMux I__13433 (
            .O(N__60292),
            .I(N__60266));
    LocalMux I__13432 (
            .O(N__60289),
            .I(N__60261));
    LocalMux I__13431 (
            .O(N__60284),
            .I(N__60261));
    InMux I__13430 (
            .O(N__60283),
            .I(N__60258));
    LocalMux I__13429 (
            .O(N__60280),
            .I(\c0.data_in_frame_0_5 ));
    Odrv4 I__13428 (
            .O(N__60277),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__13427 (
            .O(N__60274),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__13426 (
            .O(N__60269),
            .I(\c0.data_in_frame_0_5 ));
    Odrv12 I__13425 (
            .O(N__60266),
            .I(\c0.data_in_frame_0_5 ));
    Odrv4 I__13424 (
            .O(N__60261),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__13423 (
            .O(N__60258),
            .I(\c0.data_in_frame_0_5 ));
    CascadeMux I__13422 (
            .O(N__60243),
            .I(N__60240));
    InMux I__13421 (
            .O(N__60240),
            .I(N__60236));
    CascadeMux I__13420 (
            .O(N__60239),
            .I(N__60231));
    LocalMux I__13419 (
            .O(N__60236),
            .I(N__60224));
    InMux I__13418 (
            .O(N__60235),
            .I(N__60219));
    InMux I__13417 (
            .O(N__60234),
            .I(N__60219));
    InMux I__13416 (
            .O(N__60231),
            .I(N__60212));
    InMux I__13415 (
            .O(N__60230),
            .I(N__60212));
    InMux I__13414 (
            .O(N__60229),
            .I(N__60212));
    CascadeMux I__13413 (
            .O(N__60228),
            .I(N__60209));
    CascadeMux I__13412 (
            .O(N__60227),
            .I(N__60205));
    Span4Mux_v I__13411 (
            .O(N__60224),
            .I(N__60198));
    LocalMux I__13410 (
            .O(N__60219),
            .I(N__60198));
    LocalMux I__13409 (
            .O(N__60212),
            .I(N__60195));
    InMux I__13408 (
            .O(N__60209),
            .I(N__60188));
    InMux I__13407 (
            .O(N__60208),
            .I(N__60188));
    InMux I__13406 (
            .O(N__60205),
            .I(N__60188));
    InMux I__13405 (
            .O(N__60204),
            .I(N__60183));
    InMux I__13404 (
            .O(N__60203),
            .I(N__60180));
    Span4Mux_v I__13403 (
            .O(N__60198),
            .I(N__60173));
    Span4Mux_h I__13402 (
            .O(N__60195),
            .I(N__60173));
    LocalMux I__13401 (
            .O(N__60188),
            .I(N__60173));
    InMux I__13400 (
            .O(N__60187),
            .I(N__60168));
    InMux I__13399 (
            .O(N__60186),
            .I(N__60168));
    LocalMux I__13398 (
            .O(N__60183),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__13397 (
            .O(N__60180),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__13396 (
            .O(N__60173),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__13395 (
            .O(N__60168),
            .I(\c0.data_in_frame_0_7 ));
    InMux I__13394 (
            .O(N__60159),
            .I(N__60156));
    LocalMux I__13393 (
            .O(N__60156),
            .I(N__60152));
    InMux I__13392 (
            .O(N__60155),
            .I(N__60149));
    Span4Mux_v I__13391 (
            .O(N__60152),
            .I(N__60143));
    LocalMux I__13390 (
            .O(N__60149),
            .I(N__60143));
    InMux I__13389 (
            .O(N__60148),
            .I(N__60140));
    Odrv4 I__13388 (
            .O(N__60143),
            .I(\c0.n22316 ));
    LocalMux I__13387 (
            .O(N__60140),
            .I(\c0.n22316 ));
    InMux I__13386 (
            .O(N__60135),
            .I(N__60132));
    LocalMux I__13385 (
            .O(N__60132),
            .I(N__60128));
    InMux I__13384 (
            .O(N__60131),
            .I(N__60125));
    Odrv4 I__13383 (
            .O(N__60128),
            .I(\c0.n23554 ));
    LocalMux I__13382 (
            .O(N__60125),
            .I(\c0.n23554 ));
    CascadeMux I__13381 (
            .O(N__60120),
            .I(\c0.n34_cascade_ ));
    InMux I__13380 (
            .O(N__60117),
            .I(N__60113));
    InMux I__13379 (
            .O(N__60116),
            .I(N__60110));
    LocalMux I__13378 (
            .O(N__60113),
            .I(N__60107));
    LocalMux I__13377 (
            .O(N__60110),
            .I(N__60102));
    Span4Mux_h I__13376 (
            .O(N__60107),
            .I(N__60102));
    Odrv4 I__13375 (
            .O(N__60102),
            .I(\c0.n23655 ));
    InMux I__13374 (
            .O(N__60099),
            .I(N__60096));
    LocalMux I__13373 (
            .O(N__60096),
            .I(N__60093));
    Span4Mux_h I__13372 (
            .O(N__60093),
            .I(N__60090));
    Odrv4 I__13371 (
            .O(N__60090),
            .I(\c0.n53 ));
    CascadeMux I__13370 (
            .O(N__60087),
            .I(\c0.n54_cascade_ ));
    InMux I__13369 (
            .O(N__60084),
            .I(N__60081));
    LocalMux I__13368 (
            .O(N__60081),
            .I(N__60077));
    InMux I__13367 (
            .O(N__60080),
            .I(N__60074));
    Span4Mux_h I__13366 (
            .O(N__60077),
            .I(N__60071));
    LocalMux I__13365 (
            .O(N__60074),
            .I(N__60068));
    Odrv4 I__13364 (
            .O(N__60071),
            .I(\c0.n56 ));
    Odrv4 I__13363 (
            .O(N__60068),
            .I(\c0.n56 ));
    InMux I__13362 (
            .O(N__60063),
            .I(N__60057));
    InMux I__13361 (
            .O(N__60062),
            .I(N__60054));
    InMux I__13360 (
            .O(N__60061),
            .I(N__60049));
    InMux I__13359 (
            .O(N__60060),
            .I(N__60049));
    LocalMux I__13358 (
            .O(N__60057),
            .I(N__60045));
    LocalMux I__13357 (
            .O(N__60054),
            .I(N__60040));
    LocalMux I__13356 (
            .O(N__60049),
            .I(N__60040));
    InMux I__13355 (
            .O(N__60048),
            .I(N__60037));
    Span4Mux_h I__13354 (
            .O(N__60045),
            .I(N__60030));
    Span4Mux_v I__13353 (
            .O(N__60040),
            .I(N__60030));
    LocalMux I__13352 (
            .O(N__60037),
            .I(N__60030));
    Span4Mux_v I__13351 (
            .O(N__60030),
            .I(N__60026));
    InMux I__13350 (
            .O(N__60029),
            .I(N__60023));
    Span4Mux_v I__13349 (
            .O(N__60026),
            .I(N__60020));
    LocalMux I__13348 (
            .O(N__60023),
            .I(N__60017));
    Odrv4 I__13347 (
            .O(N__60020),
            .I(\c0.n13821 ));
    Odrv4 I__13346 (
            .O(N__60017),
            .I(\c0.n13821 ));
    InMux I__13345 (
            .O(N__60012),
            .I(N__60009));
    LocalMux I__13344 (
            .O(N__60009),
            .I(N__60006));
    Odrv4 I__13343 (
            .O(N__60006),
            .I(\c0.n48 ));
    CascadeMux I__13342 (
            .O(N__60003),
            .I(\c0.n24441_cascade_ ));
    InMux I__13341 (
            .O(N__60000),
            .I(N__59997));
    LocalMux I__13340 (
            .O(N__59997),
            .I(N__59994));
    Span4Mux_h I__13339 (
            .O(N__59994),
            .I(N__59991));
    Span4Mux_h I__13338 (
            .O(N__59991),
            .I(N__59988));
    Odrv4 I__13337 (
            .O(N__59988),
            .I(\c0.n30_adj_4545 ));
    InMux I__13336 (
            .O(N__59985),
            .I(N__59982));
    LocalMux I__13335 (
            .O(N__59982),
            .I(\c0.n72 ));
    InMux I__13334 (
            .O(N__59979),
            .I(N__59976));
    LocalMux I__13333 (
            .O(N__59976),
            .I(N__59973));
    Span4Mux_v I__13332 (
            .O(N__59973),
            .I(N__59970));
    Odrv4 I__13331 (
            .O(N__59970),
            .I(\c0.n24559 ));
    CascadeMux I__13330 (
            .O(N__59967),
            .I(N__59964));
    InMux I__13329 (
            .O(N__59964),
            .I(N__59961));
    LocalMux I__13328 (
            .O(N__59961),
            .I(N__59958));
    Odrv4 I__13327 (
            .O(N__59958),
            .I(\c0.n42_adj_4510 ));
    InMux I__13326 (
            .O(N__59955),
            .I(N__59952));
    LocalMux I__13325 (
            .O(N__59952),
            .I(\c0.n20_adj_4518 ));
    CascadeMux I__13324 (
            .O(N__59949),
            .I(N__59946));
    InMux I__13323 (
            .O(N__59946),
            .I(N__59943));
    LocalMux I__13322 (
            .O(N__59943),
            .I(N__59940));
    Span4Mux_h I__13321 (
            .O(N__59940),
            .I(N__59937));
    Odrv4 I__13320 (
            .O(N__59937),
            .I(\c0.n24751 ));
    CascadeMux I__13319 (
            .O(N__59934),
            .I(\c0.n14_adj_4676_cascade_ ));
    InMux I__13318 (
            .O(N__59931),
            .I(N__59928));
    LocalMux I__13317 (
            .O(N__59928),
            .I(N__59925));
    Span4Mux_h I__13316 (
            .O(N__59925),
            .I(N__59922));
    Odrv4 I__13315 (
            .O(N__59922),
            .I(\c0.data_out_frame_0__7__N_2777 ));
    InMux I__13314 (
            .O(N__59919),
            .I(N__59916));
    LocalMux I__13313 (
            .O(N__59916),
            .I(N__59913));
    Span4Mux_h I__13312 (
            .O(N__59913),
            .I(N__59909));
    InMux I__13311 (
            .O(N__59912),
            .I(N__59906));
    Odrv4 I__13310 (
            .O(N__59909),
            .I(\c0.n10_adj_4513 ));
    LocalMux I__13309 (
            .O(N__59906),
            .I(\c0.n10_adj_4513 ));
    InMux I__13308 (
            .O(N__59901),
            .I(N__59898));
    LocalMux I__13307 (
            .O(N__59898),
            .I(N__59893));
    InMux I__13306 (
            .O(N__59897),
            .I(N__59890));
    InMux I__13305 (
            .O(N__59896),
            .I(N__59887));
    Odrv4 I__13304 (
            .O(N__59893),
            .I(\c0.n15_adj_4497 ));
    LocalMux I__13303 (
            .O(N__59890),
            .I(\c0.n15_adj_4497 ));
    LocalMux I__13302 (
            .O(N__59887),
            .I(\c0.n15_adj_4497 ));
    CascadeMux I__13301 (
            .O(N__59880),
            .I(N__59877));
    InMux I__13300 (
            .O(N__59877),
            .I(N__59872));
    InMux I__13299 (
            .O(N__59876),
            .I(N__59869));
    CascadeMux I__13298 (
            .O(N__59875),
            .I(N__59864));
    LocalMux I__13297 (
            .O(N__59872),
            .I(N__59861));
    LocalMux I__13296 (
            .O(N__59869),
            .I(N__59858));
    InMux I__13295 (
            .O(N__59868),
            .I(N__59853));
    InMux I__13294 (
            .O(N__59867),
            .I(N__59853));
    InMux I__13293 (
            .O(N__59864),
            .I(N__59850));
    Span4Mux_h I__13292 (
            .O(N__59861),
            .I(N__59845));
    Span4Mux_h I__13291 (
            .O(N__59858),
            .I(N__59845));
    LocalMux I__13290 (
            .O(N__59853),
            .I(\c0.data_in_frame_25_4 ));
    LocalMux I__13289 (
            .O(N__59850),
            .I(\c0.data_in_frame_25_4 ));
    Odrv4 I__13288 (
            .O(N__59845),
            .I(\c0.data_in_frame_25_4 ));
    InMux I__13287 (
            .O(N__59838),
            .I(N__59835));
    LocalMux I__13286 (
            .O(N__59835),
            .I(N__59832));
    Span4Mux_v I__13285 (
            .O(N__59832),
            .I(N__59829));
    Odrv4 I__13284 (
            .O(N__59829),
            .I(\c0.n23_adj_4551 ));
    InMux I__13283 (
            .O(N__59826),
            .I(N__59823));
    LocalMux I__13282 (
            .O(N__59823),
            .I(\c0.n26_adj_4548 ));
    CascadeMux I__13281 (
            .O(N__59820),
            .I(\c0.n24_adj_4550_cascade_ ));
    CascadeMux I__13280 (
            .O(N__59817),
            .I(\c0.n21010_cascade_ ));
    InMux I__13279 (
            .O(N__59814),
            .I(N__59811));
    LocalMux I__13278 (
            .O(N__59811),
            .I(\c0.n53_adj_4538 ));
    InMux I__13277 (
            .O(N__59808),
            .I(N__59805));
    LocalMux I__13276 (
            .O(N__59805),
            .I(\c0.n61_adj_4543 ));
    InMux I__13275 (
            .O(N__59802),
            .I(N__59799));
    LocalMux I__13274 (
            .O(N__59799),
            .I(\c0.n42_adj_4540 ));
    CascadeMux I__13273 (
            .O(N__59796),
            .I(N__59793));
    InMux I__13272 (
            .O(N__59793),
            .I(N__59790));
    LocalMux I__13271 (
            .O(N__59790),
            .I(\c0.n62_adj_4541 ));
    CascadeMux I__13270 (
            .O(N__59787),
            .I(N__59783));
    InMux I__13269 (
            .O(N__59786),
            .I(N__59777));
    InMux I__13268 (
            .O(N__59783),
            .I(N__59777));
    InMux I__13267 (
            .O(N__59782),
            .I(N__59774));
    LocalMux I__13266 (
            .O(N__59777),
            .I(N__59771));
    LocalMux I__13265 (
            .O(N__59774),
            .I(N__59768));
    Odrv4 I__13264 (
            .O(N__59771),
            .I(\c0.n13_adj_4492 ));
    Odrv12 I__13263 (
            .O(N__59768),
            .I(\c0.n13_adj_4492 ));
    InMux I__13262 (
            .O(N__59763),
            .I(N__59760));
    LocalMux I__13261 (
            .O(N__59760),
            .I(N__59757));
    Odrv4 I__13260 (
            .O(N__59757),
            .I(\c0.n18_adj_4493 ));
    InMux I__13259 (
            .O(N__59754),
            .I(N__59751));
    LocalMux I__13258 (
            .O(N__59751),
            .I(N__59748));
    Odrv4 I__13257 (
            .O(N__59748),
            .I(\c0.n22_adj_4498 ));
    CascadeMux I__13256 (
            .O(N__59745),
            .I(\c0.n26_adj_4499_cascade_ ));
    InMux I__13255 (
            .O(N__59742),
            .I(N__59739));
    LocalMux I__13254 (
            .O(N__59739),
            .I(N__59735));
    InMux I__13253 (
            .O(N__59738),
            .I(N__59732));
    Span4Mux_v I__13252 (
            .O(N__59735),
            .I(N__59725));
    LocalMux I__13251 (
            .O(N__59732),
            .I(N__59725));
    CascadeMux I__13250 (
            .O(N__59731),
            .I(N__59721));
    InMux I__13249 (
            .O(N__59730),
            .I(N__59717));
    Span4Mux_h I__13248 (
            .O(N__59725),
            .I(N__59714));
    InMux I__13247 (
            .O(N__59724),
            .I(N__59711));
    InMux I__13246 (
            .O(N__59721),
            .I(N__59706));
    InMux I__13245 (
            .O(N__59720),
            .I(N__59706));
    LocalMux I__13244 (
            .O(N__59717),
            .I(N__59703));
    Span4Mux_v I__13243 (
            .O(N__59714),
            .I(N__59699));
    LocalMux I__13242 (
            .O(N__59711),
            .I(N__59692));
    LocalMux I__13241 (
            .O(N__59706),
            .I(N__59692));
    Sp12to4 I__13240 (
            .O(N__59703),
            .I(N__59692));
    InMux I__13239 (
            .O(N__59702),
            .I(N__59689));
    Span4Mux_v I__13238 (
            .O(N__59699),
            .I(N__59686));
    Span12Mux_v I__13237 (
            .O(N__59692),
            .I(N__59683));
    LocalMux I__13236 (
            .O(N__59689),
            .I(\c0.data_in_frame_20_4 ));
    Odrv4 I__13235 (
            .O(N__59686),
            .I(\c0.data_in_frame_20_4 ));
    Odrv12 I__13234 (
            .O(N__59683),
            .I(\c0.data_in_frame_20_4 ));
    InMux I__13233 (
            .O(N__59676),
            .I(N__59673));
    LocalMux I__13232 (
            .O(N__59673),
            .I(\c0.n30_adj_4357 ));
    CascadeMux I__13231 (
            .O(N__59670),
            .I(N__59667));
    InMux I__13230 (
            .O(N__59667),
            .I(N__59664));
    LocalMux I__13229 (
            .O(N__59664),
            .I(N__59660));
    InMux I__13228 (
            .O(N__59663),
            .I(N__59657));
    Span4Mux_h I__13227 (
            .O(N__59660),
            .I(N__59654));
    LocalMux I__13226 (
            .O(N__59657),
            .I(N__59651));
    Span4Mux_v I__13225 (
            .O(N__59654),
            .I(N__59648));
    Span4Mux_h I__13224 (
            .O(N__59651),
            .I(N__59645));
    Odrv4 I__13223 (
            .O(N__59648),
            .I(\c0.n22334 ));
    Odrv4 I__13222 (
            .O(N__59645),
            .I(\c0.n22334 ));
    CascadeMux I__13221 (
            .O(N__59640),
            .I(N__59637));
    InMux I__13220 (
            .O(N__59637),
            .I(N__59633));
    CascadeMux I__13219 (
            .O(N__59636),
            .I(N__59630));
    LocalMux I__13218 (
            .O(N__59633),
            .I(N__59625));
    InMux I__13217 (
            .O(N__59630),
            .I(N__59622));
    CascadeMux I__13216 (
            .O(N__59629),
            .I(N__59619));
    CascadeMux I__13215 (
            .O(N__59628),
            .I(N__59616));
    Span4Mux_v I__13214 (
            .O(N__59625),
            .I(N__59613));
    LocalMux I__13213 (
            .O(N__59622),
            .I(N__59610));
    InMux I__13212 (
            .O(N__59619),
            .I(N__59607));
    InMux I__13211 (
            .O(N__59616),
            .I(N__59604));
    Span4Mux_h I__13210 (
            .O(N__59613),
            .I(N__59601));
    Span4Mux_v I__13209 (
            .O(N__59610),
            .I(N__59598));
    LocalMux I__13208 (
            .O(N__59607),
            .I(\c0.data_in_frame_25_6 ));
    LocalMux I__13207 (
            .O(N__59604),
            .I(\c0.data_in_frame_25_6 ));
    Odrv4 I__13206 (
            .O(N__59601),
            .I(\c0.data_in_frame_25_6 ));
    Odrv4 I__13205 (
            .O(N__59598),
            .I(\c0.data_in_frame_25_6 ));
    InMux I__13204 (
            .O(N__59589),
            .I(N__59582));
    InMux I__13203 (
            .O(N__59588),
            .I(N__59582));
    CascadeMux I__13202 (
            .O(N__59587),
            .I(N__59579));
    LocalMux I__13201 (
            .O(N__59582),
            .I(N__59575));
    InMux I__13200 (
            .O(N__59579),
            .I(N__59570));
    InMux I__13199 (
            .O(N__59578),
            .I(N__59570));
    Span4Mux_h I__13198 (
            .O(N__59575),
            .I(N__59567));
    LocalMux I__13197 (
            .O(N__59570),
            .I(\c0.data_in_frame_24_3 ));
    Odrv4 I__13196 (
            .O(N__59567),
            .I(\c0.data_in_frame_24_3 ));
    InMux I__13195 (
            .O(N__59562),
            .I(N__59558));
    InMux I__13194 (
            .O(N__59561),
            .I(N__59553));
    LocalMux I__13193 (
            .O(N__59558),
            .I(N__59550));
    InMux I__13192 (
            .O(N__59557),
            .I(N__59545));
    InMux I__13191 (
            .O(N__59556),
            .I(N__59545));
    LocalMux I__13190 (
            .O(N__59553),
            .I(N__59542));
    Span4Mux_h I__13189 (
            .O(N__59550),
            .I(N__59539));
    LocalMux I__13188 (
            .O(N__59545),
            .I(\c0.n24547 ));
    Odrv4 I__13187 (
            .O(N__59542),
            .I(\c0.n24547 ));
    Odrv4 I__13186 (
            .O(N__59539),
            .I(\c0.n24547 ));
    CascadeMux I__13185 (
            .O(N__59532),
            .I(N__59529));
    InMux I__13184 (
            .O(N__59529),
            .I(N__59526));
    LocalMux I__13183 (
            .O(N__59526),
            .I(N__59521));
    InMux I__13182 (
            .O(N__59525),
            .I(N__59516));
    InMux I__13181 (
            .O(N__59524),
            .I(N__59516));
    Span4Mux_v I__13180 (
            .O(N__59521),
            .I(N__59513));
    LocalMux I__13179 (
            .O(N__59516),
            .I(\c0.n21353 ));
    Odrv4 I__13178 (
            .O(N__59513),
            .I(\c0.n21353 ));
    CascadeMux I__13177 (
            .O(N__59508),
            .I(\c0.n66_cascade_ ));
    InMux I__13176 (
            .O(N__59505),
            .I(N__59502));
    LocalMux I__13175 (
            .O(N__59502),
            .I(\c0.n75 ));
    InMux I__13174 (
            .O(N__59499),
            .I(N__59496));
    LocalMux I__13173 (
            .O(N__59496),
            .I(\c0.n46_adj_4461 ));
    InMux I__13172 (
            .O(N__59493),
            .I(N__59490));
    LocalMux I__13171 (
            .O(N__59490),
            .I(N__59487));
    Odrv12 I__13170 (
            .O(N__59487),
            .I(\c0.n4_adj_4347 ));
    InMux I__13169 (
            .O(N__59484),
            .I(N__59481));
    LocalMux I__13168 (
            .O(N__59481),
            .I(N__59476));
    InMux I__13167 (
            .O(N__59480),
            .I(N__59471));
    InMux I__13166 (
            .O(N__59479),
            .I(N__59471));
    Span4Mux_h I__13165 (
            .O(N__59476),
            .I(N__59468));
    LocalMux I__13164 (
            .O(N__59471),
            .I(\c0.data_in_frame_23_4 ));
    Odrv4 I__13163 (
            .O(N__59468),
            .I(\c0.data_in_frame_23_4 ));
    CascadeMux I__13162 (
            .O(N__59463),
            .I(\c0.n4_adj_4347_cascade_ ));
    CascadeMux I__13161 (
            .O(N__59460),
            .I(N__59457));
    InMux I__13160 (
            .O(N__59457),
            .I(N__59453));
    InMux I__13159 (
            .O(N__59456),
            .I(N__59450));
    LocalMux I__13158 (
            .O(N__59453),
            .I(\c0.data_in_frame_23_1 ));
    LocalMux I__13157 (
            .O(N__59450),
            .I(\c0.data_in_frame_23_1 ));
    CascadeMux I__13156 (
            .O(N__59445),
            .I(\c0.n30_adj_4357_cascade_ ));
    InMux I__13155 (
            .O(N__59442),
            .I(N__59435));
    InMux I__13154 (
            .O(N__59441),
            .I(N__59435));
    InMux I__13153 (
            .O(N__59440),
            .I(N__59430));
    LocalMux I__13152 (
            .O(N__59435),
            .I(N__59427));
    InMux I__13151 (
            .O(N__59434),
            .I(N__59424));
    InMux I__13150 (
            .O(N__59433),
            .I(N__59421));
    LocalMux I__13149 (
            .O(N__59430),
            .I(N__59418));
    Span4Mux_h I__13148 (
            .O(N__59427),
            .I(N__59415));
    LocalMux I__13147 (
            .O(N__59424),
            .I(N__59412));
    LocalMux I__13146 (
            .O(N__59421),
            .I(\c0.n14_adj_4356 ));
    Odrv4 I__13145 (
            .O(N__59418),
            .I(\c0.n14_adj_4356 ));
    Odrv4 I__13144 (
            .O(N__59415),
            .I(\c0.n14_adj_4356 ));
    Odrv4 I__13143 (
            .O(N__59412),
            .I(\c0.n14_adj_4356 ));
    InMux I__13142 (
            .O(N__59403),
            .I(N__59400));
    LocalMux I__13141 (
            .O(N__59400),
            .I(\c0.n40_adj_4359 ));
    CascadeMux I__13140 (
            .O(N__59397),
            .I(\c0.n42_adj_4358_cascade_ ));
    InMux I__13139 (
            .O(N__59394),
            .I(N__59391));
    LocalMux I__13138 (
            .O(N__59391),
            .I(N__59388));
    Odrv12 I__13137 (
            .O(N__59388),
            .I(\c0.n41_adj_4360 ));
    InMux I__13136 (
            .O(N__59385),
            .I(N__59382));
    LocalMux I__13135 (
            .O(N__59382),
            .I(\c0.n37_adj_4458 ));
    CascadeMux I__13134 (
            .O(N__59379),
            .I(\c0.n34_adj_4361_cascade_ ));
    InMux I__13133 (
            .O(N__59376),
            .I(N__59373));
    LocalMux I__13132 (
            .O(N__59373),
            .I(\c0.n14148 ));
    InMux I__13131 (
            .O(N__59370),
            .I(N__59367));
    LocalMux I__13130 (
            .O(N__59367),
            .I(N__59363));
    InMux I__13129 (
            .O(N__59366),
            .I(N__59360));
    Odrv12 I__13128 (
            .O(N__59363),
            .I(\c0.n9_adj_4208 ));
    LocalMux I__13127 (
            .O(N__59360),
            .I(\c0.n9_adj_4208 ));
    CascadeMux I__13126 (
            .O(N__59355),
            .I(\c0.n6_adj_4587_cascade_ ));
    InMux I__13125 (
            .O(N__59352),
            .I(N__59349));
    LocalMux I__13124 (
            .O(N__59349),
            .I(N__59345));
    InMux I__13123 (
            .O(N__59348),
            .I(N__59342));
    Span4Mux_h I__13122 (
            .O(N__59345),
            .I(N__59339));
    LocalMux I__13121 (
            .O(N__59342),
            .I(\c0.n13461 ));
    Odrv4 I__13120 (
            .O(N__59339),
            .I(\c0.n13461 ));
    CascadeMux I__13119 (
            .O(N__59334),
            .I(N__59330));
    InMux I__13118 (
            .O(N__59333),
            .I(N__59326));
    InMux I__13117 (
            .O(N__59330),
            .I(N__59321));
    InMux I__13116 (
            .O(N__59329),
            .I(N__59321));
    LocalMux I__13115 (
            .O(N__59326),
            .I(N__59316));
    LocalMux I__13114 (
            .O(N__59321),
            .I(N__59316));
    Sp12to4 I__13113 (
            .O(N__59316),
            .I(N__59313));
    Odrv12 I__13112 (
            .O(N__59313),
            .I(\c0.n13756 ));
    CascadeMux I__13111 (
            .O(N__59310),
            .I(\c0.n13461_cascade_ ));
    CascadeMux I__13110 (
            .O(N__59307),
            .I(\c0.n6227_cascade_ ));
    InMux I__13109 (
            .O(N__59304),
            .I(N__59301));
    LocalMux I__13108 (
            .O(N__59301),
            .I(N__59297));
    InMux I__13107 (
            .O(N__59300),
            .I(N__59294));
    Span4Mux_v I__13106 (
            .O(N__59297),
            .I(N__59289));
    LocalMux I__13105 (
            .O(N__59294),
            .I(N__59289));
    Odrv4 I__13104 (
            .O(N__59289),
            .I(\c0.n22173 ));
    InMux I__13103 (
            .O(N__59286),
            .I(N__59283));
    LocalMux I__13102 (
            .O(N__59283),
            .I(N__59277));
    InMux I__13101 (
            .O(N__59282),
            .I(N__59270));
    InMux I__13100 (
            .O(N__59281),
            .I(N__59270));
    InMux I__13099 (
            .O(N__59280),
            .I(N__59270));
    Odrv12 I__13098 (
            .O(N__59277),
            .I(\c0.n19_adj_4291 ));
    LocalMux I__13097 (
            .O(N__59270),
            .I(\c0.n19_adj_4291 ));
    CascadeMux I__13096 (
            .O(N__59265),
            .I(N__59262));
    InMux I__13095 (
            .O(N__59262),
            .I(N__59256));
    InMux I__13094 (
            .O(N__59261),
            .I(N__59253));
    InMux I__13093 (
            .O(N__59260),
            .I(N__59250));
    InMux I__13092 (
            .O(N__59259),
            .I(N__59247));
    LocalMux I__13091 (
            .O(N__59256),
            .I(N__59244));
    LocalMux I__13090 (
            .O(N__59253),
            .I(N__59240));
    LocalMux I__13089 (
            .O(N__59250),
            .I(N__59237));
    LocalMux I__13088 (
            .O(N__59247),
            .I(N__59232));
    Span4Mux_h I__13087 (
            .O(N__59244),
            .I(N__59232));
    CascadeMux I__13086 (
            .O(N__59243),
            .I(N__59228));
    Span4Mux_v I__13085 (
            .O(N__59240),
            .I(N__59225));
    Span4Mux_h I__13084 (
            .O(N__59237),
            .I(N__59220));
    Span4Mux_v I__13083 (
            .O(N__59232),
            .I(N__59220));
    InMux I__13082 (
            .O(N__59231),
            .I(N__59215));
    InMux I__13081 (
            .O(N__59228),
            .I(N__59215));
    Odrv4 I__13080 (
            .O(N__59225),
            .I(data_in_frame_14_6));
    Odrv4 I__13079 (
            .O(N__59220),
            .I(data_in_frame_14_6));
    LocalMux I__13078 (
            .O(N__59215),
            .I(data_in_frame_14_6));
    InMux I__13077 (
            .O(N__59208),
            .I(N__59202));
    InMux I__13076 (
            .O(N__59207),
            .I(N__59199));
    InMux I__13075 (
            .O(N__59206),
            .I(N__59194));
    InMux I__13074 (
            .O(N__59205),
            .I(N__59191));
    LocalMux I__13073 (
            .O(N__59202),
            .I(N__59187));
    LocalMux I__13072 (
            .O(N__59199),
            .I(N__59184));
    InMux I__13071 (
            .O(N__59198),
            .I(N__59179));
    InMux I__13070 (
            .O(N__59197),
            .I(N__59179));
    LocalMux I__13069 (
            .O(N__59194),
            .I(N__59176));
    LocalMux I__13068 (
            .O(N__59191),
            .I(N__59173));
    InMux I__13067 (
            .O(N__59190),
            .I(N__59170));
    Span4Mux_v I__13066 (
            .O(N__59187),
            .I(N__59165));
    Span4Mux_h I__13065 (
            .O(N__59184),
            .I(N__59165));
    LocalMux I__13064 (
            .O(N__59179),
            .I(N__59162));
    Span4Mux_h I__13063 (
            .O(N__59176),
            .I(N__59157));
    Span4Mux_h I__13062 (
            .O(N__59173),
            .I(N__59157));
    LocalMux I__13061 (
            .O(N__59170),
            .I(N__59154));
    Span4Mux_v I__13060 (
            .O(N__59165),
            .I(N__59149));
    Span4Mux_h I__13059 (
            .O(N__59162),
            .I(N__59149));
    Span4Mux_v I__13058 (
            .O(N__59157),
            .I(N__59143));
    Span4Mux_h I__13057 (
            .O(N__59154),
            .I(N__59143));
    Span4Mux_v I__13056 (
            .O(N__59149),
            .I(N__59140));
    InMux I__13055 (
            .O(N__59148),
            .I(N__59137));
    Odrv4 I__13054 (
            .O(N__59143),
            .I(n22118));
    Odrv4 I__13053 (
            .O(N__59140),
            .I(n22118));
    LocalMux I__13052 (
            .O(N__59137),
            .I(n22118));
    InMux I__13051 (
            .O(N__59130),
            .I(N__59126));
    InMux I__13050 (
            .O(N__59129),
            .I(N__59122));
    LocalMux I__13049 (
            .O(N__59126),
            .I(N__59119));
    InMux I__13048 (
            .O(N__59125),
            .I(N__59116));
    LocalMux I__13047 (
            .O(N__59122),
            .I(\c0.data_in_frame_19_3 ));
    Odrv4 I__13046 (
            .O(N__59119),
            .I(\c0.data_in_frame_19_3 ));
    LocalMux I__13045 (
            .O(N__59116),
            .I(\c0.data_in_frame_19_3 ));
    InMux I__13044 (
            .O(N__59109),
            .I(N__59106));
    LocalMux I__13043 (
            .O(N__59106),
            .I(N__59102));
    InMux I__13042 (
            .O(N__59105),
            .I(N__59099));
    Span4Mux_v I__13041 (
            .O(N__59102),
            .I(N__59096));
    LocalMux I__13040 (
            .O(N__59099),
            .I(N__59093));
    Odrv4 I__13039 (
            .O(N__59096),
            .I(\c0.n14088 ));
    Odrv12 I__13038 (
            .O(N__59093),
            .I(\c0.n14088 ));
    InMux I__13037 (
            .O(N__59088),
            .I(N__59085));
    LocalMux I__13036 (
            .O(N__59085),
            .I(\c0.n23300 ));
    InMux I__13035 (
            .O(N__59082),
            .I(N__59078));
    InMux I__13034 (
            .O(N__59081),
            .I(N__59075));
    LocalMux I__13033 (
            .O(N__59078),
            .I(N__59072));
    LocalMux I__13032 (
            .O(N__59075),
            .I(N__59069));
    Span4Mux_v I__13031 (
            .O(N__59072),
            .I(N__59064));
    Span4Mux_v I__13030 (
            .O(N__59069),
            .I(N__59064));
    Span4Mux_h I__13029 (
            .O(N__59064),
            .I(N__59061));
    Odrv4 I__13028 (
            .O(N__59061),
            .I(\c0.n6_adj_4577 ));
    CascadeMux I__13027 (
            .O(N__59058),
            .I(N__59054));
    InMux I__13026 (
            .O(N__59057),
            .I(N__59050));
    InMux I__13025 (
            .O(N__59054),
            .I(N__59047));
    InMux I__13024 (
            .O(N__59053),
            .I(N__59044));
    LocalMux I__13023 (
            .O(N__59050),
            .I(N__59039));
    LocalMux I__13022 (
            .O(N__59047),
            .I(N__59039));
    LocalMux I__13021 (
            .O(N__59044),
            .I(\c0.n22662 ));
    Odrv12 I__13020 (
            .O(N__59039),
            .I(\c0.n22662 ));
    CascadeMux I__13019 (
            .O(N__59034),
            .I(\c0.n23300_cascade_ ));
    InMux I__13018 (
            .O(N__59031),
            .I(N__59028));
    LocalMux I__13017 (
            .O(N__59028),
            .I(\c0.n21_adj_4594 ));
    InMux I__13016 (
            .O(N__59025),
            .I(N__59022));
    LocalMux I__13015 (
            .O(N__59022),
            .I(N__59019));
    Span4Mux_v I__13014 (
            .O(N__59019),
            .I(N__59015));
    InMux I__13013 (
            .O(N__59018),
            .I(N__59012));
    Span4Mux_h I__13012 (
            .O(N__59015),
            .I(N__59005));
    LocalMux I__13011 (
            .O(N__59012),
            .I(N__59005));
    CascadeMux I__13010 (
            .O(N__59011),
            .I(N__59002));
    InMux I__13009 (
            .O(N__59010),
            .I(N__58998));
    Span4Mux_v I__13008 (
            .O(N__59005),
            .I(N__58995));
    InMux I__13007 (
            .O(N__59002),
            .I(N__58990));
    InMux I__13006 (
            .O(N__59001),
            .I(N__58990));
    LocalMux I__13005 (
            .O(N__58998),
            .I(\c0.data_in_frame_12_4 ));
    Odrv4 I__13004 (
            .O(N__58995),
            .I(\c0.data_in_frame_12_4 ));
    LocalMux I__13003 (
            .O(N__58990),
            .I(\c0.data_in_frame_12_4 ));
    CascadeMux I__13002 (
            .O(N__58983),
            .I(\c0.n4_adj_4658_cascade_ ));
    InMux I__13001 (
            .O(N__58980),
            .I(N__58974));
    InMux I__13000 (
            .O(N__58979),
            .I(N__58974));
    LocalMux I__12999 (
            .O(N__58974),
            .I(N__58971));
    Span4Mux_v I__12998 (
            .O(N__58971),
            .I(N__58968));
    Span4Mux_h I__12997 (
            .O(N__58968),
            .I(N__58963));
    InMux I__12996 (
            .O(N__58967),
            .I(N__58960));
    InMux I__12995 (
            .O(N__58966),
            .I(N__58957));
    Span4Mux_v I__12994 (
            .O(N__58963),
            .I(N__58952));
    LocalMux I__12993 (
            .O(N__58960),
            .I(N__58952));
    LocalMux I__12992 (
            .O(N__58957),
            .I(N__58949));
    Span4Mux_v I__12991 (
            .O(N__58952),
            .I(N__58946));
    Span12Mux_h I__12990 (
            .O(N__58949),
            .I(N__58943));
    Odrv4 I__12989 (
            .O(N__58946),
            .I(\c0.n24433 ));
    Odrv12 I__12988 (
            .O(N__58943),
            .I(\c0.n24433 ));
    InMux I__12987 (
            .O(N__58938),
            .I(N__58934));
    CascadeMux I__12986 (
            .O(N__58937),
            .I(N__58931));
    LocalMux I__12985 (
            .O(N__58934),
            .I(N__58927));
    InMux I__12984 (
            .O(N__58931),
            .I(N__58924));
    CascadeMux I__12983 (
            .O(N__58930),
            .I(N__58921));
    Span4Mux_h I__12982 (
            .O(N__58927),
            .I(N__58918));
    LocalMux I__12981 (
            .O(N__58924),
            .I(N__58915));
    InMux I__12980 (
            .O(N__58921),
            .I(N__58912));
    Span4Mux_h I__12979 (
            .O(N__58918),
            .I(N__58907));
    Span4Mux_v I__12978 (
            .O(N__58915),
            .I(N__58907));
    LocalMux I__12977 (
            .O(N__58912),
            .I(\c0.data_in_frame_16_6 ));
    Odrv4 I__12976 (
            .O(N__58907),
            .I(\c0.data_in_frame_16_6 ));
    CascadeMux I__12975 (
            .O(N__58902),
            .I(\c0.n12_adj_4682_cascade_ ));
    InMux I__12974 (
            .O(N__58899),
            .I(N__58896));
    LocalMux I__12973 (
            .O(N__58896),
            .I(N__58893));
    Span4Mux_h I__12972 (
            .O(N__58893),
            .I(N__58887));
    InMux I__12971 (
            .O(N__58892),
            .I(N__58884));
    InMux I__12970 (
            .O(N__58891),
            .I(N__58879));
    InMux I__12969 (
            .O(N__58890),
            .I(N__58879));
    Odrv4 I__12968 (
            .O(N__58887),
            .I(\c0.n23390 ));
    LocalMux I__12967 (
            .O(N__58884),
            .I(\c0.n23390 ));
    LocalMux I__12966 (
            .O(N__58879),
            .I(\c0.n23390 ));
    InMux I__12965 (
            .O(N__58872),
            .I(N__58868));
    InMux I__12964 (
            .O(N__58871),
            .I(N__58865));
    LocalMux I__12963 (
            .O(N__58868),
            .I(N__58862));
    LocalMux I__12962 (
            .O(N__58865),
            .I(N__58859));
    Odrv12 I__12961 (
            .O(N__58862),
            .I(\c0.n22249 ));
    Odrv12 I__12960 (
            .O(N__58859),
            .I(\c0.n22249 ));
    InMux I__12959 (
            .O(N__58854),
            .I(N__58851));
    LocalMux I__12958 (
            .O(N__58851),
            .I(\c0.n10_adj_4315 ));
    CascadeMux I__12957 (
            .O(N__58848),
            .I(N__58844));
    InMux I__12956 (
            .O(N__58847),
            .I(N__58836));
    InMux I__12955 (
            .O(N__58844),
            .I(N__58836));
    InMux I__12954 (
            .O(N__58843),
            .I(N__58836));
    LocalMux I__12953 (
            .O(N__58836),
            .I(\c0.n24534 ));
    InMux I__12952 (
            .O(N__58833),
            .I(N__58830));
    LocalMux I__12951 (
            .O(N__58830),
            .I(N__58825));
    CascadeMux I__12950 (
            .O(N__58829),
            .I(N__58822));
    InMux I__12949 (
            .O(N__58828),
            .I(N__58818));
    Span4Mux_h I__12948 (
            .O(N__58825),
            .I(N__58815));
    InMux I__12947 (
            .O(N__58822),
            .I(N__58810));
    InMux I__12946 (
            .O(N__58821),
            .I(N__58810));
    LocalMux I__12945 (
            .O(N__58818),
            .I(\c0.data_in_frame_17_3 ));
    Odrv4 I__12944 (
            .O(N__58815),
            .I(\c0.data_in_frame_17_3 ));
    LocalMux I__12943 (
            .O(N__58810),
            .I(\c0.data_in_frame_17_3 ));
    InMux I__12942 (
            .O(N__58803),
            .I(N__58800));
    LocalMux I__12941 (
            .O(N__58800),
            .I(\c0.n4_adj_4345 ));
    CascadeMux I__12940 (
            .O(N__58797),
            .I(\c0.n24534_cascade_ ));
    InMux I__12939 (
            .O(N__58794),
            .I(N__58791));
    LocalMux I__12938 (
            .O(N__58791),
            .I(N__58788));
    Span4Mux_h I__12937 (
            .O(N__58788),
            .I(N__58785));
    Odrv4 I__12936 (
            .O(N__58785),
            .I(\c0.n12_adj_4346 ));
    CascadeMux I__12935 (
            .O(N__58782),
            .I(N__58779));
    InMux I__12934 (
            .O(N__58779),
            .I(N__58768));
    InMux I__12933 (
            .O(N__58778),
            .I(N__58768));
    InMux I__12932 (
            .O(N__58777),
            .I(N__58768));
    InMux I__12931 (
            .O(N__58776),
            .I(N__58764));
    InMux I__12930 (
            .O(N__58775),
            .I(N__58761));
    LocalMux I__12929 (
            .O(N__58768),
            .I(N__58758));
    InMux I__12928 (
            .O(N__58767),
            .I(N__58755));
    LocalMux I__12927 (
            .O(N__58764),
            .I(N__58752));
    LocalMux I__12926 (
            .O(N__58761),
            .I(N__58748));
    Span4Mux_v I__12925 (
            .O(N__58758),
            .I(N__58743));
    LocalMux I__12924 (
            .O(N__58755),
            .I(N__58743));
    Span4Mux_v I__12923 (
            .O(N__58752),
            .I(N__58740));
    InMux I__12922 (
            .O(N__58751),
            .I(N__58737));
    Span4Mux_v I__12921 (
            .O(N__58748),
            .I(N__58732));
    Span4Mux_h I__12920 (
            .O(N__58743),
            .I(N__58732));
    Odrv4 I__12919 (
            .O(N__58740),
            .I(\c0.n13329 ));
    LocalMux I__12918 (
            .O(N__58737),
            .I(\c0.n13329 ));
    Odrv4 I__12917 (
            .O(N__58732),
            .I(\c0.n13329 ));
    InMux I__12916 (
            .O(N__58725),
            .I(N__58722));
    LocalMux I__12915 (
            .O(N__58722),
            .I(\c0.n4_adj_4621 ));
    InMux I__12914 (
            .O(N__58719),
            .I(N__58716));
    LocalMux I__12913 (
            .O(N__58716),
            .I(N__58712));
    InMux I__12912 (
            .O(N__58715),
            .I(N__58709));
    Odrv4 I__12911 (
            .O(N__58712),
            .I(\c0.n12_adj_4500 ));
    LocalMux I__12910 (
            .O(N__58709),
            .I(\c0.n12_adj_4500 ));
    CascadeMux I__12909 (
            .O(N__58704),
            .I(\c0.n22514_cascade_ ));
    InMux I__12908 (
            .O(N__58701),
            .I(N__58697));
    InMux I__12907 (
            .O(N__58700),
            .I(N__58694));
    LocalMux I__12906 (
            .O(N__58697),
            .I(\c0.data_in_frame_16_1 ));
    LocalMux I__12905 (
            .O(N__58694),
            .I(\c0.data_in_frame_16_1 ));
    InMux I__12904 (
            .O(N__58689),
            .I(N__58686));
    LocalMux I__12903 (
            .O(N__58686),
            .I(N__58683));
    Span4Mux_v I__12902 (
            .O(N__58683),
            .I(N__58680));
    Span4Mux_h I__12901 (
            .O(N__58680),
            .I(N__58677));
    Odrv4 I__12900 (
            .O(N__58677),
            .I(\c0.n14_adj_4566 ));
    CascadeMux I__12899 (
            .O(N__58674),
            .I(\c0.n14165_cascade_ ));
    CascadeMux I__12898 (
            .O(N__58671),
            .I(N__58666));
    CascadeMux I__12897 (
            .O(N__58670),
            .I(N__58663));
    InMux I__12896 (
            .O(N__58669),
            .I(N__58659));
    InMux I__12895 (
            .O(N__58666),
            .I(N__58656));
    InMux I__12894 (
            .O(N__58663),
            .I(N__58651));
    InMux I__12893 (
            .O(N__58662),
            .I(N__58651));
    LocalMux I__12892 (
            .O(N__58659),
            .I(N__58646));
    LocalMux I__12891 (
            .O(N__58656),
            .I(N__58646));
    LocalMux I__12890 (
            .O(N__58651),
            .I(N__58643));
    Odrv12 I__12889 (
            .O(N__58646),
            .I(\c0.data_in_frame_17_2 ));
    Odrv4 I__12888 (
            .O(N__58643),
            .I(\c0.data_in_frame_17_2 ));
    CascadeMux I__12887 (
            .O(N__58638),
            .I(N__58635));
    InMux I__12886 (
            .O(N__58635),
            .I(N__58632));
    LocalMux I__12885 (
            .O(N__58632),
            .I(N__58629));
    Span4Mux_v I__12884 (
            .O(N__58629),
            .I(N__58626));
    Odrv4 I__12883 (
            .O(N__58626),
            .I(\c0.n22_adj_4622 ));
    CascadeMux I__12882 (
            .O(N__58623),
            .I(\c0.n22825_cascade_ ));
    InMux I__12881 (
            .O(N__58620),
            .I(N__58615));
    InMux I__12880 (
            .O(N__58619),
            .I(N__58611));
    InMux I__12879 (
            .O(N__58618),
            .I(N__58608));
    LocalMux I__12878 (
            .O(N__58615),
            .I(N__58605));
    InMux I__12877 (
            .O(N__58614),
            .I(N__58602));
    LocalMux I__12876 (
            .O(N__58611),
            .I(N__58599));
    LocalMux I__12875 (
            .O(N__58608),
            .I(N__58594));
    Span4Mux_h I__12874 (
            .O(N__58605),
            .I(N__58594));
    LocalMux I__12873 (
            .O(N__58602),
            .I(data_in_frame_14_0));
    Odrv12 I__12872 (
            .O(N__58599),
            .I(data_in_frame_14_0));
    Odrv4 I__12871 (
            .O(N__58594),
            .I(data_in_frame_14_0));
    InMux I__12870 (
            .O(N__58587),
            .I(N__58584));
    LocalMux I__12869 (
            .O(N__58584),
            .I(N__58581));
    Span4Mux_h I__12868 (
            .O(N__58581),
            .I(N__58578));
    Span4Mux_h I__12867 (
            .O(N__58578),
            .I(N__58575));
    Odrv4 I__12866 (
            .O(N__58575),
            .I(\c0.n136 ));
    CascadeMux I__12865 (
            .O(N__58572),
            .I(\c0.n22751_cascade_ ));
    InMux I__12864 (
            .O(N__58569),
            .I(N__58566));
    LocalMux I__12863 (
            .O(N__58566),
            .I(N__58563));
    Odrv4 I__12862 (
            .O(N__58563),
            .I(\c0.n107 ));
    InMux I__12861 (
            .O(N__58560),
            .I(N__58557));
    LocalMux I__12860 (
            .O(N__58557),
            .I(\c0.n149 ));
    InMux I__12859 (
            .O(N__58554),
            .I(N__58551));
    LocalMux I__12858 (
            .O(N__58551),
            .I(\c0.n140 ));
    InMux I__12857 (
            .O(N__58548),
            .I(N__58545));
    LocalMux I__12856 (
            .O(N__58545),
            .I(N__58541));
    InMux I__12855 (
            .O(N__58544),
            .I(N__58538));
    Span12Mux_h I__12854 (
            .O(N__58541),
            .I(N__58535));
    LocalMux I__12853 (
            .O(N__58538),
            .I(N__58532));
    Odrv12 I__12852 (
            .O(N__58535),
            .I(\c0.n22843 ));
    Odrv4 I__12851 (
            .O(N__58532),
            .I(\c0.n22843 ));
    InMux I__12850 (
            .O(N__58527),
            .I(N__58524));
    LocalMux I__12849 (
            .O(N__58524),
            .I(N__58520));
    InMux I__12848 (
            .O(N__58523),
            .I(N__58517));
    Span4Mux_v I__12847 (
            .O(N__58520),
            .I(N__58514));
    LocalMux I__12846 (
            .O(N__58517),
            .I(N__58511));
    Span4Mux_h I__12845 (
            .O(N__58514),
            .I(N__58506));
    Span4Mux_v I__12844 (
            .O(N__58511),
            .I(N__58506));
    Odrv4 I__12843 (
            .O(N__58506),
            .I(\c0.n22_adj_4245 ));
    CascadeMux I__12842 (
            .O(N__58503),
            .I(\c0.n23598_cascade_ ));
    InMux I__12841 (
            .O(N__58500),
            .I(N__58497));
    LocalMux I__12840 (
            .O(N__58497),
            .I(N__58493));
    InMux I__12839 (
            .O(N__58496),
            .I(N__58490));
    Odrv12 I__12838 (
            .O(N__58493),
            .I(\c0.n23611 ));
    LocalMux I__12837 (
            .O(N__58490),
            .I(\c0.n23611 ));
    CascadeMux I__12836 (
            .O(N__58485),
            .I(\c0.n9_adj_4208_cascade_ ));
    InMux I__12835 (
            .O(N__58482),
            .I(N__58479));
    LocalMux I__12834 (
            .O(N__58479),
            .I(N__58476));
    Span4Mux_v I__12833 (
            .O(N__58476),
            .I(N__58473));
    Span4Mux_h I__12832 (
            .O(N__58473),
            .I(N__58469));
    InMux I__12831 (
            .O(N__58472),
            .I(N__58466));
    Odrv4 I__12830 (
            .O(N__58469),
            .I(\c0.n22304 ));
    LocalMux I__12829 (
            .O(N__58466),
            .I(\c0.n22304 ));
    CascadeMux I__12828 (
            .O(N__58461),
            .I(\c0.n13892_cascade_ ));
    CascadeMux I__12827 (
            .O(N__58458),
            .I(N__58455));
    InMux I__12826 (
            .O(N__58455),
            .I(N__58452));
    LocalMux I__12825 (
            .O(N__58452),
            .I(N__58448));
    CascadeMux I__12824 (
            .O(N__58451),
            .I(N__58444));
    Span4Mux_v I__12823 (
            .O(N__58448),
            .I(N__58441));
    InMux I__12822 (
            .O(N__58447),
            .I(N__58438));
    InMux I__12821 (
            .O(N__58444),
            .I(N__58435));
    Span4Mux_h I__12820 (
            .O(N__58441),
            .I(N__58430));
    LocalMux I__12819 (
            .O(N__58438),
            .I(N__58430));
    LocalMux I__12818 (
            .O(N__58435),
            .I(\c0.data_in_frame_11_6 ));
    Odrv4 I__12817 (
            .O(N__58430),
            .I(\c0.data_in_frame_11_6 ));
    InMux I__12816 (
            .O(N__58425),
            .I(N__58422));
    LocalMux I__12815 (
            .O(N__58422),
            .I(\c0.n13892 ));
    InMux I__12814 (
            .O(N__58419),
            .I(N__58416));
    LocalMux I__12813 (
            .O(N__58416),
            .I(N__58413));
    Odrv12 I__12812 (
            .O(N__58413),
            .I(\c0.n31 ));
    CascadeMux I__12811 (
            .O(N__58410),
            .I(\c0.n31_cascade_ ));
    InMux I__12810 (
            .O(N__58407),
            .I(N__58404));
    LocalMux I__12809 (
            .O(N__58404),
            .I(N__58400));
    CascadeMux I__12808 (
            .O(N__58403),
            .I(N__58396));
    Span4Mux_v I__12807 (
            .O(N__58400),
            .I(N__58392));
    InMux I__12806 (
            .O(N__58399),
            .I(N__58387));
    InMux I__12805 (
            .O(N__58396),
            .I(N__58387));
    InMux I__12804 (
            .O(N__58395),
            .I(N__58384));
    Odrv4 I__12803 (
            .O(N__58392),
            .I(\c0.data_in_frame_10_0 ));
    LocalMux I__12802 (
            .O(N__58387),
            .I(\c0.data_in_frame_10_0 ));
    LocalMux I__12801 (
            .O(N__58384),
            .I(\c0.data_in_frame_10_0 ));
    InMux I__12800 (
            .O(N__58377),
            .I(N__58374));
    LocalMux I__12799 (
            .O(N__58374),
            .I(N__58369));
    InMux I__12798 (
            .O(N__58373),
            .I(N__58366));
    InMux I__12797 (
            .O(N__58372),
            .I(N__58363));
    Span4Mux_v I__12796 (
            .O(N__58369),
            .I(N__58360));
    LocalMux I__12795 (
            .O(N__58366),
            .I(N__58355));
    LocalMux I__12794 (
            .O(N__58363),
            .I(N__58355));
    Odrv4 I__12793 (
            .O(N__58360),
            .I(\c0.n28 ));
    Odrv12 I__12792 (
            .O(N__58355),
            .I(\c0.n28 ));
    CascadeMux I__12791 (
            .O(N__58350),
            .I(N__58347));
    InMux I__12790 (
            .O(N__58347),
            .I(N__58344));
    LocalMux I__12789 (
            .O(N__58344),
            .I(\c0.n24 ));
    InMux I__12788 (
            .O(N__58341),
            .I(N__58338));
    LocalMux I__12787 (
            .O(N__58338),
            .I(N__58335));
    Odrv4 I__12786 (
            .O(N__58335),
            .I(\c0.n16 ));
    InMux I__12785 (
            .O(N__58332),
            .I(N__58326));
    InMux I__12784 (
            .O(N__58331),
            .I(N__58326));
    LocalMux I__12783 (
            .O(N__58326),
            .I(data_in_frame_14_2));
    CascadeMux I__12782 (
            .O(N__58323),
            .I(N__58320));
    InMux I__12781 (
            .O(N__58320),
            .I(N__58317));
    LocalMux I__12780 (
            .O(N__58317),
            .I(\c0.n8_adj_4673 ));
    InMux I__12779 (
            .O(N__58314),
            .I(N__58308));
    InMux I__12778 (
            .O(N__58313),
            .I(N__58308));
    LocalMux I__12777 (
            .O(N__58308),
            .I(data_in_frame_6_2));
    InMux I__12776 (
            .O(N__58305),
            .I(N__58301));
    CascadeMux I__12775 (
            .O(N__58304),
            .I(N__58298));
    LocalMux I__12774 (
            .O(N__58301),
            .I(N__58295));
    InMux I__12773 (
            .O(N__58298),
            .I(N__58292));
    Span4Mux_v I__12772 (
            .O(N__58295),
            .I(N__58289));
    LocalMux I__12771 (
            .O(N__58292),
            .I(\c0.data_in_frame_13_0 ));
    Odrv4 I__12770 (
            .O(N__58289),
            .I(\c0.data_in_frame_13_0 ));
    CascadeMux I__12769 (
            .O(N__58284),
            .I(\c0.n22205_cascade_ ));
    InMux I__12768 (
            .O(N__58281),
            .I(N__58274));
    InMux I__12767 (
            .O(N__58280),
            .I(N__58274));
    InMux I__12766 (
            .O(N__58279),
            .I(N__58271));
    LocalMux I__12765 (
            .O(N__58274),
            .I(N__58268));
    LocalMux I__12764 (
            .O(N__58271),
            .I(\c0.n23491 ));
    Odrv4 I__12763 (
            .O(N__58268),
            .I(\c0.n23491 ));
    InMux I__12762 (
            .O(N__58263),
            .I(N__58260));
    LocalMux I__12761 (
            .O(N__58260),
            .I(N__58257));
    Span4Mux_h I__12760 (
            .O(N__58257),
            .I(N__58254));
    Span4Mux_v I__12759 (
            .O(N__58254),
            .I(N__58250));
    InMux I__12758 (
            .O(N__58253),
            .I(N__58247));
    Odrv4 I__12757 (
            .O(N__58250),
            .I(\c0.n17_adj_4224 ));
    LocalMux I__12756 (
            .O(N__58247),
            .I(\c0.n17_adj_4224 ));
    InMux I__12755 (
            .O(N__58242),
            .I(N__58239));
    LocalMux I__12754 (
            .O(N__58239),
            .I(N__58236));
    Span4Mux_v I__12753 (
            .O(N__58236),
            .I(N__58233));
    Odrv4 I__12752 (
            .O(N__58233),
            .I(\c0.n130 ));
    InMux I__12751 (
            .O(N__58230),
            .I(N__58227));
    LocalMux I__12750 (
            .O(N__58227),
            .I(N__58224));
    Span4Mux_v I__12749 (
            .O(N__58224),
            .I(N__58221));
    Span4Mux_h I__12748 (
            .O(N__58221),
            .I(N__58218));
    Sp12to4 I__12747 (
            .O(N__58218),
            .I(N__58215));
    Odrv12 I__12746 (
            .O(N__58215),
            .I(\c0.n14_adj_4707 ));
    InMux I__12745 (
            .O(N__58212),
            .I(N__58209));
    LocalMux I__12744 (
            .O(N__58209),
            .I(N__58206));
    Span4Mux_h I__12743 (
            .O(N__58206),
            .I(N__58203));
    Odrv4 I__12742 (
            .O(N__58203),
            .I(\c0.n15_adj_4710 ));
    CascadeMux I__12741 (
            .O(N__58200),
            .I(N__58196));
    InMux I__12740 (
            .O(N__58199),
            .I(N__58193));
    InMux I__12739 (
            .O(N__58196),
            .I(N__58190));
    LocalMux I__12738 (
            .O(N__58193),
            .I(N__58187));
    LocalMux I__12737 (
            .O(N__58190),
            .I(N__58184));
    Span4Mux_v I__12736 (
            .O(N__58187),
            .I(N__58181));
    Span12Mux_v I__12735 (
            .O(N__58184),
            .I(N__58178));
    Odrv4 I__12734 (
            .O(N__58181),
            .I(\c0.n22511 ));
    Odrv12 I__12733 (
            .O(N__58178),
            .I(\c0.n22511 ));
    CascadeMux I__12732 (
            .O(N__58173),
            .I(N__58170));
    InMux I__12731 (
            .O(N__58170),
            .I(N__58166));
    InMux I__12730 (
            .O(N__58169),
            .I(N__58163));
    LocalMux I__12729 (
            .O(N__58166),
            .I(N__58159));
    LocalMux I__12728 (
            .O(N__58163),
            .I(N__58156));
    InMux I__12727 (
            .O(N__58162),
            .I(N__58152));
    Span4Mux_v I__12726 (
            .O(N__58159),
            .I(N__58147));
    Span4Mux_v I__12725 (
            .O(N__58156),
            .I(N__58147));
    InMux I__12724 (
            .O(N__58155),
            .I(N__58144));
    LocalMux I__12723 (
            .O(N__58152),
            .I(\c0.n22_adj_4259 ));
    Odrv4 I__12722 (
            .O(N__58147),
            .I(\c0.n22_adj_4259 ));
    LocalMux I__12721 (
            .O(N__58144),
            .I(\c0.n22_adj_4259 ));
    InMux I__12720 (
            .O(N__58137),
            .I(N__58133));
    InMux I__12719 (
            .O(N__58136),
            .I(N__58129));
    LocalMux I__12718 (
            .O(N__58133),
            .I(N__58125));
    InMux I__12717 (
            .O(N__58132),
            .I(N__58122));
    LocalMux I__12716 (
            .O(N__58129),
            .I(N__58119));
    InMux I__12715 (
            .O(N__58128),
            .I(N__58116));
    Span4Mux_v I__12714 (
            .O(N__58125),
            .I(N__58113));
    LocalMux I__12713 (
            .O(N__58122),
            .I(N__58108));
    Span4Mux_v I__12712 (
            .O(N__58119),
            .I(N__58108));
    LocalMux I__12711 (
            .O(N__58116),
            .I(data_in_frame_6_1));
    Odrv4 I__12710 (
            .O(N__58113),
            .I(data_in_frame_6_1));
    Odrv4 I__12709 (
            .O(N__58108),
            .I(data_in_frame_6_1));
    CascadeMux I__12708 (
            .O(N__58101),
            .I(\c0.n18_adj_4314_cascade_ ));
    InMux I__12707 (
            .O(N__58098),
            .I(N__58094));
    InMux I__12706 (
            .O(N__58097),
            .I(N__58091));
    LocalMux I__12705 (
            .O(N__58094),
            .I(N__58087));
    LocalMux I__12704 (
            .O(N__58091),
            .I(N__58084));
    CascadeMux I__12703 (
            .O(N__58090),
            .I(N__58081));
    Span4Mux_h I__12702 (
            .O(N__58087),
            .I(N__58075));
    Span4Mux_v I__12701 (
            .O(N__58084),
            .I(N__58072));
    InMux I__12700 (
            .O(N__58081),
            .I(N__58063));
    InMux I__12699 (
            .O(N__58080),
            .I(N__58063));
    InMux I__12698 (
            .O(N__58079),
            .I(N__58063));
    InMux I__12697 (
            .O(N__58078),
            .I(N__58063));
    Odrv4 I__12696 (
            .O(N__58075),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__12695 (
            .O(N__58072),
            .I(\c0.data_in_frame_3_7 ));
    LocalMux I__12694 (
            .O(N__58063),
            .I(\c0.data_in_frame_3_7 ));
    InMux I__12693 (
            .O(N__58056),
            .I(N__58044));
    CascadeMux I__12692 (
            .O(N__58055),
            .I(N__58040));
    InMux I__12691 (
            .O(N__58054),
            .I(N__58037));
    InMux I__12690 (
            .O(N__58053),
            .I(N__58026));
    InMux I__12689 (
            .O(N__58052),
            .I(N__58026));
    InMux I__12688 (
            .O(N__58051),
            .I(N__58026));
    InMux I__12687 (
            .O(N__58050),
            .I(N__58026));
    InMux I__12686 (
            .O(N__58049),
            .I(N__58026));
    InMux I__12685 (
            .O(N__58048),
            .I(N__58021));
    InMux I__12684 (
            .O(N__58047),
            .I(N__58021));
    LocalMux I__12683 (
            .O(N__58044),
            .I(N__58018));
    InMux I__12682 (
            .O(N__58043),
            .I(N__58015));
    InMux I__12681 (
            .O(N__58040),
            .I(N__58009));
    LocalMux I__12680 (
            .O(N__58037),
            .I(N__58002));
    LocalMux I__12679 (
            .O(N__58026),
            .I(N__58002));
    LocalMux I__12678 (
            .O(N__58021),
            .I(N__58002));
    Span12Mux_h I__12677 (
            .O(N__58018),
            .I(N__57999));
    LocalMux I__12676 (
            .O(N__58015),
            .I(N__57996));
    InMux I__12675 (
            .O(N__58014),
            .I(N__57993));
    InMux I__12674 (
            .O(N__58013),
            .I(N__57988));
    InMux I__12673 (
            .O(N__58012),
            .I(N__57988));
    LocalMux I__12672 (
            .O(N__58009),
            .I(N__57983));
    Span4Mux_v I__12671 (
            .O(N__58002),
            .I(N__57983));
    Odrv12 I__12670 (
            .O(N__57999),
            .I(data_in_frame_1_6));
    Odrv4 I__12669 (
            .O(N__57996),
            .I(data_in_frame_1_6));
    LocalMux I__12668 (
            .O(N__57993),
            .I(data_in_frame_1_6));
    LocalMux I__12667 (
            .O(N__57988),
            .I(data_in_frame_1_6));
    Odrv4 I__12666 (
            .O(N__57983),
            .I(data_in_frame_1_6));
    InMux I__12665 (
            .O(N__57972),
            .I(N__57969));
    LocalMux I__12664 (
            .O(N__57969),
            .I(\c0.n38_adj_4448 ));
    InMux I__12663 (
            .O(N__57966),
            .I(N__57963));
    LocalMux I__12662 (
            .O(N__57963),
            .I(\c0.n42_adj_4449 ));
    InMux I__12661 (
            .O(N__57960),
            .I(N__57952));
    InMux I__12660 (
            .O(N__57959),
            .I(N__57952));
    InMux I__12659 (
            .O(N__57958),
            .I(N__57946));
    InMux I__12658 (
            .O(N__57957),
            .I(N__57943));
    LocalMux I__12657 (
            .O(N__57952),
            .I(N__57939));
    InMux I__12656 (
            .O(N__57951),
            .I(N__57934));
    InMux I__12655 (
            .O(N__57950),
            .I(N__57934));
    CascadeMux I__12654 (
            .O(N__57949),
            .I(N__57931));
    LocalMux I__12653 (
            .O(N__57946),
            .I(N__57925));
    LocalMux I__12652 (
            .O(N__57943),
            .I(N__57925));
    InMux I__12651 (
            .O(N__57942),
            .I(N__57922));
    Span4Mux_v I__12650 (
            .O(N__57939),
            .I(N__57917));
    LocalMux I__12649 (
            .O(N__57934),
            .I(N__57917));
    InMux I__12648 (
            .O(N__57931),
            .I(N__57912));
    InMux I__12647 (
            .O(N__57930),
            .I(N__57912));
    Span4Mux_h I__12646 (
            .O(N__57925),
            .I(N__57909));
    LocalMux I__12645 (
            .O(N__57922),
            .I(\c0.data_in_frame_3_3 ));
    Odrv4 I__12644 (
            .O(N__57917),
            .I(\c0.data_in_frame_3_3 ));
    LocalMux I__12643 (
            .O(N__57912),
            .I(\c0.data_in_frame_3_3 ));
    Odrv4 I__12642 (
            .O(N__57909),
            .I(\c0.data_in_frame_3_3 ));
    InMux I__12641 (
            .O(N__57900),
            .I(N__57897));
    LocalMux I__12640 (
            .O(N__57897),
            .I(N__57894));
    Span4Mux_h I__12639 (
            .O(N__57894),
            .I(N__57891));
    Odrv4 I__12638 (
            .O(N__57891),
            .I(\c0.n24_adj_4689 ));
    InMux I__12637 (
            .O(N__57888),
            .I(N__57883));
    InMux I__12636 (
            .O(N__57887),
            .I(N__57878));
    InMux I__12635 (
            .O(N__57886),
            .I(N__57878));
    LocalMux I__12634 (
            .O(N__57883),
            .I(N__57875));
    LocalMux I__12633 (
            .O(N__57878),
            .I(N__57872));
    Span4Mux_h I__12632 (
            .O(N__57875),
            .I(N__57869));
    Odrv4 I__12631 (
            .O(N__57872),
            .I(\c0.n13_adj_4281 ));
    Odrv4 I__12630 (
            .O(N__57869),
            .I(\c0.n13_adj_4281 ));
    InMux I__12629 (
            .O(N__57864),
            .I(N__57861));
    LocalMux I__12628 (
            .O(N__57861),
            .I(N__57858));
    Odrv4 I__12627 (
            .O(N__57858),
            .I(\c0.n102_adj_4445 ));
    InMux I__12626 (
            .O(N__57855),
            .I(N__57852));
    LocalMux I__12625 (
            .O(N__57852),
            .I(\c0.n101 ));
    InMux I__12624 (
            .O(N__57849),
            .I(N__57846));
    LocalMux I__12623 (
            .O(N__57846),
            .I(\c0.n103 ));
    InMux I__12622 (
            .O(N__57843),
            .I(N__57840));
    LocalMux I__12621 (
            .O(N__57840),
            .I(\c0.n98 ));
    InMux I__12620 (
            .O(N__57837),
            .I(N__57834));
    LocalMux I__12619 (
            .O(N__57834),
            .I(N__57831));
    Span4Mux_v I__12618 (
            .O(N__57831),
            .I(N__57828));
    Odrv4 I__12617 (
            .O(N__57828),
            .I(\c0.n97 ));
    CascadeMux I__12616 (
            .O(N__57825),
            .I(\c0.n110_cascade_ ));
    InMux I__12615 (
            .O(N__57822),
            .I(N__57819));
    LocalMux I__12614 (
            .O(N__57819),
            .I(\c0.n24465 ));
    InMux I__12613 (
            .O(N__57816),
            .I(N__57813));
    LocalMux I__12612 (
            .O(N__57813),
            .I(N__57810));
    Span4Mux_v I__12611 (
            .O(N__57810),
            .I(N__57807));
    Span4Mux_h I__12610 (
            .O(N__57807),
            .I(N__57804));
    Odrv4 I__12609 (
            .O(N__57804),
            .I(\c0.data_out_frame_0__7__N_2579 ));
    InMux I__12608 (
            .O(N__57801),
            .I(N__57797));
    CascadeMux I__12607 (
            .O(N__57800),
            .I(N__57794));
    LocalMux I__12606 (
            .O(N__57797),
            .I(N__57791));
    InMux I__12605 (
            .O(N__57794),
            .I(N__57788));
    Odrv4 I__12604 (
            .O(N__57791),
            .I(\c0.n15_adj_4450 ));
    LocalMux I__12603 (
            .O(N__57788),
            .I(\c0.n15_adj_4450 ));
    CascadeMux I__12602 (
            .O(N__57783),
            .I(N__57779));
    InMux I__12601 (
            .O(N__57782),
            .I(N__57776));
    InMux I__12600 (
            .O(N__57779),
            .I(N__57773));
    LocalMux I__12599 (
            .O(N__57776),
            .I(N__57768));
    LocalMux I__12598 (
            .O(N__57773),
            .I(N__57768));
    Odrv12 I__12597 (
            .O(N__57768),
            .I(\c0.n87 ));
    InMux I__12596 (
            .O(N__57765),
            .I(N__57762));
    LocalMux I__12595 (
            .O(N__57762),
            .I(N__57759));
    Span4Mux_v I__12594 (
            .O(N__57759),
            .I(N__57756));
    Odrv4 I__12593 (
            .O(N__57756),
            .I(\c0.n85 ));
    InMux I__12592 (
            .O(N__57753),
            .I(N__57750));
    LocalMux I__12591 (
            .O(N__57750),
            .I(N__57747));
    Span4Mux_h I__12590 (
            .O(N__57747),
            .I(N__57744));
    Odrv4 I__12589 (
            .O(N__57744),
            .I(\c0.n88 ));
    CascadeMux I__12588 (
            .O(N__57741),
            .I(\c0.n87_cascade_ ));
    InMux I__12587 (
            .O(N__57738),
            .I(N__57735));
    LocalMux I__12586 (
            .O(N__57735),
            .I(\c0.n106 ));
    InMux I__12585 (
            .O(N__57732),
            .I(N__57725));
    InMux I__12584 (
            .O(N__57731),
            .I(N__57722));
    InMux I__12583 (
            .O(N__57730),
            .I(N__57714));
    InMux I__12582 (
            .O(N__57729),
            .I(N__57714));
    InMux I__12581 (
            .O(N__57728),
            .I(N__57714));
    LocalMux I__12580 (
            .O(N__57725),
            .I(N__57711));
    LocalMux I__12579 (
            .O(N__57722),
            .I(N__57708));
    InMux I__12578 (
            .O(N__57721),
            .I(N__57705));
    LocalMux I__12577 (
            .O(N__57714),
            .I(N__57702));
    Span4Mux_v I__12576 (
            .O(N__57711),
            .I(N__57699));
    Span4Mux_v I__12575 (
            .O(N__57708),
            .I(N__57694));
    LocalMux I__12574 (
            .O(N__57705),
            .I(N__57694));
    Span4Mux_h I__12573 (
            .O(N__57702),
            .I(N__57691));
    Odrv4 I__12572 (
            .O(N__57699),
            .I(\c0.n22160 ));
    Odrv4 I__12571 (
            .O(N__57694),
            .I(\c0.n22160 ));
    Odrv4 I__12570 (
            .O(N__57691),
            .I(\c0.n22160 ));
    InMux I__12569 (
            .O(N__57684),
            .I(N__57678));
    InMux I__12568 (
            .O(N__57683),
            .I(N__57678));
    LocalMux I__12567 (
            .O(N__57678),
            .I(\c0.n7_adj_4304 ));
    CascadeMux I__12566 (
            .O(N__57675),
            .I(\c0.n7_adj_4304_cascade_ ));
    CascadeMux I__12565 (
            .O(N__57672),
            .I(N__57668));
    CascadeMux I__12564 (
            .O(N__57671),
            .I(N__57664));
    InMux I__12563 (
            .O(N__57668),
            .I(N__57658));
    InMux I__12562 (
            .O(N__57667),
            .I(N__57655));
    InMux I__12561 (
            .O(N__57664),
            .I(N__57650));
    InMux I__12560 (
            .O(N__57663),
            .I(N__57650));
    InMux I__12559 (
            .O(N__57662),
            .I(N__57647));
    InMux I__12558 (
            .O(N__57661),
            .I(N__57644));
    LocalMux I__12557 (
            .O(N__57658),
            .I(N__57639));
    LocalMux I__12556 (
            .O(N__57655),
            .I(N__57639));
    LocalMux I__12555 (
            .O(N__57650),
            .I(N__57633));
    LocalMux I__12554 (
            .O(N__57647),
            .I(N__57628));
    LocalMux I__12553 (
            .O(N__57644),
            .I(N__57628));
    Span4Mux_h I__12552 (
            .O(N__57639),
            .I(N__57625));
    InMux I__12551 (
            .O(N__57638),
            .I(N__57620));
    InMux I__12550 (
            .O(N__57637),
            .I(N__57620));
    InMux I__12549 (
            .O(N__57636),
            .I(N__57617));
    Odrv12 I__12548 (
            .O(N__57633),
            .I(data_in_frame_5_7));
    Odrv12 I__12547 (
            .O(N__57628),
            .I(data_in_frame_5_7));
    Odrv4 I__12546 (
            .O(N__57625),
            .I(data_in_frame_5_7));
    LocalMux I__12545 (
            .O(N__57620),
            .I(data_in_frame_5_7));
    LocalMux I__12544 (
            .O(N__57617),
            .I(data_in_frame_5_7));
    InMux I__12543 (
            .O(N__57606),
            .I(N__57603));
    LocalMux I__12542 (
            .O(N__57603),
            .I(N__57600));
    Span4Mux_h I__12541 (
            .O(N__57600),
            .I(N__57597));
    Sp12to4 I__12540 (
            .O(N__57597),
            .I(N__57594));
    Span12Mux_v I__12539 (
            .O(N__57594),
            .I(N__57589));
    InMux I__12538 (
            .O(N__57593),
            .I(N__57584));
    InMux I__12537 (
            .O(N__57592),
            .I(N__57584));
    Odrv12 I__12536 (
            .O(N__57589),
            .I(data_in_frame_6_0));
    LocalMux I__12535 (
            .O(N__57584),
            .I(data_in_frame_6_0));
    InMux I__12534 (
            .O(N__57579),
            .I(N__57576));
    LocalMux I__12533 (
            .O(N__57576),
            .I(N__57573));
    Span4Mux_v I__12532 (
            .O(N__57573),
            .I(N__57570));
    Span4Mux_h I__12531 (
            .O(N__57570),
            .I(N__57567));
    Odrv4 I__12530 (
            .O(N__57567),
            .I(\c0.n27_adj_4725 ));
    InMux I__12529 (
            .O(N__57564),
            .I(N__57559));
    InMux I__12528 (
            .O(N__57563),
            .I(N__57554));
    InMux I__12527 (
            .O(N__57562),
            .I(N__57554));
    LocalMux I__12526 (
            .O(N__57559),
            .I(N__57551));
    LocalMux I__12525 (
            .O(N__57554),
            .I(N__57548));
    Span4Mux_h I__12524 (
            .O(N__57551),
            .I(N__57545));
    Span4Mux_v I__12523 (
            .O(N__57548),
            .I(N__57542));
    Odrv4 I__12522 (
            .O(N__57545),
            .I(\c0.n13453 ));
    Odrv4 I__12521 (
            .O(N__57542),
            .I(\c0.n13453 ));
    InMux I__12520 (
            .O(N__57537),
            .I(N__57532));
    InMux I__12519 (
            .O(N__57536),
            .I(N__57529));
    CascadeMux I__12518 (
            .O(N__57535),
            .I(N__57526));
    LocalMux I__12517 (
            .O(N__57532),
            .I(N__57523));
    LocalMux I__12516 (
            .O(N__57529),
            .I(N__57520));
    InMux I__12515 (
            .O(N__57526),
            .I(N__57517));
    Odrv4 I__12514 (
            .O(N__57523),
            .I(\c0.n13_adj_4584 ));
    Odrv12 I__12513 (
            .O(N__57520),
            .I(\c0.n13_adj_4584 ));
    LocalMux I__12512 (
            .O(N__57517),
            .I(\c0.n13_adj_4584 ));
    CascadeMux I__12511 (
            .O(N__57510),
            .I(\c0.n15_adj_4444_cascade_ ));
    InMux I__12510 (
            .O(N__57507),
            .I(N__57504));
    LocalMux I__12509 (
            .O(N__57504),
            .I(N__57501));
    Span4Mux_h I__12508 (
            .O(N__57501),
            .I(N__57498));
    Odrv4 I__12507 (
            .O(N__57498),
            .I(\c0.n11_adj_4656 ));
    InMux I__12506 (
            .O(N__57495),
            .I(N__57489));
    InMux I__12505 (
            .O(N__57494),
            .I(N__57489));
    LocalMux I__12504 (
            .O(N__57489),
            .I(N__57485));
    CascadeMux I__12503 (
            .O(N__57488),
            .I(N__57480));
    Span4Mux_h I__12502 (
            .O(N__57485),
            .I(N__57477));
    InMux I__12501 (
            .O(N__57484),
            .I(N__57474));
    InMux I__12500 (
            .O(N__57483),
            .I(N__57469));
    InMux I__12499 (
            .O(N__57480),
            .I(N__57469));
    Odrv4 I__12498 (
            .O(N__57477),
            .I(\c0.data_in_frame_3_2 ));
    LocalMux I__12497 (
            .O(N__57474),
            .I(\c0.data_in_frame_3_2 ));
    LocalMux I__12496 (
            .O(N__57469),
            .I(\c0.data_in_frame_3_2 ));
    CascadeMux I__12495 (
            .O(N__57462),
            .I(N__57457));
    InMux I__12494 (
            .O(N__57461),
            .I(N__57450));
    InMux I__12493 (
            .O(N__57460),
            .I(N__57450));
    InMux I__12492 (
            .O(N__57457),
            .I(N__57450));
    LocalMux I__12491 (
            .O(N__57450),
            .I(data_in_frame_5_4));
    CascadeMux I__12490 (
            .O(N__57447),
            .I(N__57444));
    InMux I__12489 (
            .O(N__57444),
            .I(N__57441));
    LocalMux I__12488 (
            .O(N__57441),
            .I(\c0.n6_adj_4611 ));
    CascadeMux I__12487 (
            .O(N__57438),
            .I(\c0.n6_adj_4611_cascade_ ));
    InMux I__12486 (
            .O(N__57435),
            .I(N__57432));
    LocalMux I__12485 (
            .O(N__57432),
            .I(N__57429));
    Span4Mux_v I__12484 (
            .O(N__57429),
            .I(N__57425));
    InMux I__12483 (
            .O(N__57428),
            .I(N__57422));
    Odrv4 I__12482 (
            .O(N__57425),
            .I(\c0.n91 ));
    LocalMux I__12481 (
            .O(N__57422),
            .I(\c0.n91 ));
    CascadeMux I__12480 (
            .O(N__57417),
            .I(N__57413));
    InMux I__12479 (
            .O(N__57416),
            .I(N__57410));
    InMux I__12478 (
            .O(N__57413),
            .I(N__57406));
    LocalMux I__12477 (
            .O(N__57410),
            .I(N__57403));
    CascadeMux I__12476 (
            .O(N__57409),
            .I(N__57400));
    LocalMux I__12475 (
            .O(N__57406),
            .I(N__57396));
    Span4Mux_v I__12474 (
            .O(N__57403),
            .I(N__57393));
    InMux I__12473 (
            .O(N__57400),
            .I(N__57388));
    InMux I__12472 (
            .O(N__57399),
            .I(N__57388));
    Odrv4 I__12471 (
            .O(N__57396),
            .I(\c0.data_in_frame_9_6 ));
    Odrv4 I__12470 (
            .O(N__57393),
            .I(\c0.data_in_frame_9_6 ));
    LocalMux I__12469 (
            .O(N__57388),
            .I(\c0.data_in_frame_9_6 ));
    InMux I__12468 (
            .O(N__57381),
            .I(N__57378));
    LocalMux I__12467 (
            .O(N__57378),
            .I(N__57373));
    InMux I__12466 (
            .O(N__57377),
            .I(N__57370));
    CascadeMux I__12465 (
            .O(N__57376),
            .I(N__57367));
    Span4Mux_h I__12464 (
            .O(N__57373),
            .I(N__57362));
    LocalMux I__12463 (
            .O(N__57370),
            .I(N__57359));
    InMux I__12462 (
            .O(N__57367),
            .I(N__57356));
    InMux I__12461 (
            .O(N__57366),
            .I(N__57352));
    InMux I__12460 (
            .O(N__57365),
            .I(N__57349));
    Span4Mux_v I__12459 (
            .O(N__57362),
            .I(N__57346));
    Span4Mux_v I__12458 (
            .O(N__57359),
            .I(N__57343));
    LocalMux I__12457 (
            .O(N__57356),
            .I(N__57340));
    InMux I__12456 (
            .O(N__57355),
            .I(N__57337));
    LocalMux I__12455 (
            .O(N__57352),
            .I(data_in_frame_5_3));
    LocalMux I__12454 (
            .O(N__57349),
            .I(data_in_frame_5_3));
    Odrv4 I__12453 (
            .O(N__57346),
            .I(data_in_frame_5_3));
    Odrv4 I__12452 (
            .O(N__57343),
            .I(data_in_frame_5_3));
    Odrv12 I__12451 (
            .O(N__57340),
            .I(data_in_frame_5_3));
    LocalMux I__12450 (
            .O(N__57337),
            .I(data_in_frame_5_3));
    InMux I__12449 (
            .O(N__57324),
            .I(N__57319));
    InMux I__12448 (
            .O(N__57323),
            .I(N__57314));
    InMux I__12447 (
            .O(N__57322),
            .I(N__57314));
    LocalMux I__12446 (
            .O(N__57319),
            .I(data_in_frame_5_2));
    LocalMux I__12445 (
            .O(N__57314),
            .I(data_in_frame_5_2));
    CascadeMux I__12444 (
            .O(N__57309),
            .I(N__57305));
    CascadeMux I__12443 (
            .O(N__57308),
            .I(N__57302));
    InMux I__12442 (
            .O(N__57305),
            .I(N__57299));
    InMux I__12441 (
            .O(N__57302),
            .I(N__57294));
    LocalMux I__12440 (
            .O(N__57299),
            .I(N__57291));
    InMux I__12439 (
            .O(N__57298),
            .I(N__57286));
    InMux I__12438 (
            .O(N__57297),
            .I(N__57286));
    LocalMux I__12437 (
            .O(N__57294),
            .I(N__57283));
    Span4Mux_h I__12436 (
            .O(N__57291),
            .I(N__57280));
    LocalMux I__12435 (
            .O(N__57286),
            .I(N__57277));
    Odrv4 I__12434 (
            .O(N__57283),
            .I(\c0.data_in_frame_7_6 ));
    Odrv4 I__12433 (
            .O(N__57280),
            .I(\c0.data_in_frame_7_6 ));
    Odrv12 I__12432 (
            .O(N__57277),
            .I(\c0.data_in_frame_7_6 ));
    InMux I__12431 (
            .O(N__57270),
            .I(N__57267));
    LocalMux I__12430 (
            .O(N__57267),
            .I(N__57264));
    Span4Mux_v I__12429 (
            .O(N__57264),
            .I(N__57260));
    CascadeMux I__12428 (
            .O(N__57263),
            .I(N__57257));
    Span4Mux_h I__12427 (
            .O(N__57260),
            .I(N__57254));
    InMux I__12426 (
            .O(N__57257),
            .I(N__57251));
    Span4Mux_v I__12425 (
            .O(N__57254),
            .I(N__57246));
    LocalMux I__12424 (
            .O(N__57251),
            .I(N__57246));
    Span4Mux_v I__12423 (
            .O(N__57246),
            .I(N__57240));
    InMux I__12422 (
            .O(N__57245),
            .I(N__57237));
    CascadeMux I__12421 (
            .O(N__57244),
            .I(N__57229));
    InMux I__12420 (
            .O(N__57243),
            .I(N__57225));
    Sp12to4 I__12419 (
            .O(N__57240),
            .I(N__57220));
    LocalMux I__12418 (
            .O(N__57237),
            .I(N__57220));
    InMux I__12417 (
            .O(N__57236),
            .I(N__57213));
    InMux I__12416 (
            .O(N__57235),
            .I(N__57213));
    InMux I__12415 (
            .O(N__57234),
            .I(N__57213));
    InMux I__12414 (
            .O(N__57233),
            .I(N__57208));
    InMux I__12413 (
            .O(N__57232),
            .I(N__57208));
    InMux I__12412 (
            .O(N__57229),
            .I(N__57203));
    InMux I__12411 (
            .O(N__57228),
            .I(N__57203));
    LocalMux I__12410 (
            .O(N__57225),
            .I(data_in_frame_1_2));
    Odrv12 I__12409 (
            .O(N__57220),
            .I(data_in_frame_1_2));
    LocalMux I__12408 (
            .O(N__57213),
            .I(data_in_frame_1_2));
    LocalMux I__12407 (
            .O(N__57208),
            .I(data_in_frame_1_2));
    LocalMux I__12406 (
            .O(N__57203),
            .I(data_in_frame_1_2));
    InMux I__12405 (
            .O(N__57192),
            .I(N__57189));
    LocalMux I__12404 (
            .O(N__57189),
            .I(\c0.n12_adj_4612 ));
    InMux I__12403 (
            .O(N__57186),
            .I(N__57183));
    LocalMux I__12402 (
            .O(N__57183),
            .I(N__57180));
    Span4Mux_h I__12401 (
            .O(N__57180),
            .I(N__57177));
    Odrv4 I__12400 (
            .O(N__57177),
            .I(\c0.n15_adj_4444 ));
    InMux I__12399 (
            .O(N__57174),
            .I(N__57171));
    LocalMux I__12398 (
            .O(N__57171),
            .I(N__57168));
    Span4Mux_h I__12397 (
            .O(N__57168),
            .I(N__57165));
    Odrv4 I__12396 (
            .O(N__57165),
            .I(\c0.n70_adj_4514 ));
    CascadeMux I__12395 (
            .O(N__57162),
            .I(\c0.n71_cascade_ ));
    CascadeMux I__12394 (
            .O(N__57159),
            .I(N__57156));
    InMux I__12393 (
            .O(N__57156),
            .I(N__57152));
    InMux I__12392 (
            .O(N__57155),
            .I(N__57149));
    LocalMux I__12391 (
            .O(N__57152),
            .I(N__57146));
    LocalMux I__12390 (
            .O(N__57149),
            .I(N__57143));
    Span4Mux_h I__12389 (
            .O(N__57146),
            .I(N__57140));
    Span12Mux_v I__12388 (
            .O(N__57143),
            .I(N__57137));
    Span4Mux_h I__12387 (
            .O(N__57140),
            .I(N__57134));
    Odrv12 I__12386 (
            .O(N__57137),
            .I(\c0.n17537 ));
    Odrv4 I__12385 (
            .O(N__57134),
            .I(\c0.n17537 ));
    CascadeMux I__12384 (
            .O(N__57129),
            .I(\c0.n81_cascade_ ));
    InMux I__12383 (
            .O(N__57126),
            .I(N__57123));
    LocalMux I__12382 (
            .O(N__57123),
            .I(\c0.n82_adj_4517 ));
    InMux I__12381 (
            .O(N__57120),
            .I(N__57117));
    LocalMux I__12380 (
            .O(N__57117),
            .I(\c0.n28_adj_4523 ));
    InMux I__12379 (
            .O(N__57114),
            .I(N__57109));
    InMux I__12378 (
            .O(N__57113),
            .I(N__57106));
    CascadeMux I__12377 (
            .O(N__57112),
            .I(N__57103));
    LocalMux I__12376 (
            .O(N__57109),
            .I(N__57099));
    LocalMux I__12375 (
            .O(N__57106),
            .I(N__57096));
    InMux I__12374 (
            .O(N__57103),
            .I(N__57091));
    InMux I__12373 (
            .O(N__57102),
            .I(N__57091));
    Span4Mux_h I__12372 (
            .O(N__57099),
            .I(N__57088));
    Odrv12 I__12371 (
            .O(N__57096),
            .I(\c0.data_in_frame_27_3 ));
    LocalMux I__12370 (
            .O(N__57091),
            .I(\c0.data_in_frame_27_3 ));
    Odrv4 I__12369 (
            .O(N__57088),
            .I(\c0.data_in_frame_27_3 ));
    CascadeMux I__12368 (
            .O(N__57081),
            .I(N__57077));
    InMux I__12367 (
            .O(N__57080),
            .I(N__57073));
    InMux I__12366 (
            .O(N__57077),
            .I(N__57069));
    InMux I__12365 (
            .O(N__57076),
            .I(N__57066));
    LocalMux I__12364 (
            .O(N__57073),
            .I(N__57063));
    InMux I__12363 (
            .O(N__57072),
            .I(N__57060));
    LocalMux I__12362 (
            .O(N__57069),
            .I(N__57053));
    LocalMux I__12361 (
            .O(N__57066),
            .I(N__57053));
    Span4Mux_v I__12360 (
            .O(N__57063),
            .I(N__57053));
    LocalMux I__12359 (
            .O(N__57060),
            .I(\c0.data_in_frame_27_4 ));
    Odrv4 I__12358 (
            .O(N__57053),
            .I(\c0.data_in_frame_27_4 ));
    CascadeMux I__12357 (
            .O(N__57048),
            .I(\c0.n23_adj_4532_cascade_ ));
    InMux I__12356 (
            .O(N__57045),
            .I(N__57042));
    LocalMux I__12355 (
            .O(N__57042),
            .I(\c0.n31_adj_4542 ));
    CascadeMux I__12354 (
            .O(N__57039),
            .I(\c0.n38_adj_4535_cascade_ ));
    InMux I__12353 (
            .O(N__57036),
            .I(N__57033));
    LocalMux I__12352 (
            .O(N__57033),
            .I(\c0.n32_adj_4534 ));
    InMux I__12351 (
            .O(N__57030),
            .I(N__57027));
    LocalMux I__12350 (
            .O(N__57027),
            .I(N__57024));
    Odrv4 I__12349 (
            .O(N__57024),
            .I(\c0.n8_adj_4677 ));
    CascadeMux I__12348 (
            .O(N__57021),
            .I(N__57018));
    InMux I__12347 (
            .O(N__57018),
            .I(N__57011));
    InMux I__12346 (
            .O(N__57017),
            .I(N__57002));
    InMux I__12345 (
            .O(N__57016),
            .I(N__57002));
    InMux I__12344 (
            .O(N__57015),
            .I(N__57002));
    InMux I__12343 (
            .O(N__57014),
            .I(N__57002));
    LocalMux I__12342 (
            .O(N__57011),
            .I(N__56998));
    LocalMux I__12341 (
            .O(N__57002),
            .I(N__56995));
    CascadeMux I__12340 (
            .O(N__57001),
            .I(N__56991));
    Span4Mux_v I__12339 (
            .O(N__56998),
            .I(N__56988));
    Span4Mux_v I__12338 (
            .O(N__56995),
            .I(N__56985));
    InMux I__12337 (
            .O(N__56994),
            .I(N__56980));
    InMux I__12336 (
            .O(N__56991),
            .I(N__56980));
    Odrv4 I__12335 (
            .O(N__56988),
            .I(\c0.data_in_frame_25_0 ));
    Odrv4 I__12334 (
            .O(N__56985),
            .I(\c0.data_in_frame_25_0 ));
    LocalMux I__12333 (
            .O(N__56980),
            .I(\c0.data_in_frame_25_0 ));
    InMux I__12332 (
            .O(N__56973),
            .I(N__56970));
    LocalMux I__12331 (
            .O(N__56970),
            .I(N__56967));
    Odrv4 I__12330 (
            .O(N__56967),
            .I(\c0.n64_adj_4539 ));
    InMux I__12329 (
            .O(N__56964),
            .I(N__56961));
    LocalMux I__12328 (
            .O(N__56961),
            .I(N__56958));
    Odrv4 I__12327 (
            .O(N__56958),
            .I(\c0.n10_adj_4544 ));
    InMux I__12326 (
            .O(N__56955),
            .I(N__56952));
    LocalMux I__12325 (
            .O(N__56952),
            .I(\c0.n13911 ));
    CascadeMux I__12324 (
            .O(N__56949),
            .I(\c0.n23921_cascade_ ));
    InMux I__12323 (
            .O(N__56946),
            .I(N__56943));
    LocalMux I__12322 (
            .O(N__56943),
            .I(N__56940));
    Span4Mux_h I__12321 (
            .O(N__56940),
            .I(N__56937));
    Odrv4 I__12320 (
            .O(N__56937),
            .I(\c0.n21_adj_4547 ));
    InMux I__12319 (
            .O(N__56934),
            .I(N__56931));
    LocalMux I__12318 (
            .O(N__56931),
            .I(N__56928));
    Odrv12 I__12317 (
            .O(N__56928),
            .I(\c0.n23975 ));
    CascadeMux I__12316 (
            .O(N__56925),
            .I(N__56922));
    InMux I__12315 (
            .O(N__56922),
            .I(N__56919));
    LocalMux I__12314 (
            .O(N__56919),
            .I(N__56916));
    Span4Mux_h I__12313 (
            .O(N__56916),
            .I(N__56913));
    Odrv4 I__12312 (
            .O(N__56913),
            .I(\c0.n32_adj_4533 ));
    InMux I__12311 (
            .O(N__56910),
            .I(N__56907));
    LocalMux I__12310 (
            .O(N__56907),
            .I(\c0.n74 ));
    InMux I__12309 (
            .O(N__56904),
            .I(N__56898));
    InMux I__12308 (
            .O(N__56903),
            .I(N__56898));
    LocalMux I__12307 (
            .O(N__56898),
            .I(\c0.data_in_frame_29_7 ));
    InMux I__12306 (
            .O(N__56895),
            .I(N__56890));
    InMux I__12305 (
            .O(N__56894),
            .I(N__56887));
    InMux I__12304 (
            .O(N__56893),
            .I(N__56883));
    LocalMux I__12303 (
            .O(N__56890),
            .I(N__56878));
    LocalMux I__12302 (
            .O(N__56887),
            .I(N__56878));
    InMux I__12301 (
            .O(N__56886),
            .I(N__56875));
    LocalMux I__12300 (
            .O(N__56883),
            .I(N__56872));
    Span4Mux_v I__12299 (
            .O(N__56878),
            .I(N__56869));
    LocalMux I__12298 (
            .O(N__56875),
            .I(\c0.data_in_frame_27_5 ));
    Odrv4 I__12297 (
            .O(N__56872),
            .I(\c0.data_in_frame_27_5 ));
    Odrv4 I__12296 (
            .O(N__56869),
            .I(\c0.data_in_frame_27_5 ));
    InMux I__12295 (
            .O(N__56862),
            .I(N__56859));
    LocalMux I__12294 (
            .O(N__56859),
            .I(N__56855));
    InMux I__12293 (
            .O(N__56858),
            .I(N__56850));
    Span4Mux_v I__12292 (
            .O(N__56855),
            .I(N__56847));
    InMux I__12291 (
            .O(N__56854),
            .I(N__56844));
    CascadeMux I__12290 (
            .O(N__56853),
            .I(N__56841));
    LocalMux I__12289 (
            .O(N__56850),
            .I(N__56836));
    Span4Mux_h I__12288 (
            .O(N__56847),
            .I(N__56836));
    LocalMux I__12287 (
            .O(N__56844),
            .I(N__56833));
    InMux I__12286 (
            .O(N__56841),
            .I(N__56830));
    Span4Mux_h I__12285 (
            .O(N__56836),
            .I(N__56827));
    Span4Mux_v I__12284 (
            .O(N__56833),
            .I(N__56824));
    LocalMux I__12283 (
            .O(N__56830),
            .I(\c0.data_in_frame_27_6 ));
    Odrv4 I__12282 (
            .O(N__56827),
            .I(\c0.data_in_frame_27_6 ));
    Odrv4 I__12281 (
            .O(N__56824),
            .I(\c0.data_in_frame_27_6 ));
    InMux I__12280 (
            .O(N__56817),
            .I(N__56811));
    CascadeMux I__12279 (
            .O(N__56816),
            .I(N__56808));
    InMux I__12278 (
            .O(N__56815),
            .I(N__56805));
    InMux I__12277 (
            .O(N__56814),
            .I(N__56802));
    LocalMux I__12276 (
            .O(N__56811),
            .I(N__56799));
    InMux I__12275 (
            .O(N__56808),
            .I(N__56794));
    LocalMux I__12274 (
            .O(N__56805),
            .I(N__56791));
    LocalMux I__12273 (
            .O(N__56802),
            .I(N__56788));
    Span4Mux_v I__12272 (
            .O(N__56799),
            .I(N__56785));
    InMux I__12271 (
            .O(N__56798),
            .I(N__56780));
    InMux I__12270 (
            .O(N__56797),
            .I(N__56780));
    LocalMux I__12269 (
            .O(N__56794),
            .I(N__56773));
    Span4Mux_v I__12268 (
            .O(N__56791),
            .I(N__56773));
    Span4Mux_h I__12267 (
            .O(N__56788),
            .I(N__56773));
    Odrv4 I__12266 (
            .O(N__56785),
            .I(\c0.data_in_frame_25_5 ));
    LocalMux I__12265 (
            .O(N__56780),
            .I(\c0.data_in_frame_25_5 ));
    Odrv4 I__12264 (
            .O(N__56773),
            .I(\c0.data_in_frame_25_5 ));
    InMux I__12263 (
            .O(N__56766),
            .I(N__56763));
    LocalMux I__12262 (
            .O(N__56763),
            .I(\c0.n12_adj_4466 ));
    CascadeMux I__12261 (
            .O(N__56760),
            .I(\c0.n11_adj_4474_cascade_ ));
    InMux I__12260 (
            .O(N__56757),
            .I(N__56754));
    LocalMux I__12259 (
            .O(N__56754),
            .I(N__56748));
    InMux I__12258 (
            .O(N__56753),
            .I(N__56745));
    InMux I__12257 (
            .O(N__56752),
            .I(N__56742));
    InMux I__12256 (
            .O(N__56751),
            .I(N__56739));
    Span4Mux_h I__12255 (
            .O(N__56748),
            .I(N__56733));
    LocalMux I__12254 (
            .O(N__56745),
            .I(N__56726));
    LocalMux I__12253 (
            .O(N__56742),
            .I(N__56726));
    LocalMux I__12252 (
            .O(N__56739),
            .I(N__56726));
    InMux I__12251 (
            .O(N__56738),
            .I(N__56719));
    InMux I__12250 (
            .O(N__56737),
            .I(N__56719));
    InMux I__12249 (
            .O(N__56736),
            .I(N__56719));
    Odrv4 I__12248 (
            .O(N__56733),
            .I(\c0.n21280 ));
    Odrv4 I__12247 (
            .O(N__56726),
            .I(\c0.n21280 ));
    LocalMux I__12246 (
            .O(N__56719),
            .I(\c0.n21280 ));
    CascadeMux I__12245 (
            .O(N__56712),
            .I(N__56709));
    InMux I__12244 (
            .O(N__56709),
            .I(N__56706));
    LocalMux I__12243 (
            .O(N__56706),
            .I(N__56702));
    InMux I__12242 (
            .O(N__56705),
            .I(N__56699));
    Span4Mux_v I__12241 (
            .O(N__56702),
            .I(N__56696));
    LocalMux I__12240 (
            .O(N__56699),
            .I(\c0.data_in_frame_29_2 ));
    Odrv4 I__12239 (
            .O(N__56696),
            .I(\c0.data_in_frame_29_2 ));
    InMux I__12238 (
            .O(N__56691),
            .I(N__56688));
    LocalMux I__12237 (
            .O(N__56688),
            .I(\c0.n25446 ));
    CascadeMux I__12236 (
            .O(N__56685),
            .I(N__56681));
    InMux I__12235 (
            .O(N__56684),
            .I(N__56678));
    InMux I__12234 (
            .O(N__56681),
            .I(N__56675));
    LocalMux I__12233 (
            .O(N__56678),
            .I(\c0.data_in_frame_29_0 ));
    LocalMux I__12232 (
            .O(N__56675),
            .I(\c0.data_in_frame_29_0 ));
    InMux I__12231 (
            .O(N__56670),
            .I(N__56666));
    InMux I__12230 (
            .O(N__56669),
            .I(N__56663));
    LocalMux I__12229 (
            .O(N__56666),
            .I(N__56658));
    LocalMux I__12228 (
            .O(N__56663),
            .I(N__56658));
    Odrv4 I__12227 (
            .O(N__56658),
            .I(\c0.n10874 ));
    CascadeMux I__12226 (
            .O(N__56655),
            .I(\c0.n43_adj_4463_cascade_ ));
    InMux I__12225 (
            .O(N__56652),
            .I(N__56642));
    InMux I__12224 (
            .O(N__56651),
            .I(N__56642));
    InMux I__12223 (
            .O(N__56650),
            .I(N__56642));
    CascadeMux I__12222 (
            .O(N__56649),
            .I(N__56639));
    LocalMux I__12221 (
            .O(N__56642),
            .I(N__56636));
    InMux I__12220 (
            .O(N__56639),
            .I(N__56633));
    Span4Mux_v I__12219 (
            .O(N__56636),
            .I(N__56629));
    LocalMux I__12218 (
            .O(N__56633),
            .I(N__56626));
    InMux I__12217 (
            .O(N__56632),
            .I(N__56623));
    Span4Mux_h I__12216 (
            .O(N__56629),
            .I(N__56620));
    Span4Mux_v I__12215 (
            .O(N__56626),
            .I(N__56617));
    LocalMux I__12214 (
            .O(N__56623),
            .I(\c0.n21389 ));
    Odrv4 I__12213 (
            .O(N__56620),
            .I(\c0.n21389 ));
    Odrv4 I__12212 (
            .O(N__56617),
            .I(\c0.n21389 ));
    InMux I__12211 (
            .O(N__56610),
            .I(N__56607));
    LocalMux I__12210 (
            .O(N__56607),
            .I(\c0.n9_adj_4521 ));
    InMux I__12209 (
            .O(N__56604),
            .I(N__56601));
    LocalMux I__12208 (
            .O(N__56601),
            .I(\c0.n20_adj_4596 ));
    CascadeMux I__12207 (
            .O(N__56598),
            .I(\c0.n23733_cascade_ ));
    InMux I__12206 (
            .O(N__56595),
            .I(N__56589));
    InMux I__12205 (
            .O(N__56594),
            .I(N__56589));
    LocalMux I__12204 (
            .O(N__56589),
            .I(N__56585));
    InMux I__12203 (
            .O(N__56588),
            .I(N__56582));
    Span4Mux_v I__12202 (
            .O(N__56585),
            .I(N__56579));
    LocalMux I__12201 (
            .O(N__56582),
            .I(\c0.data_in_frame_26_0 ));
    Odrv4 I__12200 (
            .O(N__56579),
            .I(\c0.data_in_frame_26_0 ));
    CascadeMux I__12199 (
            .O(N__56574),
            .I(N__56569));
    InMux I__12198 (
            .O(N__56573),
            .I(N__56564));
    InMux I__12197 (
            .O(N__56572),
            .I(N__56564));
    InMux I__12196 (
            .O(N__56569),
            .I(N__56561));
    LocalMux I__12195 (
            .O(N__56564),
            .I(N__56557));
    LocalMux I__12194 (
            .O(N__56561),
            .I(N__56554));
    CascadeMux I__12193 (
            .O(N__56560),
            .I(N__56551));
    Span4Mux_v I__12192 (
            .O(N__56557),
            .I(N__56548));
    Span4Mux_h I__12191 (
            .O(N__56554),
            .I(N__56545));
    InMux I__12190 (
            .O(N__56551),
            .I(N__56542));
    Span4Mux_h I__12189 (
            .O(N__56548),
            .I(N__56539));
    Span4Mux_v I__12188 (
            .O(N__56545),
            .I(N__56536));
    LocalMux I__12187 (
            .O(N__56542),
            .I(\c0.data_in_frame_27_7 ));
    Odrv4 I__12186 (
            .O(N__56539),
            .I(\c0.data_in_frame_27_7 ));
    Odrv4 I__12185 (
            .O(N__56536),
            .I(\c0.data_in_frame_27_7 ));
    CascadeMux I__12184 (
            .O(N__56529),
            .I(\c0.n20314_cascade_ ));
    InMux I__12183 (
            .O(N__56526),
            .I(N__56523));
    LocalMux I__12182 (
            .O(N__56523),
            .I(N__56519));
    InMux I__12181 (
            .O(N__56522),
            .I(N__56516));
    Span4Mux_v I__12180 (
            .O(N__56519),
            .I(N__56512));
    LocalMux I__12179 (
            .O(N__56516),
            .I(N__56509));
    InMux I__12178 (
            .O(N__56515),
            .I(N__56506));
    Odrv4 I__12177 (
            .O(N__56512),
            .I(\c0.n21325 ));
    Odrv12 I__12176 (
            .O(N__56509),
            .I(\c0.n21325 ));
    LocalMux I__12175 (
            .O(N__56506),
            .I(\c0.n21325 ));
    InMux I__12174 (
            .O(N__56499),
            .I(N__56496));
    LocalMux I__12173 (
            .O(N__56496),
            .I(\c0.n20314 ));
    InMux I__12172 (
            .O(N__56493),
            .I(N__56490));
    LocalMux I__12171 (
            .O(N__56490),
            .I(\c0.n22_adj_4597 ));
    InMux I__12170 (
            .O(N__56487),
            .I(N__56484));
    LocalMux I__12169 (
            .O(N__56484),
            .I(N__56476));
    InMux I__12168 (
            .O(N__56483),
            .I(N__56471));
    InMux I__12167 (
            .O(N__56482),
            .I(N__56471));
    InMux I__12166 (
            .O(N__56481),
            .I(N__56468));
    InMux I__12165 (
            .O(N__56480),
            .I(N__56465));
    CascadeMux I__12164 (
            .O(N__56479),
            .I(N__56462));
    Span4Mux_h I__12163 (
            .O(N__56476),
            .I(N__56456));
    LocalMux I__12162 (
            .O(N__56471),
            .I(N__56456));
    LocalMux I__12161 (
            .O(N__56468),
            .I(N__56453));
    LocalMux I__12160 (
            .O(N__56465),
            .I(N__56450));
    InMux I__12159 (
            .O(N__56462),
            .I(N__56445));
    InMux I__12158 (
            .O(N__56461),
            .I(N__56445));
    Span4Mux_h I__12157 (
            .O(N__56456),
            .I(N__56438));
    Span4Mux_v I__12156 (
            .O(N__56453),
            .I(N__56438));
    Span4Mux_v I__12155 (
            .O(N__56450),
            .I(N__56438));
    LocalMux I__12154 (
            .O(N__56445),
            .I(N__56435));
    Span4Mux_h I__12153 (
            .O(N__56438),
            .I(N__56432));
    Odrv4 I__12152 (
            .O(N__56435),
            .I(\c0.n12_adj_4671 ));
    Odrv4 I__12151 (
            .O(N__56432),
            .I(\c0.n12_adj_4671 ));
    InMux I__12150 (
            .O(N__56427),
            .I(N__56424));
    LocalMux I__12149 (
            .O(N__56424),
            .I(N__56421));
    Odrv12 I__12148 (
            .O(N__56421),
            .I(\c0.n22_adj_4350 ));
    CascadeMux I__12147 (
            .O(N__56418),
            .I(\c0.n22_adj_4350_cascade_ ));
    InMux I__12146 (
            .O(N__56415),
            .I(N__56412));
    LocalMux I__12145 (
            .O(N__56412),
            .I(N__56408));
    CascadeMux I__12144 (
            .O(N__56411),
            .I(N__56403));
    Span4Mux_h I__12143 (
            .O(N__56408),
            .I(N__56400));
    CascadeMux I__12142 (
            .O(N__56407),
            .I(N__56397));
    InMux I__12141 (
            .O(N__56406),
            .I(N__56393));
    InMux I__12140 (
            .O(N__56403),
            .I(N__56390));
    Span4Mux_v I__12139 (
            .O(N__56400),
            .I(N__56387));
    InMux I__12138 (
            .O(N__56397),
            .I(N__56382));
    InMux I__12137 (
            .O(N__56396),
            .I(N__56382));
    LocalMux I__12136 (
            .O(N__56393),
            .I(\c0.data_in_frame_20_6 ));
    LocalMux I__12135 (
            .O(N__56390),
            .I(\c0.data_in_frame_20_6 ));
    Odrv4 I__12134 (
            .O(N__56387),
            .I(\c0.data_in_frame_20_6 ));
    LocalMux I__12133 (
            .O(N__56382),
            .I(\c0.data_in_frame_20_6 ));
    InMux I__12132 (
            .O(N__56373),
            .I(N__56366));
    InMux I__12131 (
            .O(N__56372),
            .I(N__56361));
    InMux I__12130 (
            .O(N__56371),
            .I(N__56361));
    CascadeMux I__12129 (
            .O(N__56370),
            .I(N__56358));
    InMux I__12128 (
            .O(N__56369),
            .I(N__56355));
    LocalMux I__12127 (
            .O(N__56366),
            .I(N__56351));
    LocalMux I__12126 (
            .O(N__56361),
            .I(N__56348));
    InMux I__12125 (
            .O(N__56358),
            .I(N__56345));
    LocalMux I__12124 (
            .O(N__56355),
            .I(N__56342));
    InMux I__12123 (
            .O(N__56354),
            .I(N__56339));
    Span4Mux_h I__12122 (
            .O(N__56351),
            .I(N__56334));
    Span4Mux_v I__12121 (
            .O(N__56348),
            .I(N__56334));
    LocalMux I__12120 (
            .O(N__56345),
            .I(\c0.data_in_frame_20_7 ));
    Odrv12 I__12119 (
            .O(N__56342),
            .I(\c0.data_in_frame_20_7 ));
    LocalMux I__12118 (
            .O(N__56339),
            .I(\c0.data_in_frame_20_7 ));
    Odrv4 I__12117 (
            .O(N__56334),
            .I(\c0.data_in_frame_20_7 ));
    InMux I__12116 (
            .O(N__56325),
            .I(N__56317));
    InMux I__12115 (
            .O(N__56324),
            .I(N__56317));
    InMux I__12114 (
            .O(N__56323),
            .I(N__56312));
    InMux I__12113 (
            .O(N__56322),
            .I(N__56312));
    LocalMux I__12112 (
            .O(N__56317),
            .I(N__56309));
    LocalMux I__12111 (
            .O(N__56312),
            .I(N__56306));
    Span4Mux_v I__12110 (
            .O(N__56309),
            .I(N__56303));
    Odrv4 I__12109 (
            .O(N__56306),
            .I(\c0.n21_adj_4225 ));
    Odrv4 I__12108 (
            .O(N__56303),
            .I(\c0.n21_adj_4225 ));
    CascadeMux I__12107 (
            .O(N__56298),
            .I(N__56295));
    InMux I__12106 (
            .O(N__56295),
            .I(N__56292));
    LocalMux I__12105 (
            .O(N__56292),
            .I(N__56289));
    Span4Mux_h I__12104 (
            .O(N__56289),
            .I(N__56286));
    Span4Mux_h I__12103 (
            .O(N__56286),
            .I(N__56283));
    Odrv4 I__12102 (
            .O(N__56283),
            .I(\c0.n22227 ));
    InMux I__12101 (
            .O(N__56280),
            .I(N__56277));
    LocalMux I__12100 (
            .O(N__56277),
            .I(N__56273));
    InMux I__12099 (
            .O(N__56276),
            .I(N__56269));
    Span4Mux_h I__12098 (
            .O(N__56273),
            .I(N__56265));
    InMux I__12097 (
            .O(N__56272),
            .I(N__56262));
    LocalMux I__12096 (
            .O(N__56269),
            .I(N__56259));
    InMux I__12095 (
            .O(N__56268),
            .I(N__56256));
    Odrv4 I__12094 (
            .O(N__56265),
            .I(\c0.n23863 ));
    LocalMux I__12093 (
            .O(N__56262),
            .I(\c0.n23863 ));
    Odrv4 I__12092 (
            .O(N__56259),
            .I(\c0.n23863 ));
    LocalMux I__12091 (
            .O(N__56256),
            .I(\c0.n23863 ));
    InMux I__12090 (
            .O(N__56247),
            .I(N__56244));
    LocalMux I__12089 (
            .O(N__56244),
            .I(\c0.n160 ));
    InMux I__12088 (
            .O(N__56241),
            .I(N__56236));
    InMux I__12087 (
            .O(N__56240),
            .I(N__56233));
    InMux I__12086 (
            .O(N__56239),
            .I(N__56230));
    LocalMux I__12085 (
            .O(N__56236),
            .I(N__56227));
    LocalMux I__12084 (
            .O(N__56233),
            .I(N__56224));
    LocalMux I__12083 (
            .O(N__56230),
            .I(N__56220));
    Span4Mux_h I__12082 (
            .O(N__56227),
            .I(N__56217));
    Span4Mux_h I__12081 (
            .O(N__56224),
            .I(N__56214));
    InMux I__12080 (
            .O(N__56223),
            .I(N__56211));
    Span4Mux_v I__12079 (
            .O(N__56220),
            .I(N__56208));
    Span4Mux_v I__12078 (
            .O(N__56217),
            .I(N__56203));
    Span4Mux_v I__12077 (
            .O(N__56214),
            .I(N__56203));
    LocalMux I__12076 (
            .O(N__56211),
            .I(\c0.n12989 ));
    Odrv4 I__12075 (
            .O(N__56208),
            .I(\c0.n12989 ));
    Odrv4 I__12074 (
            .O(N__56203),
            .I(\c0.n12989 ));
    CascadeMux I__12073 (
            .O(N__56196),
            .I(\c0.n22104_cascade_ ));
    InMux I__12072 (
            .O(N__56193),
            .I(N__56189));
    InMux I__12071 (
            .O(N__56192),
            .I(N__56186));
    LocalMux I__12070 (
            .O(N__56189),
            .I(N__56182));
    LocalMux I__12069 (
            .O(N__56186),
            .I(N__56179));
    InMux I__12068 (
            .O(N__56185),
            .I(N__56176));
    Span4Mux_v I__12067 (
            .O(N__56182),
            .I(N__56171));
    Span4Mux_h I__12066 (
            .O(N__56179),
            .I(N__56171));
    LocalMux I__12065 (
            .O(N__56176),
            .I(\c0.data_in_frame_19_4 ));
    Odrv4 I__12064 (
            .O(N__56171),
            .I(\c0.data_in_frame_19_4 ));
    CascadeMux I__12063 (
            .O(N__56166),
            .I(\c0.n22347_cascade_ ));
    InMux I__12062 (
            .O(N__56163),
            .I(N__56160));
    LocalMux I__12061 (
            .O(N__56160),
            .I(N__56156));
    InMux I__12060 (
            .O(N__56159),
            .I(N__56153));
    Odrv4 I__12059 (
            .O(N__56156),
            .I(\c0.n24520 ));
    LocalMux I__12058 (
            .O(N__56153),
            .I(\c0.n24520 ));
    InMux I__12057 (
            .O(N__56148),
            .I(N__56144));
    InMux I__12056 (
            .O(N__56147),
            .I(N__56140));
    LocalMux I__12055 (
            .O(N__56144),
            .I(N__56136));
    InMux I__12054 (
            .O(N__56143),
            .I(N__56133));
    LocalMux I__12053 (
            .O(N__56140),
            .I(N__56130));
    InMux I__12052 (
            .O(N__56139),
            .I(N__56127));
    Span4Mux_v I__12051 (
            .O(N__56136),
            .I(N__56124));
    LocalMux I__12050 (
            .O(N__56133),
            .I(N__56119));
    Span4Mux_v I__12049 (
            .O(N__56130),
            .I(N__56119));
    LocalMux I__12048 (
            .O(N__56127),
            .I(\c0.data_in_frame_20_5 ));
    Odrv4 I__12047 (
            .O(N__56124),
            .I(\c0.data_in_frame_20_5 ));
    Odrv4 I__12046 (
            .O(N__56119),
            .I(\c0.data_in_frame_20_5 ));
    InMux I__12045 (
            .O(N__56112),
            .I(N__56109));
    LocalMux I__12044 (
            .O(N__56109),
            .I(N__56106));
    Odrv4 I__12043 (
            .O(N__56106),
            .I(\c0.n33 ));
    CascadeMux I__12042 (
            .O(N__56103),
            .I(\c0.n34_adj_4600_cascade_ ));
    InMux I__12041 (
            .O(N__56100),
            .I(N__56097));
    LocalMux I__12040 (
            .O(N__56097),
            .I(N__56094));
    Span4Mux_v I__12039 (
            .O(N__56094),
            .I(N__56091));
    Odrv4 I__12038 (
            .O(N__56091),
            .I(\c0.n38_adj_4573 ));
    CascadeMux I__12037 (
            .O(N__56088),
            .I(\c0.n24333_cascade_ ));
    InMux I__12036 (
            .O(N__56085),
            .I(N__56079));
    InMux I__12035 (
            .O(N__56084),
            .I(N__56079));
    LocalMux I__12034 (
            .O(N__56079),
            .I(N__56076));
    Odrv4 I__12033 (
            .O(N__56076),
            .I(\c0.n23661 ));
    CascadeMux I__12032 (
            .O(N__56073),
            .I(N__56069));
    CascadeMux I__12031 (
            .O(N__56072),
            .I(N__56066));
    InMux I__12030 (
            .O(N__56069),
            .I(N__56063));
    InMux I__12029 (
            .O(N__56066),
            .I(N__56060));
    LocalMux I__12028 (
            .O(N__56063),
            .I(N__56057));
    LocalMux I__12027 (
            .O(N__56060),
            .I(N__56051));
    Span4Mux_h I__12026 (
            .O(N__56057),
            .I(N__56051));
    InMux I__12025 (
            .O(N__56056),
            .I(N__56048));
    Odrv4 I__12024 (
            .O(N__56051),
            .I(\c0.data_in_frame_18_5 ));
    LocalMux I__12023 (
            .O(N__56048),
            .I(\c0.data_in_frame_18_5 ));
    InMux I__12022 (
            .O(N__56043),
            .I(N__56040));
    LocalMux I__12021 (
            .O(N__56040),
            .I(N__56035));
    InMux I__12020 (
            .O(N__56039),
            .I(N__56030));
    InMux I__12019 (
            .O(N__56038),
            .I(N__56030));
    Span4Mux_h I__12018 (
            .O(N__56035),
            .I(N__56027));
    LocalMux I__12017 (
            .O(N__56030),
            .I(\c0.data_in_frame_16_3 ));
    Odrv4 I__12016 (
            .O(N__56027),
            .I(\c0.data_in_frame_16_3 ));
    InMux I__12015 (
            .O(N__56022),
            .I(N__56019));
    LocalMux I__12014 (
            .O(N__56019),
            .I(N__56016));
    Odrv12 I__12013 (
            .O(N__56016),
            .I(\c0.n155 ));
    InMux I__12012 (
            .O(N__56013),
            .I(N__56010));
    LocalMux I__12011 (
            .O(N__56010),
            .I(N__56006));
    CascadeMux I__12010 (
            .O(N__56009),
            .I(N__56002));
    Span4Mux_v I__12009 (
            .O(N__56006),
            .I(N__55999));
    InMux I__12008 (
            .O(N__56005),
            .I(N__55994));
    InMux I__12007 (
            .O(N__56002),
            .I(N__55994));
    Span4Mux_v I__12006 (
            .O(N__55999),
            .I(N__55991));
    LocalMux I__12005 (
            .O(N__55994),
            .I(N__55988));
    Odrv4 I__12004 (
            .O(N__55991),
            .I(\c0.n5_adj_4311 ));
    Odrv4 I__12003 (
            .O(N__55988),
            .I(\c0.n5_adj_4311 ));
    CascadeMux I__12002 (
            .O(N__55983),
            .I(\c0.n5_adj_4311_cascade_ ));
    InMux I__12001 (
            .O(N__55980),
            .I(N__55977));
    LocalMux I__12000 (
            .O(N__55977),
            .I(N__55973));
    InMux I__11999 (
            .O(N__55976),
            .I(N__55969));
    Span4Mux_h I__11998 (
            .O(N__55973),
            .I(N__55966));
    InMux I__11997 (
            .O(N__55972),
            .I(N__55962));
    LocalMux I__11996 (
            .O(N__55969),
            .I(N__55959));
    Span4Mux_v I__11995 (
            .O(N__55966),
            .I(N__55956));
    InMux I__11994 (
            .O(N__55965),
            .I(N__55953));
    LocalMux I__11993 (
            .O(N__55962),
            .I(\c0.data_in_frame_10_3 ));
    Odrv4 I__11992 (
            .O(N__55959),
            .I(\c0.data_in_frame_10_3 ));
    Odrv4 I__11991 (
            .O(N__55956),
            .I(\c0.data_in_frame_10_3 ));
    LocalMux I__11990 (
            .O(N__55953),
            .I(\c0.data_in_frame_10_3 ));
    InMux I__11989 (
            .O(N__55944),
            .I(N__55938));
    InMux I__11988 (
            .O(N__55943),
            .I(N__55938));
    LocalMux I__11987 (
            .O(N__55938),
            .I(N__55935));
    Odrv12 I__11986 (
            .O(N__55935),
            .I(\c0.n23677 ));
    CascadeMux I__11985 (
            .O(N__55932),
            .I(N__55928));
    InMux I__11984 (
            .O(N__55931),
            .I(N__55923));
    InMux I__11983 (
            .O(N__55928),
            .I(N__55923));
    LocalMux I__11982 (
            .O(N__55923),
            .I(N__55920));
    Span4Mux_h I__11981 (
            .O(N__55920),
            .I(N__55916));
    InMux I__11980 (
            .O(N__55919),
            .I(N__55913));
    Span4Mux_v I__11979 (
            .O(N__55916),
            .I(N__55910));
    LocalMux I__11978 (
            .O(N__55913),
            .I(data_in_frame_14_4));
    Odrv4 I__11977 (
            .O(N__55910),
            .I(data_in_frame_14_4));
    CascadeMux I__11976 (
            .O(N__55905),
            .I(N__55902));
    InMux I__11975 (
            .O(N__55902),
            .I(N__55889));
    InMux I__11974 (
            .O(N__55901),
            .I(N__55889));
    InMux I__11973 (
            .O(N__55900),
            .I(N__55889));
    InMux I__11972 (
            .O(N__55899),
            .I(N__55889));
    CascadeMux I__11971 (
            .O(N__55898),
            .I(N__55886));
    LocalMux I__11970 (
            .O(N__55889),
            .I(N__55883));
    InMux I__11969 (
            .O(N__55886),
            .I(N__55879));
    Span4Mux_h I__11968 (
            .O(N__55883),
            .I(N__55876));
    InMux I__11967 (
            .O(N__55882),
            .I(N__55873));
    LocalMux I__11966 (
            .O(N__55879),
            .I(\c0.data_in_frame_8_2 ));
    Odrv4 I__11965 (
            .O(N__55876),
            .I(\c0.data_in_frame_8_2 ));
    LocalMux I__11964 (
            .O(N__55873),
            .I(\c0.data_in_frame_8_2 ));
    CascadeMux I__11963 (
            .O(N__55866),
            .I(\c0.n120_cascade_ ));
    InMux I__11962 (
            .O(N__55863),
            .I(N__55860));
    LocalMux I__11961 (
            .O(N__55860),
            .I(N__55857));
    Span4Mux_v I__11960 (
            .O(N__55857),
            .I(N__55854));
    Odrv4 I__11959 (
            .O(N__55854),
            .I(\c0.n142 ));
    CascadeMux I__11958 (
            .O(N__55851),
            .I(\c0.n152_cascade_ ));
    InMux I__11957 (
            .O(N__55848),
            .I(N__55845));
    LocalMux I__11956 (
            .O(N__55845),
            .I(N__55842));
    Odrv4 I__11955 (
            .O(N__55842),
            .I(\c0.n158 ));
    InMux I__11954 (
            .O(N__55839),
            .I(N__55835));
    InMux I__11953 (
            .O(N__55838),
            .I(N__55832));
    LocalMux I__11952 (
            .O(N__55835),
            .I(N__55827));
    LocalMux I__11951 (
            .O(N__55832),
            .I(N__55827));
    Odrv12 I__11950 (
            .O(N__55827),
            .I(\c0.n22472 ));
    InMux I__11949 (
            .O(N__55824),
            .I(N__55820));
    CascadeMux I__11948 (
            .O(N__55823),
            .I(N__55817));
    LocalMux I__11947 (
            .O(N__55820),
            .I(N__55814));
    InMux I__11946 (
            .O(N__55817),
            .I(N__55811));
    Span4Mux_h I__11945 (
            .O(N__55814),
            .I(N__55808));
    LocalMux I__11944 (
            .O(N__55811),
            .I(data_in_frame_14_3));
    Odrv4 I__11943 (
            .O(N__55808),
            .I(data_in_frame_14_3));
    CascadeMux I__11942 (
            .O(N__55803),
            .I(\c0.n30_adj_4571_cascade_ ));
    InMux I__11941 (
            .O(N__55800),
            .I(N__55790));
    InMux I__11940 (
            .O(N__55799),
            .I(N__55790));
    InMux I__11939 (
            .O(N__55798),
            .I(N__55790));
    InMux I__11938 (
            .O(N__55797),
            .I(N__55787));
    LocalMux I__11937 (
            .O(N__55790),
            .I(N__55782));
    LocalMux I__11936 (
            .O(N__55787),
            .I(N__55782));
    Odrv4 I__11935 (
            .O(N__55782),
            .I(\c0.data_in_frame_4_1 ));
    CascadeMux I__11934 (
            .O(N__55779),
            .I(N__55776));
    InMux I__11933 (
            .O(N__55776),
            .I(N__55770));
    InMux I__11932 (
            .O(N__55775),
            .I(N__55770));
    LocalMux I__11931 (
            .O(N__55770),
            .I(\c0.data_in_frame_10_4 ));
    InMux I__11930 (
            .O(N__55767),
            .I(N__55761));
    InMux I__11929 (
            .O(N__55766),
            .I(N__55761));
    LocalMux I__11928 (
            .O(N__55761),
            .I(N__55757));
    InMux I__11927 (
            .O(N__55760),
            .I(N__55754));
    Span4Mux_h I__11926 (
            .O(N__55757),
            .I(N__55751));
    LocalMux I__11925 (
            .O(N__55754),
            .I(\c0.n22455 ));
    Odrv4 I__11924 (
            .O(N__55751),
            .I(\c0.n22455 ));
    CascadeMux I__11923 (
            .O(N__55746),
            .I(N__55743));
    InMux I__11922 (
            .O(N__55743),
            .I(N__55737));
    CascadeMux I__11921 (
            .O(N__55742),
            .I(N__55734));
    InMux I__11920 (
            .O(N__55741),
            .I(N__55731));
    InMux I__11919 (
            .O(N__55740),
            .I(N__55728));
    LocalMux I__11918 (
            .O(N__55737),
            .I(N__55724));
    InMux I__11917 (
            .O(N__55734),
            .I(N__55721));
    LocalMux I__11916 (
            .O(N__55731),
            .I(N__55718));
    LocalMux I__11915 (
            .O(N__55728),
            .I(N__55715));
    InMux I__11914 (
            .O(N__55727),
            .I(N__55712));
    Span4Mux_h I__11913 (
            .O(N__55724),
            .I(N__55709));
    LocalMux I__11912 (
            .O(N__55721),
            .I(N__55704));
    Span4Mux_v I__11911 (
            .O(N__55718),
            .I(N__55704));
    Span4Mux_h I__11910 (
            .O(N__55715),
            .I(N__55701));
    LocalMux I__11909 (
            .O(N__55712),
            .I(N__55698));
    Span4Mux_v I__11908 (
            .O(N__55709),
            .I(N__55695));
    Odrv4 I__11907 (
            .O(N__55704),
            .I(\c0.data_in_frame_12_5 ));
    Odrv4 I__11906 (
            .O(N__55701),
            .I(\c0.data_in_frame_12_5 ));
    Odrv4 I__11905 (
            .O(N__55698),
            .I(\c0.data_in_frame_12_5 ));
    Odrv4 I__11904 (
            .O(N__55695),
            .I(\c0.data_in_frame_12_5 ));
    InMux I__11903 (
            .O(N__55686),
            .I(N__55683));
    LocalMux I__11902 (
            .O(N__55683),
            .I(N__55679));
    CascadeMux I__11901 (
            .O(N__55682),
            .I(N__55676));
    Span4Mux_h I__11900 (
            .O(N__55679),
            .I(N__55673));
    InMux I__11899 (
            .O(N__55676),
            .I(N__55670));
    Sp12to4 I__11898 (
            .O(N__55673),
            .I(N__55665));
    LocalMux I__11897 (
            .O(N__55670),
            .I(N__55665));
    Span12Mux_v I__11896 (
            .O(N__55665),
            .I(N__55661));
    InMux I__11895 (
            .O(N__55664),
            .I(N__55658));
    Odrv12 I__11894 (
            .O(N__55661),
            .I(\c0.n42 ));
    LocalMux I__11893 (
            .O(N__55658),
            .I(\c0.n42 ));
    InMux I__11892 (
            .O(N__55653),
            .I(N__55650));
    LocalMux I__11891 (
            .O(N__55650),
            .I(N__55647));
    Odrv4 I__11890 (
            .O(N__55647),
            .I(\c0.n58 ));
    InMux I__11889 (
            .O(N__55644),
            .I(N__55641));
    LocalMux I__11888 (
            .O(N__55641),
            .I(N__55638));
    Odrv4 I__11887 (
            .O(N__55638),
            .I(\c0.n127 ));
    CascadeMux I__11886 (
            .O(N__55635),
            .I(\c0.n41_adj_4452_cascade_ ));
    InMux I__11885 (
            .O(N__55632),
            .I(N__55627));
    InMux I__11884 (
            .O(N__55631),
            .I(N__55624));
    InMux I__11883 (
            .O(N__55630),
            .I(N__55621));
    LocalMux I__11882 (
            .O(N__55627),
            .I(N__55618));
    LocalMux I__11881 (
            .O(N__55624),
            .I(N__55615));
    LocalMux I__11880 (
            .O(N__55621),
            .I(N__55612));
    Span4Mux_h I__11879 (
            .O(N__55618),
            .I(N__55604));
    Span4Mux_v I__11878 (
            .O(N__55615),
            .I(N__55604));
    Span4Mux_v I__11877 (
            .O(N__55612),
            .I(N__55604));
    InMux I__11876 (
            .O(N__55611),
            .I(N__55601));
    Span4Mux_h I__11875 (
            .O(N__55604),
            .I(N__55598));
    LocalMux I__11874 (
            .O(N__55601),
            .I(\c0.data_in_frame_11_7 ));
    Odrv4 I__11873 (
            .O(N__55598),
            .I(\c0.data_in_frame_11_7 ));
    InMux I__11872 (
            .O(N__55593),
            .I(N__55590));
    LocalMux I__11871 (
            .O(N__55590),
            .I(\c0.n39_adj_4453 ));
    InMux I__11870 (
            .O(N__55587),
            .I(N__55584));
    LocalMux I__11869 (
            .O(N__55584),
            .I(\c0.n40_adj_4451 ));
    CascadeMux I__11868 (
            .O(N__55581),
            .I(N__55578));
    InMux I__11867 (
            .O(N__55578),
            .I(N__55575));
    LocalMux I__11866 (
            .O(N__55575),
            .I(N__55572));
    Span4Mux_h I__11865 (
            .O(N__55572),
            .I(N__55569));
    Odrv4 I__11864 (
            .O(N__55569),
            .I(\c0.n14016 ));
    InMux I__11863 (
            .O(N__55566),
            .I(N__55561));
    InMux I__11862 (
            .O(N__55565),
            .I(N__55558));
    CascadeMux I__11861 (
            .O(N__55564),
            .I(N__55555));
    LocalMux I__11860 (
            .O(N__55561),
            .I(N__55552));
    LocalMux I__11859 (
            .O(N__55558),
            .I(N__55549));
    InMux I__11858 (
            .O(N__55555),
            .I(N__55546));
    Span4Mux_v I__11857 (
            .O(N__55552),
            .I(N__55543));
    Span4Mux_v I__11856 (
            .O(N__55549),
            .I(N__55538));
    LocalMux I__11855 (
            .O(N__55546),
            .I(N__55538));
    Odrv4 I__11854 (
            .O(N__55543),
            .I(\c0.n13223 ));
    Odrv4 I__11853 (
            .O(N__55538),
            .I(\c0.n13223 ));
    InMux I__11852 (
            .O(N__55533),
            .I(N__55530));
    LocalMux I__11851 (
            .O(N__55530),
            .I(N__55527));
    Odrv4 I__11850 (
            .O(N__55527),
            .I(\c0.n16_adj_4608 ));
    InMux I__11849 (
            .O(N__55524),
            .I(N__55520));
    InMux I__11848 (
            .O(N__55523),
            .I(N__55517));
    LocalMux I__11847 (
            .O(N__55520),
            .I(N__55514));
    LocalMux I__11846 (
            .O(N__55517),
            .I(N__55509));
    Span4Mux_h I__11845 (
            .O(N__55514),
            .I(N__55505));
    InMux I__11844 (
            .O(N__55513),
            .I(N__55500));
    InMux I__11843 (
            .O(N__55512),
            .I(N__55500));
    Span12Mux_v I__11842 (
            .O(N__55509),
            .I(N__55497));
    InMux I__11841 (
            .O(N__55508),
            .I(N__55494));
    Sp12to4 I__11840 (
            .O(N__55505),
            .I(N__55489));
    LocalMux I__11839 (
            .O(N__55500),
            .I(N__55489));
    Odrv12 I__11838 (
            .O(N__55497),
            .I(\c0.n21 ));
    LocalMux I__11837 (
            .O(N__55494),
            .I(\c0.n21 ));
    Odrv12 I__11836 (
            .O(N__55489),
            .I(\c0.n21 ));
    CascadeMux I__11835 (
            .O(N__55482),
            .I(N__55479));
    InMux I__11834 (
            .O(N__55479),
            .I(N__55475));
    InMux I__11833 (
            .O(N__55478),
            .I(N__55472));
    LocalMux I__11832 (
            .O(N__55475),
            .I(N__55469));
    LocalMux I__11831 (
            .O(N__55472),
            .I(N__55466));
    Span4Mux_h I__11830 (
            .O(N__55469),
            .I(N__55463));
    Span4Mux_h I__11829 (
            .O(N__55466),
            .I(N__55460));
    Odrv4 I__11828 (
            .O(N__55463),
            .I(\c0.n20 ));
    Odrv4 I__11827 (
            .O(N__55460),
            .I(\c0.n20 ));
    InMux I__11826 (
            .O(N__55455),
            .I(N__55451));
    InMux I__11825 (
            .O(N__55454),
            .I(N__55448));
    LocalMux I__11824 (
            .O(N__55451),
            .I(N__55445));
    LocalMux I__11823 (
            .O(N__55448),
            .I(N__55442));
    Span4Mux_v I__11822 (
            .O(N__55445),
            .I(N__55439));
    Odrv12 I__11821 (
            .O(N__55442),
            .I(\c0.n13_adj_4610 ));
    Odrv4 I__11820 (
            .O(N__55439),
            .I(\c0.n13_adj_4610 ));
    InMux I__11819 (
            .O(N__55434),
            .I(N__55431));
    LocalMux I__11818 (
            .O(N__55431),
            .I(N__55426));
    InMux I__11817 (
            .O(N__55430),
            .I(N__55423));
    InMux I__11816 (
            .O(N__55429),
            .I(N__55420));
    Span4Mux_h I__11815 (
            .O(N__55426),
            .I(N__55415));
    LocalMux I__11814 (
            .O(N__55423),
            .I(N__55415));
    LocalMux I__11813 (
            .O(N__55420),
            .I(data_in_frame_14_1));
    Odrv4 I__11812 (
            .O(N__55415),
            .I(data_in_frame_14_1));
    InMux I__11811 (
            .O(N__55410),
            .I(N__55407));
    LocalMux I__11810 (
            .O(N__55407),
            .I(N__55404));
    Odrv4 I__11809 (
            .O(N__55404),
            .I(\c0.n102 ));
    CascadeMux I__11808 (
            .O(N__55401),
            .I(\c0.n147_cascade_ ));
    InMux I__11807 (
            .O(N__55398),
            .I(N__55395));
    LocalMux I__11806 (
            .O(N__55395),
            .I(\c0.n134 ));
    CascadeMux I__11805 (
            .O(N__55392),
            .I(N__55389));
    InMux I__11804 (
            .O(N__55389),
            .I(N__55386));
    LocalMux I__11803 (
            .O(N__55386),
            .I(\c0.n131 ));
    CascadeMux I__11802 (
            .O(N__55383),
            .I(N__55380));
    InMux I__11801 (
            .O(N__55380),
            .I(N__55377));
    LocalMux I__11800 (
            .O(N__55377),
            .I(N__55374));
    Span4Mux_h I__11799 (
            .O(N__55374),
            .I(N__55371));
    Odrv4 I__11798 (
            .O(N__55371),
            .I(\c0.n31_adj_4284 ));
    InMux I__11797 (
            .O(N__55368),
            .I(N__55365));
    LocalMux I__11796 (
            .O(N__55365),
            .I(\c0.n36_adj_4447 ));
    InMux I__11795 (
            .O(N__55362),
            .I(N__55359));
    LocalMux I__11794 (
            .O(N__55359),
            .I(N__55356));
    Span4Mux_v I__11793 (
            .O(N__55356),
            .I(N__55353));
    Odrv4 I__11792 (
            .O(N__55353),
            .I(\c0.n5_adj_4268 ));
    InMux I__11791 (
            .O(N__55350),
            .I(N__55347));
    LocalMux I__11790 (
            .O(N__55347),
            .I(N__55344));
    Span4Mux_h I__11789 (
            .O(N__55344),
            .I(N__55341));
    Odrv4 I__11788 (
            .O(N__55341),
            .I(\c0.n4_adj_4267 ));
    InMux I__11787 (
            .O(N__55338),
            .I(N__55335));
    LocalMux I__11786 (
            .O(N__55335),
            .I(\c0.n4_adj_4269 ));
    InMux I__11785 (
            .O(N__55332),
            .I(N__55326));
    InMux I__11784 (
            .O(N__55331),
            .I(N__55323));
    InMux I__11783 (
            .O(N__55330),
            .I(N__55319));
    CascadeMux I__11782 (
            .O(N__55329),
            .I(N__55316));
    LocalMux I__11781 (
            .O(N__55326),
            .I(N__55311));
    LocalMux I__11780 (
            .O(N__55323),
            .I(N__55311));
    InMux I__11779 (
            .O(N__55322),
            .I(N__55308));
    LocalMux I__11778 (
            .O(N__55319),
            .I(N__55305));
    InMux I__11777 (
            .O(N__55316),
            .I(N__55302));
    Span4Mux_v I__11776 (
            .O(N__55311),
            .I(N__55297));
    LocalMux I__11775 (
            .O(N__55308),
            .I(N__55297));
    Odrv4 I__11774 (
            .O(N__55305),
            .I(\c0.n22196 ));
    LocalMux I__11773 (
            .O(N__55302),
            .I(\c0.n22196 ));
    Odrv4 I__11772 (
            .O(N__55297),
            .I(\c0.n22196 ));
    CascadeMux I__11771 (
            .O(N__55290),
            .I(\c0.n4_adj_4269_cascade_ ));
    InMux I__11770 (
            .O(N__55287),
            .I(N__55284));
    LocalMux I__11769 (
            .O(N__55284),
            .I(\c0.n68 ));
    CascadeMux I__11768 (
            .O(N__55281),
            .I(\c0.n89_cascade_ ));
    CascadeMux I__11767 (
            .O(N__55278),
            .I(\c0.n23_cascade_ ));
    CascadeMux I__11766 (
            .O(N__55275),
            .I(N__55272));
    InMux I__11765 (
            .O(N__55272),
            .I(N__55269));
    LocalMux I__11764 (
            .O(N__55269),
            .I(N__55266));
    Span4Mux_v I__11763 (
            .O(N__55266),
            .I(N__55263));
    Span4Mux_v I__11762 (
            .O(N__55263),
            .I(N__55260));
    Odrv4 I__11761 (
            .O(N__55260),
            .I(\c0.n26 ));
    CascadeMux I__11760 (
            .O(N__55257),
            .I(\c0.n13075_cascade_ ));
    CascadeMux I__11759 (
            .O(N__55254),
            .I(\c0.n93_cascade_ ));
    InMux I__11758 (
            .O(N__55251),
            .I(N__55248));
    LocalMux I__11757 (
            .O(N__55248),
            .I(\c0.n12_adj_4299 ));
    CascadeMux I__11756 (
            .O(N__55245),
            .I(\c0.n7_adj_4300_cascade_ ));
    InMux I__11755 (
            .O(N__55242),
            .I(N__55238));
    CascadeMux I__11754 (
            .O(N__55241),
            .I(N__55235));
    LocalMux I__11753 (
            .O(N__55238),
            .I(N__55232));
    InMux I__11752 (
            .O(N__55235),
            .I(N__55229));
    Span4Mux_v I__11751 (
            .O(N__55232),
            .I(N__55226));
    LocalMux I__11750 (
            .O(N__55229),
            .I(\c0.n11_adj_4280 ));
    Odrv4 I__11749 (
            .O(N__55226),
            .I(\c0.n11_adj_4280 ));
    InMux I__11748 (
            .O(N__55221),
            .I(N__55217));
    InMux I__11747 (
            .O(N__55220),
            .I(N__55214));
    LocalMux I__11746 (
            .O(N__55217),
            .I(N__55211));
    LocalMux I__11745 (
            .O(N__55214),
            .I(N__55208));
    Span4Mux_h I__11744 (
            .O(N__55211),
            .I(N__55203));
    Span4Mux_h I__11743 (
            .O(N__55208),
            .I(N__55200));
    InMux I__11742 (
            .O(N__55207),
            .I(N__55195));
    InMux I__11741 (
            .O(N__55206),
            .I(N__55195));
    Odrv4 I__11740 (
            .O(N__55203),
            .I(\c0.n23251 ));
    Odrv4 I__11739 (
            .O(N__55200),
            .I(\c0.n23251 ));
    LocalMux I__11738 (
            .O(N__55195),
            .I(\c0.n23251 ));
    InMux I__11737 (
            .O(N__55188),
            .I(N__55179));
    InMux I__11736 (
            .O(N__55187),
            .I(N__55179));
    InMux I__11735 (
            .O(N__55186),
            .I(N__55174));
    InMux I__11734 (
            .O(N__55185),
            .I(N__55174));
    InMux I__11733 (
            .O(N__55184),
            .I(N__55171));
    LocalMux I__11732 (
            .O(N__55179),
            .I(N__55168));
    LocalMux I__11731 (
            .O(N__55174),
            .I(N__55165));
    LocalMux I__11730 (
            .O(N__55171),
            .I(N__55162));
    Span4Mux_h I__11729 (
            .O(N__55168),
            .I(N__55157));
    Span4Mux_v I__11728 (
            .O(N__55165),
            .I(N__55157));
    Odrv4 I__11727 (
            .O(N__55162),
            .I(\c0.n23305 ));
    Odrv4 I__11726 (
            .O(N__55157),
            .I(\c0.n23305 ));
    CascadeMux I__11725 (
            .O(N__55152),
            .I(\c0.n23251_cascade_ ));
    InMux I__11724 (
            .O(N__55149),
            .I(N__55146));
    LocalMux I__11723 (
            .O(N__55146),
            .I(N__55143));
    Span4Mux_v I__11722 (
            .O(N__55143),
            .I(N__55140));
    Odrv4 I__11721 (
            .O(N__55140),
            .I(\c0.n23574 ));
    CascadeMux I__11720 (
            .O(N__55137),
            .I(\c0.n7_adj_4282_cascade_ ));
    InMux I__11719 (
            .O(N__55134),
            .I(N__55128));
    InMux I__11718 (
            .O(N__55133),
            .I(N__55128));
    LocalMux I__11717 (
            .O(N__55128),
            .I(\c0.n10_adj_4283 ));
    InMux I__11716 (
            .O(N__55125),
            .I(N__55121));
    InMux I__11715 (
            .O(N__55124),
            .I(N__55118));
    LocalMux I__11714 (
            .O(N__55121),
            .I(N__55115));
    LocalMux I__11713 (
            .O(N__55118),
            .I(N__55110));
    Span4Mux_h I__11712 (
            .O(N__55115),
            .I(N__55107));
    InMux I__11711 (
            .O(N__55114),
            .I(N__55104));
    CascadeMux I__11710 (
            .O(N__55113),
            .I(N__55101));
    Span4Mux_h I__11709 (
            .O(N__55110),
            .I(N__55097));
    Span4Mux_v I__11708 (
            .O(N__55107),
            .I(N__55092));
    LocalMux I__11707 (
            .O(N__55104),
            .I(N__55092));
    InMux I__11706 (
            .O(N__55101),
            .I(N__55087));
    InMux I__11705 (
            .O(N__55100),
            .I(N__55087));
    Odrv4 I__11704 (
            .O(N__55097),
            .I(\c0.data_in_frame_8_1 ));
    Odrv4 I__11703 (
            .O(N__55092),
            .I(\c0.data_in_frame_8_1 ));
    LocalMux I__11702 (
            .O(N__55087),
            .I(\c0.data_in_frame_8_1 ));
    CascadeMux I__11701 (
            .O(N__55080),
            .I(\c0.n13_adj_4638_cascade_ ));
    InMux I__11700 (
            .O(N__55077),
            .I(N__55074));
    LocalMux I__11699 (
            .O(N__55074),
            .I(N__55071));
    Span4Mux_h I__11698 (
            .O(N__55071),
            .I(N__55066));
    InMux I__11697 (
            .O(N__55070),
            .I(N__55063));
    InMux I__11696 (
            .O(N__55069),
            .I(N__55060));
    Span4Mux_h I__11695 (
            .O(N__55066),
            .I(N__55057));
    LocalMux I__11694 (
            .O(N__55063),
            .I(\c0.data_in_frame_10_1 ));
    LocalMux I__11693 (
            .O(N__55060),
            .I(\c0.data_in_frame_10_1 ));
    Odrv4 I__11692 (
            .O(N__55057),
            .I(\c0.data_in_frame_10_1 ));
    CascadeMux I__11691 (
            .O(N__55050),
            .I(N__55046));
    InMux I__11690 (
            .O(N__55049),
            .I(N__55040));
    InMux I__11689 (
            .O(N__55046),
            .I(N__55040));
    CascadeMux I__11688 (
            .O(N__55045),
            .I(N__55037));
    LocalMux I__11687 (
            .O(N__55040),
            .I(N__55034));
    InMux I__11686 (
            .O(N__55037),
            .I(N__55031));
    Span4Mux_v I__11685 (
            .O(N__55034),
            .I(N__55028));
    LocalMux I__11684 (
            .O(N__55031),
            .I(\c0.data_in_frame_10_2 ));
    Odrv4 I__11683 (
            .O(N__55028),
            .I(\c0.data_in_frame_10_2 ));
    CascadeMux I__11682 (
            .O(N__55023),
            .I(N__55017));
    InMux I__11681 (
            .O(N__55022),
            .I(N__55014));
    InMux I__11680 (
            .O(N__55021),
            .I(N__55009));
    InMux I__11679 (
            .O(N__55020),
            .I(N__55009));
    InMux I__11678 (
            .O(N__55017),
            .I(N__55006));
    LocalMux I__11677 (
            .O(N__55014),
            .I(N__55003));
    LocalMux I__11676 (
            .O(N__55009),
            .I(N__55000));
    LocalMux I__11675 (
            .O(N__55006),
            .I(N__54995));
    Span4Mux_v I__11674 (
            .O(N__55003),
            .I(N__54995));
    Span4Mux_h I__11673 (
            .O(N__55000),
            .I(N__54992));
    Odrv4 I__11672 (
            .O(N__54995),
            .I(\c0.data_in_frame_9_7 ));
    Odrv4 I__11671 (
            .O(N__54992),
            .I(\c0.data_in_frame_9_7 ));
    CascadeMux I__11670 (
            .O(N__54987),
            .I(\c0.n22196_cascade_ ));
    InMux I__11669 (
            .O(N__54984),
            .I(N__54981));
    LocalMux I__11668 (
            .O(N__54981),
            .I(N__54978));
    Span4Mux_h I__11667 (
            .O(N__54978),
            .I(N__54975));
    Span4Mux_v I__11666 (
            .O(N__54975),
            .I(N__54972));
    Odrv4 I__11665 (
            .O(N__54972),
            .I(\c0.n12_adj_4258 ));
    InMux I__11664 (
            .O(N__54969),
            .I(N__54963));
    InMux I__11663 (
            .O(N__54968),
            .I(N__54963));
    LocalMux I__11662 (
            .O(N__54963),
            .I(\c0.data_in_frame_3_0 ));
    CascadeMux I__11661 (
            .O(N__54960),
            .I(N__54957));
    InMux I__11660 (
            .O(N__54957),
            .I(N__54954));
    LocalMux I__11659 (
            .O(N__54954),
            .I(\c0.n10_adj_4615 ));
    InMux I__11658 (
            .O(N__54951),
            .I(N__54947));
    CascadeMux I__11657 (
            .O(N__54950),
            .I(N__54944));
    LocalMux I__11656 (
            .O(N__54947),
            .I(N__54940));
    InMux I__11655 (
            .O(N__54944),
            .I(N__54937));
    InMux I__11654 (
            .O(N__54943),
            .I(N__54933));
    Span4Mux_h I__11653 (
            .O(N__54940),
            .I(N__54930));
    LocalMux I__11652 (
            .O(N__54937),
            .I(N__54927));
    InMux I__11651 (
            .O(N__54936),
            .I(N__54924));
    LocalMux I__11650 (
            .O(N__54933),
            .I(N__54921));
    Span4Mux_v I__11649 (
            .O(N__54930),
            .I(N__54918));
    Odrv4 I__11648 (
            .O(N__54927),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__11647 (
            .O(N__54924),
            .I(\c0.data_in_frame_3_1 ));
    Odrv12 I__11646 (
            .O(N__54921),
            .I(\c0.data_in_frame_3_1 ));
    Odrv4 I__11645 (
            .O(N__54918),
            .I(\c0.data_in_frame_3_1 ));
    InMux I__11644 (
            .O(N__54909),
            .I(N__54906));
    LocalMux I__11643 (
            .O(N__54906),
            .I(\c0.n7_adj_4300 ));
    SRMux I__11642 (
            .O(N__54903),
            .I(N__54900));
    LocalMux I__11641 (
            .O(N__54900),
            .I(N__54897));
    Odrv4 I__11640 (
            .O(N__54897),
            .I(\c0.n3_adj_4436 ));
    SRMux I__11639 (
            .O(N__54894),
            .I(N__54891));
    LocalMux I__11638 (
            .O(N__54891),
            .I(N__54888));
    Odrv4 I__11637 (
            .O(N__54888),
            .I(\c0.n3_adj_4376 ));
    InMux I__11636 (
            .O(N__54885),
            .I(N__54872));
    InMux I__11635 (
            .O(N__54884),
            .I(N__54872));
    InMux I__11634 (
            .O(N__54883),
            .I(N__54872));
    InMux I__11633 (
            .O(N__54882),
            .I(N__54863));
    InMux I__11632 (
            .O(N__54881),
            .I(N__54863));
    InMux I__11631 (
            .O(N__54880),
            .I(N__54863));
    InMux I__11630 (
            .O(N__54879),
            .I(N__54863));
    LocalMux I__11629 (
            .O(N__54872),
            .I(N__54822));
    LocalMux I__11628 (
            .O(N__54863),
            .I(N__54822));
    InMux I__11627 (
            .O(N__54862),
            .I(N__54815));
    InMux I__11626 (
            .O(N__54861),
            .I(N__54815));
    InMux I__11625 (
            .O(N__54860),
            .I(N__54815));
    InMux I__11624 (
            .O(N__54859),
            .I(N__54806));
    InMux I__11623 (
            .O(N__54858),
            .I(N__54806));
    InMux I__11622 (
            .O(N__54857),
            .I(N__54806));
    InMux I__11621 (
            .O(N__54856),
            .I(N__54806));
    InMux I__11620 (
            .O(N__54855),
            .I(N__54799));
    InMux I__11619 (
            .O(N__54854),
            .I(N__54799));
    InMux I__11618 (
            .O(N__54853),
            .I(N__54799));
    InMux I__11617 (
            .O(N__54852),
            .I(N__54790));
    InMux I__11616 (
            .O(N__54851),
            .I(N__54790));
    InMux I__11615 (
            .O(N__54850),
            .I(N__54790));
    InMux I__11614 (
            .O(N__54849),
            .I(N__54790));
    InMux I__11613 (
            .O(N__54848),
            .I(N__54783));
    InMux I__11612 (
            .O(N__54847),
            .I(N__54783));
    InMux I__11611 (
            .O(N__54846),
            .I(N__54783));
    InMux I__11610 (
            .O(N__54845),
            .I(N__54774));
    InMux I__11609 (
            .O(N__54844),
            .I(N__54774));
    InMux I__11608 (
            .O(N__54843),
            .I(N__54774));
    InMux I__11607 (
            .O(N__54842),
            .I(N__54774));
    InMux I__11606 (
            .O(N__54841),
            .I(N__54767));
    InMux I__11605 (
            .O(N__54840),
            .I(N__54767));
    InMux I__11604 (
            .O(N__54839),
            .I(N__54767));
    InMux I__11603 (
            .O(N__54838),
            .I(N__54758));
    InMux I__11602 (
            .O(N__54837),
            .I(N__54758));
    InMux I__11601 (
            .O(N__54836),
            .I(N__54758));
    InMux I__11600 (
            .O(N__54835),
            .I(N__54758));
    CascadeMux I__11599 (
            .O(N__54834),
            .I(N__54755));
    CascadeMux I__11598 (
            .O(N__54833),
            .I(N__54751));
    CascadeMux I__11597 (
            .O(N__54832),
            .I(N__54747));
    CascadeMux I__11596 (
            .O(N__54831),
            .I(N__54743));
    CascadeMux I__11595 (
            .O(N__54830),
            .I(N__54733));
    CascadeMux I__11594 (
            .O(N__54829),
            .I(N__54729));
    CascadeMux I__11593 (
            .O(N__54828),
            .I(N__54725));
    CascadeMux I__11592 (
            .O(N__54827),
            .I(N__54721));
    Span4Mux_s3_v I__11591 (
            .O(N__54822),
            .I(N__54695));
    LocalMux I__11590 (
            .O(N__54815),
            .I(N__54695));
    LocalMux I__11589 (
            .O(N__54806),
            .I(N__54695));
    LocalMux I__11588 (
            .O(N__54799),
            .I(N__54695));
    LocalMux I__11587 (
            .O(N__54790),
            .I(N__54695));
    LocalMux I__11586 (
            .O(N__54783),
            .I(N__54695));
    LocalMux I__11585 (
            .O(N__54774),
            .I(N__54695));
    LocalMux I__11584 (
            .O(N__54767),
            .I(N__54695));
    LocalMux I__11583 (
            .O(N__54758),
            .I(N__54695));
    InMux I__11582 (
            .O(N__54755),
            .I(N__54680));
    InMux I__11581 (
            .O(N__54754),
            .I(N__54680));
    InMux I__11580 (
            .O(N__54751),
            .I(N__54680));
    InMux I__11579 (
            .O(N__54750),
            .I(N__54680));
    InMux I__11578 (
            .O(N__54747),
            .I(N__54680));
    InMux I__11577 (
            .O(N__54746),
            .I(N__54680));
    InMux I__11576 (
            .O(N__54743),
            .I(N__54680));
    InMux I__11575 (
            .O(N__54742),
            .I(N__54673));
    InMux I__11574 (
            .O(N__54741),
            .I(N__54673));
    InMux I__11573 (
            .O(N__54740),
            .I(N__54673));
    InMux I__11572 (
            .O(N__54739),
            .I(N__54664));
    InMux I__11571 (
            .O(N__54738),
            .I(N__54664));
    InMux I__11570 (
            .O(N__54737),
            .I(N__54664));
    InMux I__11569 (
            .O(N__54736),
            .I(N__54664));
    InMux I__11568 (
            .O(N__54733),
            .I(N__54649));
    InMux I__11567 (
            .O(N__54732),
            .I(N__54649));
    InMux I__11566 (
            .O(N__54729),
            .I(N__54649));
    InMux I__11565 (
            .O(N__54728),
            .I(N__54649));
    InMux I__11564 (
            .O(N__54725),
            .I(N__54649));
    InMux I__11563 (
            .O(N__54724),
            .I(N__54649));
    InMux I__11562 (
            .O(N__54721),
            .I(N__54649));
    InMux I__11561 (
            .O(N__54720),
            .I(N__54642));
    InMux I__11560 (
            .O(N__54719),
            .I(N__54642));
    InMux I__11559 (
            .O(N__54718),
            .I(N__54642));
    InMux I__11558 (
            .O(N__54717),
            .I(N__54633));
    InMux I__11557 (
            .O(N__54716),
            .I(N__54633));
    InMux I__11556 (
            .O(N__54715),
            .I(N__54633));
    InMux I__11555 (
            .O(N__54714),
            .I(N__54633));
    Span4Mux_v I__11554 (
            .O(N__54695),
            .I(N__54615));
    LocalMux I__11553 (
            .O(N__54680),
            .I(N__54615));
    LocalMux I__11552 (
            .O(N__54673),
            .I(N__54615));
    LocalMux I__11551 (
            .O(N__54664),
            .I(N__54615));
    LocalMux I__11550 (
            .O(N__54649),
            .I(N__54615));
    LocalMux I__11549 (
            .O(N__54642),
            .I(N__54615));
    LocalMux I__11548 (
            .O(N__54633),
            .I(N__54615));
    CascadeMux I__11547 (
            .O(N__54632),
            .I(N__54590));
    CascadeMux I__11546 (
            .O(N__54631),
            .I(N__54586));
    CascadeMux I__11545 (
            .O(N__54630),
            .I(N__54582));
    Span4Mux_v I__11544 (
            .O(N__54615),
            .I(N__54566));
    InMux I__11543 (
            .O(N__54614),
            .I(N__54559));
    InMux I__11542 (
            .O(N__54613),
            .I(N__54559));
    InMux I__11541 (
            .O(N__54612),
            .I(N__54559));
    InMux I__11540 (
            .O(N__54611),
            .I(N__54550));
    InMux I__11539 (
            .O(N__54610),
            .I(N__54550));
    InMux I__11538 (
            .O(N__54609),
            .I(N__54550));
    InMux I__11537 (
            .O(N__54608),
            .I(N__54550));
    InMux I__11536 (
            .O(N__54607),
            .I(N__54543));
    InMux I__11535 (
            .O(N__54606),
            .I(N__54543));
    InMux I__11534 (
            .O(N__54605),
            .I(N__54543));
    InMux I__11533 (
            .O(N__54604),
            .I(N__54534));
    InMux I__11532 (
            .O(N__54603),
            .I(N__54534));
    InMux I__11531 (
            .O(N__54602),
            .I(N__54534));
    InMux I__11530 (
            .O(N__54601),
            .I(N__54534));
    InMux I__11529 (
            .O(N__54600),
            .I(N__54527));
    InMux I__11528 (
            .O(N__54599),
            .I(N__54527));
    InMux I__11527 (
            .O(N__54598),
            .I(N__54527));
    InMux I__11526 (
            .O(N__54597),
            .I(N__54518));
    InMux I__11525 (
            .O(N__54596),
            .I(N__54518));
    InMux I__11524 (
            .O(N__54595),
            .I(N__54518));
    InMux I__11523 (
            .O(N__54594),
            .I(N__54518));
    InMux I__11522 (
            .O(N__54593),
            .I(N__54475));
    InMux I__11521 (
            .O(N__54590),
            .I(N__54475));
    InMux I__11520 (
            .O(N__54589),
            .I(N__54475));
    InMux I__11519 (
            .O(N__54586),
            .I(N__54475));
    InMux I__11518 (
            .O(N__54585),
            .I(N__54475));
    InMux I__11517 (
            .O(N__54582),
            .I(N__54475));
    InMux I__11516 (
            .O(N__54581),
            .I(N__54475));
    CascadeMux I__11515 (
            .O(N__54580),
            .I(N__54471));
    CascadeMux I__11514 (
            .O(N__54579),
            .I(N__54467));
    CascadeMux I__11513 (
            .O(N__54578),
            .I(N__54463));
    CascadeMux I__11512 (
            .O(N__54577),
            .I(N__54458));
    CascadeMux I__11511 (
            .O(N__54576),
            .I(N__54454));
    CascadeMux I__11510 (
            .O(N__54575),
            .I(N__54450));
    CascadeMux I__11509 (
            .O(N__54574),
            .I(N__54445));
    CascadeMux I__11508 (
            .O(N__54573),
            .I(N__54441));
    CascadeMux I__11507 (
            .O(N__54572),
            .I(N__54437));
    CascadeMux I__11506 (
            .O(N__54571),
            .I(N__54432));
    CascadeMux I__11505 (
            .O(N__54570),
            .I(N__54428));
    CascadeMux I__11504 (
            .O(N__54569),
            .I(N__54424));
    Span4Mux_h I__11503 (
            .O(N__54566),
            .I(N__54402));
    LocalMux I__11502 (
            .O(N__54559),
            .I(N__54402));
    LocalMux I__11501 (
            .O(N__54550),
            .I(N__54402));
    LocalMux I__11500 (
            .O(N__54543),
            .I(N__54402));
    LocalMux I__11499 (
            .O(N__54534),
            .I(N__54402));
    LocalMux I__11498 (
            .O(N__54527),
            .I(N__54402));
    LocalMux I__11497 (
            .O(N__54518),
            .I(N__54402));
    InMux I__11496 (
            .O(N__54517),
            .I(N__54395));
    InMux I__11495 (
            .O(N__54516),
            .I(N__54395));
    InMux I__11494 (
            .O(N__54515),
            .I(N__54395));
    InMux I__11493 (
            .O(N__54514),
            .I(N__54386));
    InMux I__11492 (
            .O(N__54513),
            .I(N__54386));
    InMux I__11491 (
            .O(N__54512),
            .I(N__54386));
    InMux I__11490 (
            .O(N__54511),
            .I(N__54386));
    InMux I__11489 (
            .O(N__54510),
            .I(N__54379));
    InMux I__11488 (
            .O(N__54509),
            .I(N__54379));
    InMux I__11487 (
            .O(N__54508),
            .I(N__54379));
    InMux I__11486 (
            .O(N__54507),
            .I(N__54370));
    InMux I__11485 (
            .O(N__54506),
            .I(N__54370));
    InMux I__11484 (
            .O(N__54505),
            .I(N__54370));
    InMux I__11483 (
            .O(N__54504),
            .I(N__54370));
    InMux I__11482 (
            .O(N__54503),
            .I(N__54363));
    InMux I__11481 (
            .O(N__54502),
            .I(N__54363));
    InMux I__11480 (
            .O(N__54501),
            .I(N__54363));
    InMux I__11479 (
            .O(N__54500),
            .I(N__54354));
    InMux I__11478 (
            .O(N__54499),
            .I(N__54354));
    InMux I__11477 (
            .O(N__54498),
            .I(N__54354));
    InMux I__11476 (
            .O(N__54497),
            .I(N__54354));
    InMux I__11475 (
            .O(N__54496),
            .I(N__54347));
    InMux I__11474 (
            .O(N__54495),
            .I(N__54347));
    InMux I__11473 (
            .O(N__54494),
            .I(N__54347));
    InMux I__11472 (
            .O(N__54493),
            .I(N__54338));
    InMux I__11471 (
            .O(N__54492),
            .I(N__54338));
    InMux I__11470 (
            .O(N__54491),
            .I(N__54338));
    InMux I__11469 (
            .O(N__54490),
            .I(N__54338));
    LocalMux I__11468 (
            .O(N__54475),
            .I(N__54304));
    InMux I__11467 (
            .O(N__54474),
            .I(N__54289));
    InMux I__11466 (
            .O(N__54471),
            .I(N__54289));
    InMux I__11465 (
            .O(N__54470),
            .I(N__54289));
    InMux I__11464 (
            .O(N__54467),
            .I(N__54289));
    InMux I__11463 (
            .O(N__54466),
            .I(N__54289));
    InMux I__11462 (
            .O(N__54463),
            .I(N__54289));
    InMux I__11461 (
            .O(N__54462),
            .I(N__54289));
    InMux I__11460 (
            .O(N__54461),
            .I(N__54274));
    InMux I__11459 (
            .O(N__54458),
            .I(N__54274));
    InMux I__11458 (
            .O(N__54457),
            .I(N__54274));
    InMux I__11457 (
            .O(N__54454),
            .I(N__54274));
    InMux I__11456 (
            .O(N__54453),
            .I(N__54274));
    InMux I__11455 (
            .O(N__54450),
            .I(N__54274));
    InMux I__11454 (
            .O(N__54449),
            .I(N__54274));
    InMux I__11453 (
            .O(N__54448),
            .I(N__54259));
    InMux I__11452 (
            .O(N__54445),
            .I(N__54259));
    InMux I__11451 (
            .O(N__54444),
            .I(N__54259));
    InMux I__11450 (
            .O(N__54441),
            .I(N__54259));
    InMux I__11449 (
            .O(N__54440),
            .I(N__54259));
    InMux I__11448 (
            .O(N__54437),
            .I(N__54259));
    InMux I__11447 (
            .O(N__54436),
            .I(N__54259));
    InMux I__11446 (
            .O(N__54435),
            .I(N__54244));
    InMux I__11445 (
            .O(N__54432),
            .I(N__54244));
    InMux I__11444 (
            .O(N__54431),
            .I(N__54244));
    InMux I__11443 (
            .O(N__54428),
            .I(N__54244));
    InMux I__11442 (
            .O(N__54427),
            .I(N__54244));
    InMux I__11441 (
            .O(N__54424),
            .I(N__54244));
    InMux I__11440 (
            .O(N__54423),
            .I(N__54244));
    CascadeMux I__11439 (
            .O(N__54422),
            .I(N__54240));
    CascadeMux I__11438 (
            .O(N__54421),
            .I(N__54236));
    CascadeMux I__11437 (
            .O(N__54420),
            .I(N__54232));
    CascadeMux I__11436 (
            .O(N__54419),
            .I(N__54227));
    CascadeMux I__11435 (
            .O(N__54418),
            .I(N__54223));
    CascadeMux I__11434 (
            .O(N__54417),
            .I(N__54219));
    Span4Mux_v I__11433 (
            .O(N__54402),
            .I(N__54199));
    LocalMux I__11432 (
            .O(N__54395),
            .I(N__54199));
    LocalMux I__11431 (
            .O(N__54386),
            .I(N__54199));
    LocalMux I__11430 (
            .O(N__54379),
            .I(N__54199));
    LocalMux I__11429 (
            .O(N__54370),
            .I(N__54199));
    LocalMux I__11428 (
            .O(N__54363),
            .I(N__54199));
    LocalMux I__11427 (
            .O(N__54354),
            .I(N__54199));
    LocalMux I__11426 (
            .O(N__54347),
            .I(N__54199));
    LocalMux I__11425 (
            .O(N__54338),
            .I(N__54199));
    InMux I__11424 (
            .O(N__54337),
            .I(N__54192));
    InMux I__11423 (
            .O(N__54336),
            .I(N__54192));
    InMux I__11422 (
            .O(N__54335),
            .I(N__54192));
    InMux I__11421 (
            .O(N__54334),
            .I(N__54183));
    InMux I__11420 (
            .O(N__54333),
            .I(N__54183));
    InMux I__11419 (
            .O(N__54332),
            .I(N__54183));
    InMux I__11418 (
            .O(N__54331),
            .I(N__54183));
    InMux I__11417 (
            .O(N__54330),
            .I(N__54176));
    InMux I__11416 (
            .O(N__54329),
            .I(N__54176));
    InMux I__11415 (
            .O(N__54328),
            .I(N__54176));
    InMux I__11414 (
            .O(N__54327),
            .I(N__54167));
    InMux I__11413 (
            .O(N__54326),
            .I(N__54167));
    InMux I__11412 (
            .O(N__54325),
            .I(N__54167));
    InMux I__11411 (
            .O(N__54324),
            .I(N__54167));
    InMux I__11410 (
            .O(N__54323),
            .I(N__54160));
    InMux I__11409 (
            .O(N__54322),
            .I(N__54160));
    InMux I__11408 (
            .O(N__54321),
            .I(N__54160));
    InMux I__11407 (
            .O(N__54320),
            .I(N__54151));
    InMux I__11406 (
            .O(N__54319),
            .I(N__54151));
    InMux I__11405 (
            .O(N__54318),
            .I(N__54151));
    InMux I__11404 (
            .O(N__54317),
            .I(N__54151));
    CascadeMux I__11403 (
            .O(N__54316),
            .I(N__54147));
    CascadeMux I__11402 (
            .O(N__54315),
            .I(N__54143));
    CascadeMux I__11401 (
            .O(N__54314),
            .I(N__54139));
    InMux I__11400 (
            .O(N__54313),
            .I(N__54124));
    InMux I__11399 (
            .O(N__54312),
            .I(N__54124));
    InMux I__11398 (
            .O(N__54311),
            .I(N__54124));
    InMux I__11397 (
            .O(N__54310),
            .I(N__54115));
    InMux I__11396 (
            .O(N__54309),
            .I(N__54115));
    InMux I__11395 (
            .O(N__54308),
            .I(N__54115));
    InMux I__11394 (
            .O(N__54307),
            .I(N__54115));
    Span4Mux_s0_v I__11393 (
            .O(N__54304),
            .I(N__54106));
    LocalMux I__11392 (
            .O(N__54289),
            .I(N__54106));
    LocalMux I__11391 (
            .O(N__54274),
            .I(N__54106));
    LocalMux I__11390 (
            .O(N__54259),
            .I(N__54106));
    LocalMux I__11389 (
            .O(N__54244),
            .I(N__54103));
    InMux I__11388 (
            .O(N__54243),
            .I(N__54088));
    InMux I__11387 (
            .O(N__54240),
            .I(N__54088));
    InMux I__11386 (
            .O(N__54239),
            .I(N__54088));
    InMux I__11385 (
            .O(N__54236),
            .I(N__54088));
    InMux I__11384 (
            .O(N__54235),
            .I(N__54088));
    InMux I__11383 (
            .O(N__54232),
            .I(N__54088));
    InMux I__11382 (
            .O(N__54231),
            .I(N__54088));
    InMux I__11381 (
            .O(N__54230),
            .I(N__54073));
    InMux I__11380 (
            .O(N__54227),
            .I(N__54073));
    InMux I__11379 (
            .O(N__54226),
            .I(N__54073));
    InMux I__11378 (
            .O(N__54223),
            .I(N__54073));
    InMux I__11377 (
            .O(N__54222),
            .I(N__54073));
    InMux I__11376 (
            .O(N__54219),
            .I(N__54073));
    InMux I__11375 (
            .O(N__54218),
            .I(N__54073));
    Span4Mux_v I__11374 (
            .O(N__54199),
            .I(N__54058));
    LocalMux I__11373 (
            .O(N__54192),
            .I(N__54058));
    LocalMux I__11372 (
            .O(N__54183),
            .I(N__54058));
    LocalMux I__11371 (
            .O(N__54176),
            .I(N__54058));
    LocalMux I__11370 (
            .O(N__54167),
            .I(N__54058));
    LocalMux I__11369 (
            .O(N__54160),
            .I(N__54058));
    LocalMux I__11368 (
            .O(N__54151),
            .I(N__54058));
    InMux I__11367 (
            .O(N__54150),
            .I(N__54043));
    InMux I__11366 (
            .O(N__54147),
            .I(N__54043));
    InMux I__11365 (
            .O(N__54146),
            .I(N__54043));
    InMux I__11364 (
            .O(N__54143),
            .I(N__54043));
    InMux I__11363 (
            .O(N__54142),
            .I(N__54043));
    InMux I__11362 (
            .O(N__54139),
            .I(N__54043));
    InMux I__11361 (
            .O(N__54138),
            .I(N__54043));
    InMux I__11360 (
            .O(N__54137),
            .I(N__54036));
    InMux I__11359 (
            .O(N__54136),
            .I(N__54036));
    InMux I__11358 (
            .O(N__54135),
            .I(N__54036));
    InMux I__11357 (
            .O(N__54134),
            .I(N__54027));
    InMux I__11356 (
            .O(N__54133),
            .I(N__54027));
    InMux I__11355 (
            .O(N__54132),
            .I(N__54027));
    InMux I__11354 (
            .O(N__54131),
            .I(N__54027));
    LocalMux I__11353 (
            .O(N__54124),
            .I(N__54015));
    LocalMux I__11352 (
            .O(N__54115),
            .I(N__54015));
    Span4Mux_v I__11351 (
            .O(N__54106),
            .I(N__54002));
    Span4Mux_h I__11350 (
            .O(N__54103),
            .I(N__54002));
    LocalMux I__11349 (
            .O(N__54088),
            .I(N__54002));
    LocalMux I__11348 (
            .O(N__54073),
            .I(N__54002));
    Span4Mux_v I__11347 (
            .O(N__54058),
            .I(N__54002));
    LocalMux I__11346 (
            .O(N__54043),
            .I(N__54002));
    LocalMux I__11345 (
            .O(N__54036),
            .I(N__53990));
    LocalMux I__11344 (
            .O(N__54027),
            .I(N__53990));
    InMux I__11343 (
            .O(N__54026),
            .I(N__53983));
    InMux I__11342 (
            .O(N__54025),
            .I(N__53983));
    InMux I__11341 (
            .O(N__54024),
            .I(N__53983));
    InMux I__11340 (
            .O(N__54023),
            .I(N__53974));
    InMux I__11339 (
            .O(N__54022),
            .I(N__53974));
    InMux I__11338 (
            .O(N__54021),
            .I(N__53974));
    InMux I__11337 (
            .O(N__54020),
            .I(N__53974));
    Span4Mux_h I__11336 (
            .O(N__54015),
            .I(N__53971));
    Span4Mux_v I__11335 (
            .O(N__54002),
            .I(N__53968));
    InMux I__11334 (
            .O(N__54001),
            .I(N__53961));
    InMux I__11333 (
            .O(N__54000),
            .I(N__53961));
    InMux I__11332 (
            .O(N__53999),
            .I(N__53961));
    InMux I__11331 (
            .O(N__53998),
            .I(N__53952));
    InMux I__11330 (
            .O(N__53997),
            .I(N__53952));
    InMux I__11329 (
            .O(N__53996),
            .I(N__53952));
    InMux I__11328 (
            .O(N__53995),
            .I(N__53952));
    Span12Mux_h I__11327 (
            .O(N__53990),
            .I(N__53949));
    LocalMux I__11326 (
            .O(N__53983),
            .I(N__53944));
    LocalMux I__11325 (
            .O(N__53974),
            .I(N__53944));
    Sp12to4 I__11324 (
            .O(N__53971),
            .I(N__53941));
    Sp12to4 I__11323 (
            .O(N__53968),
            .I(N__53934));
    LocalMux I__11322 (
            .O(N__53961),
            .I(N__53934));
    LocalMux I__11321 (
            .O(N__53952),
            .I(N__53934));
    Span12Mux_v I__11320 (
            .O(N__53949),
            .I(N__53929));
    Span12Mux_h I__11319 (
            .O(N__53944),
            .I(N__53929));
    Span12Mux_s8_v I__11318 (
            .O(N__53941),
            .I(N__53924));
    Span12Mux_h I__11317 (
            .O(N__53934),
            .I(N__53924));
    Odrv12 I__11316 (
            .O(N__53929),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__11315 (
            .O(N__53924),
            .I(CONSTANT_ONE_NET));
    InMux I__11314 (
            .O(N__53919),
            .I(bfn_19_32_0_));
    CascadeMux I__11313 (
            .O(N__53916),
            .I(N__53912));
    InMux I__11312 (
            .O(N__53915),
            .I(N__53905));
    InMux I__11311 (
            .O(N__53912),
            .I(N__53902));
    InMux I__11310 (
            .O(N__53911),
            .I(N__53895));
    InMux I__11309 (
            .O(N__53910),
            .I(N__53895));
    InMux I__11308 (
            .O(N__53909),
            .I(N__53895));
    InMux I__11307 (
            .O(N__53908),
            .I(N__53891));
    LocalMux I__11306 (
            .O(N__53905),
            .I(N__53888));
    LocalMux I__11305 (
            .O(N__53902),
            .I(N__53885));
    LocalMux I__11304 (
            .O(N__53895),
            .I(N__53882));
    InMux I__11303 (
            .O(N__53894),
            .I(N__53878));
    LocalMux I__11302 (
            .O(N__53891),
            .I(N__53874));
    Span4Mux_v I__11301 (
            .O(N__53888),
            .I(N__53871));
    Span4Mux_h I__11300 (
            .O(N__53885),
            .I(N__53866));
    Span4Mux_v I__11299 (
            .O(N__53882),
            .I(N__53866));
    InMux I__11298 (
            .O(N__53881),
            .I(N__53863));
    LocalMux I__11297 (
            .O(N__53878),
            .I(N__53860));
    InMux I__11296 (
            .O(N__53877),
            .I(N__53857));
    Span4Mux_v I__11295 (
            .O(N__53874),
            .I(N__53854));
    Span4Mux_v I__11294 (
            .O(N__53871),
            .I(N__53851));
    Span4Mux_v I__11293 (
            .O(N__53866),
            .I(N__53848));
    LocalMux I__11292 (
            .O(N__53863),
            .I(N__53843));
    Span12Mux_v I__11291 (
            .O(N__53860),
            .I(N__53843));
    LocalMux I__11290 (
            .O(N__53857),
            .I(N__53838));
    Span4Mux_v I__11289 (
            .O(N__53854),
            .I(N__53838));
    Span4Mux_h I__11288 (
            .O(N__53851),
            .I(N__53835));
    Span4Mux_h I__11287 (
            .O(N__53848),
            .I(N__53832));
    Odrv12 I__11286 (
            .O(N__53843),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__11285 (
            .O(N__53838),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__11284 (
            .O(N__53835),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__11283 (
            .O(N__53832),
            .I(\c0.FRAME_MATCHER_i_31 ));
    SRMux I__11282 (
            .O(N__53823),
            .I(N__53820));
    LocalMux I__11281 (
            .O(N__53820),
            .I(N__53817));
    Odrv12 I__11280 (
            .O(N__53817),
            .I(\c0.n3_adj_4373 ));
    InMux I__11279 (
            .O(N__53814),
            .I(N__53811));
    LocalMux I__11278 (
            .O(N__53811),
            .I(N__53808));
    Span4Mux_h I__11277 (
            .O(N__53808),
            .I(N__53804));
    InMux I__11276 (
            .O(N__53807),
            .I(N__53799));
    Span4Mux_v I__11275 (
            .O(N__53804),
            .I(N__53796));
    InMux I__11274 (
            .O(N__53803),
            .I(N__53793));
    InMux I__11273 (
            .O(N__53802),
            .I(N__53790));
    LocalMux I__11272 (
            .O(N__53799),
            .I(N__53787));
    Span4Mux_v I__11271 (
            .O(N__53796),
            .I(N__53782));
    LocalMux I__11270 (
            .O(N__53793),
            .I(N__53782));
    LocalMux I__11269 (
            .O(N__53790),
            .I(N__53779));
    Span4Mux_h I__11268 (
            .O(N__53787),
            .I(N__53776));
    Odrv4 I__11267 (
            .O(N__53782),
            .I(\c0.n17856 ));
    Odrv4 I__11266 (
            .O(N__53779),
            .I(\c0.n17856 ));
    Odrv4 I__11265 (
            .O(N__53776),
            .I(\c0.n17856 ));
    InMux I__11264 (
            .O(N__53769),
            .I(N__53761));
    InMux I__11263 (
            .O(N__53768),
            .I(N__53756));
    InMux I__11262 (
            .O(N__53767),
            .I(N__53753));
    InMux I__11261 (
            .O(N__53766),
            .I(N__53750));
    InMux I__11260 (
            .O(N__53765),
            .I(N__53737));
    InMux I__11259 (
            .O(N__53764),
            .I(N__53734));
    LocalMux I__11258 (
            .O(N__53761),
            .I(N__53731));
    InMux I__11257 (
            .O(N__53760),
            .I(N__53728));
    InMux I__11256 (
            .O(N__53759),
            .I(N__53725));
    LocalMux I__11255 (
            .O(N__53756),
            .I(N__53717));
    LocalMux I__11254 (
            .O(N__53753),
            .I(N__53717));
    LocalMux I__11253 (
            .O(N__53750),
            .I(N__53717));
    InMux I__11252 (
            .O(N__53749),
            .I(N__53714));
    InMux I__11251 (
            .O(N__53748),
            .I(N__53709));
    InMux I__11250 (
            .O(N__53747),
            .I(N__53706));
    InMux I__11249 (
            .O(N__53746),
            .I(N__53703));
    InMux I__11248 (
            .O(N__53745),
            .I(N__53700));
    InMux I__11247 (
            .O(N__53744),
            .I(N__53689));
    InMux I__11246 (
            .O(N__53743),
            .I(N__53686));
    InMux I__11245 (
            .O(N__53742),
            .I(N__53683));
    InMux I__11244 (
            .O(N__53741),
            .I(N__53680));
    InMux I__11243 (
            .O(N__53740),
            .I(N__53677));
    LocalMux I__11242 (
            .O(N__53737),
            .I(N__53666));
    LocalMux I__11241 (
            .O(N__53734),
            .I(N__53666));
    Sp12to4 I__11240 (
            .O(N__53731),
            .I(N__53666));
    LocalMux I__11239 (
            .O(N__53728),
            .I(N__53666));
    LocalMux I__11238 (
            .O(N__53725),
            .I(N__53666));
    InMux I__11237 (
            .O(N__53724),
            .I(N__53662));
    Span4Mux_v I__11236 (
            .O(N__53717),
            .I(N__53657));
    LocalMux I__11235 (
            .O(N__53714),
            .I(N__53657));
    InMux I__11234 (
            .O(N__53713),
            .I(N__53654));
    InMux I__11233 (
            .O(N__53712),
            .I(N__53651));
    LocalMux I__11232 (
            .O(N__53709),
            .I(N__53642));
    LocalMux I__11231 (
            .O(N__53706),
            .I(N__53642));
    LocalMux I__11230 (
            .O(N__53703),
            .I(N__53642));
    LocalMux I__11229 (
            .O(N__53700),
            .I(N__53642));
    InMux I__11228 (
            .O(N__53699),
            .I(N__53637));
    InMux I__11227 (
            .O(N__53698),
            .I(N__53634));
    InMux I__11226 (
            .O(N__53697),
            .I(N__53631));
    InMux I__11225 (
            .O(N__53696),
            .I(N__53628));
    InMux I__11224 (
            .O(N__53695),
            .I(N__53625));
    InMux I__11223 (
            .O(N__53694),
            .I(N__53622));
    InMux I__11222 (
            .O(N__53693),
            .I(N__53619));
    InMux I__11221 (
            .O(N__53692),
            .I(N__53616));
    LocalMux I__11220 (
            .O(N__53689),
            .I(N__53603));
    LocalMux I__11219 (
            .O(N__53686),
            .I(N__53603));
    LocalMux I__11218 (
            .O(N__53683),
            .I(N__53603));
    LocalMux I__11217 (
            .O(N__53680),
            .I(N__53603));
    LocalMux I__11216 (
            .O(N__53677),
            .I(N__53603));
    Span12Mux_s8_v I__11215 (
            .O(N__53666),
            .I(N__53603));
    InMux I__11214 (
            .O(N__53665),
            .I(N__53600));
    LocalMux I__11213 (
            .O(N__53662),
            .I(N__53589));
    Sp12to4 I__11212 (
            .O(N__53657),
            .I(N__53589));
    LocalMux I__11211 (
            .O(N__53654),
            .I(N__53589));
    LocalMux I__11210 (
            .O(N__53651),
            .I(N__53589));
    Span12Mux_v I__11209 (
            .O(N__53642),
            .I(N__53589));
    InMux I__11208 (
            .O(N__53641),
            .I(N__53586));
    InMux I__11207 (
            .O(N__53640),
            .I(N__53583));
    LocalMux I__11206 (
            .O(N__53637),
            .I(N__53580));
    LocalMux I__11205 (
            .O(N__53634),
            .I(N__53563));
    LocalMux I__11204 (
            .O(N__53631),
            .I(N__53563));
    LocalMux I__11203 (
            .O(N__53628),
            .I(N__53563));
    LocalMux I__11202 (
            .O(N__53625),
            .I(N__53563));
    LocalMux I__11201 (
            .O(N__53622),
            .I(N__53563));
    LocalMux I__11200 (
            .O(N__53619),
            .I(N__53563));
    LocalMux I__11199 (
            .O(N__53616),
            .I(N__53563));
    Span12Mux_v I__11198 (
            .O(N__53603),
            .I(N__53563));
    LocalMux I__11197 (
            .O(N__53600),
            .I(N__53558));
    Span12Mux_v I__11196 (
            .O(N__53589),
            .I(N__53558));
    LocalMux I__11195 (
            .O(N__53586),
            .I(\c0.n1306 ));
    LocalMux I__11194 (
            .O(N__53583),
            .I(\c0.n1306 ));
    Odrv4 I__11193 (
            .O(N__53580),
            .I(\c0.n1306 ));
    Odrv12 I__11192 (
            .O(N__53563),
            .I(\c0.n1306 ));
    Odrv12 I__11191 (
            .O(N__53558),
            .I(\c0.n1306 ));
    InMux I__11190 (
            .O(N__53547),
            .I(N__53544));
    LocalMux I__11189 (
            .O(N__53544),
            .I(N__53539));
    InMux I__11188 (
            .O(N__53543),
            .I(N__53536));
    InMux I__11187 (
            .O(N__53542),
            .I(N__53533));
    Span4Mux_h I__11186 (
            .O(N__53539),
            .I(N__53530));
    LocalMux I__11185 (
            .O(N__53536),
            .I(\c0.FRAME_MATCHER_i_29 ));
    LocalMux I__11184 (
            .O(N__53533),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__11183 (
            .O(N__53530),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__11182 (
            .O(N__53523),
            .I(bfn_19_30_0_));
    SRMux I__11181 (
            .O(N__53520),
            .I(N__53517));
    LocalMux I__11180 (
            .O(N__53517),
            .I(\c0.n3_adj_4378 ));
    InMux I__11179 (
            .O(N__53514),
            .I(N__53511));
    LocalMux I__11178 (
            .O(N__53511),
            .I(N__53506));
    InMux I__11177 (
            .O(N__53510),
            .I(N__53503));
    InMux I__11176 (
            .O(N__53509),
            .I(N__53500));
    Span4Mux_v I__11175 (
            .O(N__53506),
            .I(N__53497));
    LocalMux I__11174 (
            .O(N__53503),
            .I(\c0.FRAME_MATCHER_i_30 ));
    LocalMux I__11173 (
            .O(N__53500),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__11172 (
            .O(N__53497),
            .I(\c0.FRAME_MATCHER_i_30 ));
    InMux I__11171 (
            .O(N__53490),
            .I(bfn_19_31_0_));
    CascadeMux I__11170 (
            .O(N__53487),
            .I(N__53484));
    InMux I__11169 (
            .O(N__53484),
            .I(N__53481));
    LocalMux I__11168 (
            .O(N__53481),
            .I(N__53476));
    InMux I__11167 (
            .O(N__53480),
            .I(N__53473));
    InMux I__11166 (
            .O(N__53479),
            .I(N__53470));
    Span4Mux_h I__11165 (
            .O(N__53476),
            .I(N__53467));
    LocalMux I__11164 (
            .O(N__53473),
            .I(\c0.FRAME_MATCHER_i_28 ));
    LocalMux I__11163 (
            .O(N__53470),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__11162 (
            .O(N__53467),
            .I(\c0.FRAME_MATCHER_i_28 ));
    InMux I__11161 (
            .O(N__53460),
            .I(bfn_19_29_0_));
    SRMux I__11160 (
            .O(N__53457),
            .I(N__53454));
    LocalMux I__11159 (
            .O(N__53454),
            .I(N__53451));
    Odrv12 I__11158 (
            .O(N__53451),
            .I(\c0.n3_adj_4380 ));
    InMux I__11157 (
            .O(N__53448),
            .I(N__53445));
    LocalMux I__11156 (
            .O(N__53445),
            .I(N__53442));
    Span4Mux_v I__11155 (
            .O(N__53442),
            .I(N__53437));
    InMux I__11154 (
            .O(N__53441),
            .I(N__53434));
    InMux I__11153 (
            .O(N__53440),
            .I(N__53431));
    Span4Mux_h I__11152 (
            .O(N__53437),
            .I(N__53428));
    LocalMux I__11151 (
            .O(N__53434),
            .I(\c0.FRAME_MATCHER_i_27 ));
    LocalMux I__11150 (
            .O(N__53431),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv4 I__11149 (
            .O(N__53428),
            .I(\c0.FRAME_MATCHER_i_27 ));
    InMux I__11148 (
            .O(N__53421),
            .I(bfn_19_28_0_));
    SRMux I__11147 (
            .O(N__53418),
            .I(N__53415));
    LocalMux I__11146 (
            .O(N__53415),
            .I(N__53412));
    Odrv4 I__11145 (
            .O(N__53412),
            .I(\c0.n3_adj_4382 ));
    InMux I__11144 (
            .O(N__53409),
            .I(N__53405));
    InMux I__11143 (
            .O(N__53408),
            .I(N__53401));
    LocalMux I__11142 (
            .O(N__53405),
            .I(N__53398));
    InMux I__11141 (
            .O(N__53404),
            .I(N__53395));
    LocalMux I__11140 (
            .O(N__53401),
            .I(N__53390));
    Span4Mux_v I__11139 (
            .O(N__53398),
            .I(N__53390));
    LocalMux I__11138 (
            .O(N__53395),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__11137 (
            .O(N__53390),
            .I(\c0.FRAME_MATCHER_i_26 ));
    InMux I__11136 (
            .O(N__53385),
            .I(bfn_19_27_0_));
    SRMux I__11135 (
            .O(N__53382),
            .I(N__53379));
    LocalMux I__11134 (
            .O(N__53379),
            .I(\c0.n3_adj_4384 ));
    InMux I__11133 (
            .O(N__53376),
            .I(N__53371));
    InMux I__11132 (
            .O(N__53375),
            .I(N__53368));
    InMux I__11131 (
            .O(N__53374),
            .I(N__53365));
    LocalMux I__11130 (
            .O(N__53371),
            .I(N__53362));
    LocalMux I__11129 (
            .O(N__53368),
            .I(\c0.FRAME_MATCHER_i_25 ));
    LocalMux I__11128 (
            .O(N__53365),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__11127 (
            .O(N__53362),
            .I(\c0.FRAME_MATCHER_i_25 ));
    InMux I__11126 (
            .O(N__53355),
            .I(bfn_19_26_0_));
    SRMux I__11125 (
            .O(N__53352),
            .I(N__53349));
    LocalMux I__11124 (
            .O(N__53349),
            .I(\c0.n3_adj_4386 ));
    InMux I__11123 (
            .O(N__53346),
            .I(N__53343));
    LocalMux I__11122 (
            .O(N__53343),
            .I(N__53338));
    InMux I__11121 (
            .O(N__53342),
            .I(N__53335));
    InMux I__11120 (
            .O(N__53341),
            .I(N__53332));
    Odrv4 I__11119 (
            .O(N__53338),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__11118 (
            .O(N__53335),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__11117 (
            .O(N__53332),
            .I(\c0.FRAME_MATCHER_i_24 ));
    InMux I__11116 (
            .O(N__53325),
            .I(bfn_19_25_0_));
    SRMux I__11115 (
            .O(N__53322),
            .I(N__53319));
    LocalMux I__11114 (
            .O(N__53319),
            .I(N__53316));
    Odrv12 I__11113 (
            .O(N__53316),
            .I(\c0.n3_adj_4388 ));
    CascadeMux I__11112 (
            .O(N__53313),
            .I(N__53310));
    InMux I__11111 (
            .O(N__53310),
            .I(N__53306));
    InMux I__11110 (
            .O(N__53309),
            .I(N__53303));
    LocalMux I__11109 (
            .O(N__53306),
            .I(N__53299));
    LocalMux I__11108 (
            .O(N__53303),
            .I(N__53296));
    InMux I__11107 (
            .O(N__53302),
            .I(N__53293));
    Span4Mux_h I__11106 (
            .O(N__53299),
            .I(N__53290));
    Odrv4 I__11105 (
            .O(N__53296),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__11104 (
            .O(N__53293),
            .I(\c0.FRAME_MATCHER_i_23 ));
    Odrv4 I__11103 (
            .O(N__53290),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__11102 (
            .O(N__53283),
            .I(bfn_19_24_0_));
    SRMux I__11101 (
            .O(N__53280),
            .I(N__53277));
    LocalMux I__11100 (
            .O(N__53277),
            .I(N__53274));
    Odrv12 I__11099 (
            .O(N__53274),
            .I(\c0.n3_adj_4390 ));
    InMux I__11098 (
            .O(N__53271),
            .I(N__53267));
    InMux I__11097 (
            .O(N__53270),
            .I(N__53264));
    LocalMux I__11096 (
            .O(N__53267),
            .I(N__53258));
    LocalMux I__11095 (
            .O(N__53264),
            .I(N__53258));
    InMux I__11094 (
            .O(N__53263),
            .I(N__53255));
    Span4Mux_v I__11093 (
            .O(N__53258),
            .I(N__53252));
    LocalMux I__11092 (
            .O(N__53255),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__11091 (
            .O(N__53252),
            .I(\c0.FRAME_MATCHER_i_22 ));
    InMux I__11090 (
            .O(N__53247),
            .I(bfn_19_23_0_));
    SRMux I__11089 (
            .O(N__53244),
            .I(N__53241));
    LocalMux I__11088 (
            .O(N__53241),
            .I(N__53238));
    Span4Mux_h I__11087 (
            .O(N__53238),
            .I(N__53235));
    Odrv4 I__11086 (
            .O(N__53235),
            .I(\c0.n3_adj_4392 ));
    SRMux I__11085 (
            .O(N__53232),
            .I(N__53229));
    LocalMux I__11084 (
            .O(N__53229),
            .I(N__53226));
    Span4Mux_v I__11083 (
            .O(N__53226),
            .I(N__53223));
    Odrv4 I__11082 (
            .O(N__53223),
            .I(\c0.n3_adj_4396 ));
    InMux I__11081 (
            .O(N__53220),
            .I(N__53216));
    InMux I__11080 (
            .O(N__53219),
            .I(N__53213));
    LocalMux I__11079 (
            .O(N__53216),
            .I(N__53207));
    LocalMux I__11078 (
            .O(N__53213),
            .I(N__53207));
    InMux I__11077 (
            .O(N__53212),
            .I(N__53204));
    Span4Mux_v I__11076 (
            .O(N__53207),
            .I(N__53201));
    LocalMux I__11075 (
            .O(N__53204),
            .I(\c0.FRAME_MATCHER_i_21 ));
    Odrv4 I__11074 (
            .O(N__53201),
            .I(\c0.FRAME_MATCHER_i_21 ));
    InMux I__11073 (
            .O(N__53196),
            .I(bfn_19_22_0_));
    SRMux I__11072 (
            .O(N__53193),
            .I(N__53190));
    LocalMux I__11071 (
            .O(N__53190),
            .I(N__53187));
    Span4Mux_h I__11070 (
            .O(N__53187),
            .I(N__53184));
    Odrv4 I__11069 (
            .O(N__53184),
            .I(\c0.n3_adj_4394 ));
    CascadeMux I__11068 (
            .O(N__53181),
            .I(N__53177));
    InMux I__11067 (
            .O(N__53180),
            .I(N__53174));
    InMux I__11066 (
            .O(N__53177),
            .I(N__53171));
    LocalMux I__11065 (
            .O(N__53174),
            .I(N__53165));
    LocalMux I__11064 (
            .O(N__53171),
            .I(N__53165));
    InMux I__11063 (
            .O(N__53170),
            .I(N__53162));
    Span4Mux_v I__11062 (
            .O(N__53165),
            .I(N__53159));
    LocalMux I__11061 (
            .O(N__53162),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv4 I__11060 (
            .O(N__53159),
            .I(\c0.FRAME_MATCHER_i_19 ));
    InMux I__11059 (
            .O(N__53154),
            .I(bfn_19_20_0_));
    SRMux I__11058 (
            .O(N__53151),
            .I(N__53148));
    LocalMux I__11057 (
            .O(N__53148),
            .I(N__53145));
    Span4Mux_v I__11056 (
            .O(N__53145),
            .I(N__53142));
    Span4Mux_h I__11055 (
            .O(N__53142),
            .I(N__53139));
    Odrv4 I__11054 (
            .O(N__53139),
            .I(\c0.n3_adj_4398 ));
    InMux I__11053 (
            .O(N__53136),
            .I(N__53133));
    LocalMux I__11052 (
            .O(N__53133),
            .I(N__53129));
    InMux I__11051 (
            .O(N__53132),
            .I(N__53126));
    Span4Mux_v I__11050 (
            .O(N__53129),
            .I(N__53120));
    LocalMux I__11049 (
            .O(N__53126),
            .I(N__53120));
    InMux I__11048 (
            .O(N__53125),
            .I(N__53117));
    Sp12to4 I__11047 (
            .O(N__53120),
            .I(N__53114));
    LocalMux I__11046 (
            .O(N__53117),
            .I(\c0.FRAME_MATCHER_i_20 ));
    Odrv12 I__11045 (
            .O(N__53114),
            .I(\c0.FRAME_MATCHER_i_20 ));
    InMux I__11044 (
            .O(N__53109),
            .I(bfn_19_21_0_));
    InMux I__11043 (
            .O(N__53106),
            .I(bfn_19_19_0_));
    CascadeMux I__11042 (
            .O(N__53103),
            .I(N__53100));
    InMux I__11041 (
            .O(N__53100),
            .I(N__53096));
    InMux I__11040 (
            .O(N__53099),
            .I(N__53093));
    LocalMux I__11039 (
            .O(N__53096),
            .I(N__53090));
    LocalMux I__11038 (
            .O(N__53093),
            .I(N__53084));
    Span4Mux_v I__11037 (
            .O(N__53090),
            .I(N__53084));
    InMux I__11036 (
            .O(N__53089),
            .I(N__53081));
    Span4Mux_v I__11035 (
            .O(N__53084),
            .I(N__53078));
    LocalMux I__11034 (
            .O(N__53081),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__11033 (
            .O(N__53078),
            .I(\c0.FRAME_MATCHER_i_17 ));
    InMux I__11032 (
            .O(N__53073),
            .I(bfn_19_18_0_));
    SRMux I__11031 (
            .O(N__53070),
            .I(N__53067));
    LocalMux I__11030 (
            .O(N__53067),
            .I(N__53064));
    Span4Mux_v I__11029 (
            .O(N__53064),
            .I(N__53061));
    Odrv4 I__11028 (
            .O(N__53061),
            .I(\c0.n3_adj_4402 ));
    CascadeMux I__11027 (
            .O(N__53058),
            .I(N__53055));
    InMux I__11026 (
            .O(N__53055),
            .I(N__53051));
    InMux I__11025 (
            .O(N__53054),
            .I(N__53048));
    LocalMux I__11024 (
            .O(N__53051),
            .I(N__53045));
    LocalMux I__11023 (
            .O(N__53048),
            .I(N__53042));
    Span4Mux_h I__11022 (
            .O(N__53045),
            .I(N__53039));
    Span4Mux_h I__11021 (
            .O(N__53042),
            .I(N__53033));
    Span4Mux_v I__11020 (
            .O(N__53039),
            .I(N__53033));
    InMux I__11019 (
            .O(N__53038),
            .I(N__53030));
    Span4Mux_v I__11018 (
            .O(N__53033),
            .I(N__53027));
    LocalMux I__11017 (
            .O(N__53030),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__11016 (
            .O(N__53027),
            .I(\c0.FRAME_MATCHER_i_16 ));
    InMux I__11015 (
            .O(N__53022),
            .I(bfn_19_17_0_));
    SRMux I__11014 (
            .O(N__53019),
            .I(N__53016));
    LocalMux I__11013 (
            .O(N__53016),
            .I(N__53013));
    Span4Mux_h I__11012 (
            .O(N__53013),
            .I(N__53010));
    Odrv4 I__11011 (
            .O(N__53010),
            .I(\c0.n3_adj_4404 ));
    InMux I__11010 (
            .O(N__53007),
            .I(N__53003));
    InMux I__11009 (
            .O(N__53006),
            .I(N__53000));
    LocalMux I__11008 (
            .O(N__53003),
            .I(N__52997));
    LocalMux I__11007 (
            .O(N__53000),
            .I(N__52993));
    Span4Mux_v I__11006 (
            .O(N__52997),
            .I(N__52990));
    InMux I__11005 (
            .O(N__52996),
            .I(N__52987));
    Span12Mux_h I__11004 (
            .O(N__52993),
            .I(N__52982));
    Sp12to4 I__11003 (
            .O(N__52990),
            .I(N__52982));
    LocalMux I__11002 (
            .O(N__52987),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv12 I__11001 (
            .O(N__52982),
            .I(\c0.FRAME_MATCHER_i_15 ));
    InMux I__11000 (
            .O(N__52977),
            .I(bfn_19_16_0_));
    SRMux I__10999 (
            .O(N__52974),
            .I(N__52971));
    LocalMux I__10998 (
            .O(N__52971),
            .I(N__52968));
    Span4Mux_h I__10997 (
            .O(N__52968),
            .I(N__52965));
    Span4Mux_v I__10996 (
            .O(N__52965),
            .I(N__52962));
    Odrv4 I__10995 (
            .O(N__52962),
            .I(\c0.n3_adj_4406 ));
    CascadeMux I__10994 (
            .O(N__52959),
            .I(N__52956));
    InMux I__10993 (
            .O(N__52956),
            .I(N__52952));
    InMux I__10992 (
            .O(N__52955),
            .I(N__52949));
    LocalMux I__10991 (
            .O(N__52952),
            .I(N__52946));
    LocalMux I__10990 (
            .O(N__52949),
            .I(N__52943));
    Sp12to4 I__10989 (
            .O(N__52946),
            .I(N__52939));
    Span4Mux_v I__10988 (
            .O(N__52943),
            .I(N__52936));
    InMux I__10987 (
            .O(N__52942),
            .I(N__52933));
    Span12Mux_s9_v I__10986 (
            .O(N__52939),
            .I(N__52930));
    Odrv4 I__10985 (
            .O(N__52936),
            .I(\c0.FRAME_MATCHER_i_14 ));
    LocalMux I__10984 (
            .O(N__52933),
            .I(\c0.FRAME_MATCHER_i_14 ));
    Odrv12 I__10983 (
            .O(N__52930),
            .I(\c0.FRAME_MATCHER_i_14 ));
    InMux I__10982 (
            .O(N__52923),
            .I(bfn_19_15_0_));
    SRMux I__10981 (
            .O(N__52920),
            .I(N__52917));
    LocalMux I__10980 (
            .O(N__52917),
            .I(N__52914));
    Span4Mux_v I__10979 (
            .O(N__52914),
            .I(N__52911));
    Odrv4 I__10978 (
            .O(N__52911),
            .I(\c0.n3_adj_4408 ));
    InMux I__10977 (
            .O(N__52908),
            .I(bfn_19_14_0_));
    InMux I__10976 (
            .O(N__52905),
            .I(N__52901));
    InMux I__10975 (
            .O(N__52904),
            .I(N__52898));
    LocalMux I__10974 (
            .O(N__52901),
            .I(N__52895));
    LocalMux I__10973 (
            .O(N__52898),
            .I(N__52892));
    Sp12to4 I__10972 (
            .O(N__52895),
            .I(N__52886));
    Sp12to4 I__10971 (
            .O(N__52892),
            .I(N__52886));
    InMux I__10970 (
            .O(N__52891),
            .I(N__52883));
    Span12Mux_s11_v I__10969 (
            .O(N__52886),
            .I(N__52880));
    LocalMux I__10968 (
            .O(N__52883),
            .I(\c0.FRAME_MATCHER_i_12 ));
    Odrv12 I__10967 (
            .O(N__52880),
            .I(\c0.FRAME_MATCHER_i_12 ));
    InMux I__10966 (
            .O(N__52875),
            .I(bfn_19_13_0_));
    SRMux I__10965 (
            .O(N__52872),
            .I(N__52869));
    LocalMux I__10964 (
            .O(N__52869),
            .I(N__52866));
    Span4Mux_v I__10963 (
            .O(N__52866),
            .I(N__52863));
    Span4Mux_v I__10962 (
            .O(N__52863),
            .I(N__52860));
    Span4Mux_v I__10961 (
            .O(N__52860),
            .I(N__52857));
    Odrv4 I__10960 (
            .O(N__52857),
            .I(\c0.n3_adj_4412 ));
    SRMux I__10959 (
            .O(N__52854),
            .I(N__52851));
    LocalMux I__10958 (
            .O(N__52851),
            .I(N__52848));
    Span4Mux_v I__10957 (
            .O(N__52848),
            .I(N__52845));
    Span4Mux_v I__10956 (
            .O(N__52845),
            .I(N__52842));
    Span4Mux_v I__10955 (
            .O(N__52842),
            .I(N__52839));
    Odrv4 I__10954 (
            .O(N__52839),
            .I(\c0.n3_adj_4416 ));
    InMux I__10953 (
            .O(N__52836),
            .I(N__52832));
    InMux I__10952 (
            .O(N__52835),
            .I(N__52829));
    LocalMux I__10951 (
            .O(N__52832),
            .I(N__52826));
    LocalMux I__10950 (
            .O(N__52829),
            .I(N__52823));
    Span4Mux_h I__10949 (
            .O(N__52826),
            .I(N__52820));
    Span4Mux_h I__10948 (
            .O(N__52823),
            .I(N__52817));
    Sp12to4 I__10947 (
            .O(N__52820),
            .I(N__52811));
    Sp12to4 I__10946 (
            .O(N__52817),
            .I(N__52811));
    InMux I__10945 (
            .O(N__52816),
            .I(N__52808));
    Span12Mux_v I__10944 (
            .O(N__52811),
            .I(N__52805));
    LocalMux I__10943 (
            .O(N__52808),
            .I(\c0.FRAME_MATCHER_i_11 ));
    Odrv12 I__10942 (
            .O(N__52805),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__10941 (
            .O(N__52800),
            .I(bfn_19_12_0_));
    SRMux I__10940 (
            .O(N__52797),
            .I(N__52794));
    LocalMux I__10939 (
            .O(N__52794),
            .I(N__52791));
    Span4Mux_h I__10938 (
            .O(N__52791),
            .I(N__52788));
    Span4Mux_v I__10937 (
            .O(N__52788),
            .I(N__52785));
    Span4Mux_v I__10936 (
            .O(N__52785),
            .I(N__52782));
    Span4Mux_h I__10935 (
            .O(N__52782),
            .I(N__52779));
    Odrv4 I__10934 (
            .O(N__52779),
            .I(\c0.n3_adj_4414 ));
    InMux I__10933 (
            .O(N__52776),
            .I(N__52773));
    LocalMux I__10932 (
            .O(N__52773),
            .I(N__52770));
    Span4Mux_h I__10931 (
            .O(N__52770),
            .I(N__52766));
    InMux I__10930 (
            .O(N__52769),
            .I(N__52763));
    Span4Mux_v I__10929 (
            .O(N__52766),
            .I(N__52760));
    LocalMux I__10928 (
            .O(N__52763),
            .I(N__52757));
    Sp12to4 I__10927 (
            .O(N__52760),
            .I(N__52751));
    Span12Mux_h I__10926 (
            .O(N__52757),
            .I(N__52751));
    InMux I__10925 (
            .O(N__52756),
            .I(N__52748));
    Span12Mux_v I__10924 (
            .O(N__52751),
            .I(N__52745));
    LocalMux I__10923 (
            .O(N__52748),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv12 I__10922 (
            .O(N__52745),
            .I(\c0.FRAME_MATCHER_i_9 ));
    InMux I__10921 (
            .O(N__52740),
            .I(bfn_19_10_0_));
    SRMux I__10920 (
            .O(N__52737),
            .I(N__52734));
    LocalMux I__10919 (
            .O(N__52734),
            .I(N__52731));
    Span4Mux_v I__10918 (
            .O(N__52731),
            .I(N__52728));
    Span4Mux_v I__10917 (
            .O(N__52728),
            .I(N__52725));
    Odrv4 I__10916 (
            .O(N__52725),
            .I(\c0.n3_adj_4418 ));
    InMux I__10915 (
            .O(N__52722),
            .I(N__52716));
    InMux I__10914 (
            .O(N__52721),
            .I(N__52716));
    LocalMux I__10913 (
            .O(N__52716),
            .I(N__52713));
    Sp12to4 I__10912 (
            .O(N__52713),
            .I(N__52709));
    InMux I__10911 (
            .O(N__52712),
            .I(N__52706));
    Span12Mux_v I__10910 (
            .O(N__52709),
            .I(N__52703));
    LocalMux I__10909 (
            .O(N__52706),
            .I(\c0.FRAME_MATCHER_i_10 ));
    Odrv12 I__10908 (
            .O(N__52703),
            .I(\c0.FRAME_MATCHER_i_10 ));
    InMux I__10907 (
            .O(N__52698),
            .I(bfn_19_11_0_));
    InMux I__10906 (
            .O(N__52695),
            .I(N__52691));
    InMux I__10905 (
            .O(N__52694),
            .I(N__52688));
    LocalMux I__10904 (
            .O(N__52691),
            .I(N__52685));
    LocalMux I__10903 (
            .O(N__52688),
            .I(N__52682));
    Span4Mux_v I__10902 (
            .O(N__52685),
            .I(N__52679));
    Span4Mux_v I__10901 (
            .O(N__52682),
            .I(N__52676));
    Span4Mux_h I__10900 (
            .O(N__52679),
            .I(N__52673));
    Span4Mux_v I__10899 (
            .O(N__52676),
            .I(N__52670));
    Span4Mux_v I__10898 (
            .O(N__52673),
            .I(N__52666));
    Sp12to4 I__10897 (
            .O(N__52670),
            .I(N__52663));
    InMux I__10896 (
            .O(N__52669),
            .I(N__52660));
    Odrv4 I__10895 (
            .O(N__52666),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv12 I__10894 (
            .O(N__52663),
            .I(\c0.FRAME_MATCHER_i_8 ));
    LocalMux I__10893 (
            .O(N__52660),
            .I(\c0.FRAME_MATCHER_i_8 ));
    InMux I__10892 (
            .O(N__52653),
            .I(bfn_19_9_0_));
    SRMux I__10891 (
            .O(N__52650),
            .I(N__52647));
    LocalMux I__10890 (
            .O(N__52647),
            .I(N__52644));
    Span4Mux_h I__10889 (
            .O(N__52644),
            .I(N__52641));
    Span4Mux_h I__10888 (
            .O(N__52641),
            .I(N__52638));
    Span4Mux_v I__10887 (
            .O(N__52638),
            .I(N__52635));
    Odrv4 I__10886 (
            .O(N__52635),
            .I(\c0.n3_adj_4420 ));
    InMux I__10885 (
            .O(N__52632),
            .I(N__52629));
    LocalMux I__10884 (
            .O(N__52629),
            .I(N__52625));
    InMux I__10883 (
            .O(N__52628),
            .I(N__52622));
    Span4Mux_h I__10882 (
            .O(N__52625),
            .I(N__52619));
    LocalMux I__10881 (
            .O(N__52622),
            .I(N__52616));
    Sp12to4 I__10880 (
            .O(N__52619),
            .I(N__52610));
    Sp12to4 I__10879 (
            .O(N__52616),
            .I(N__52610));
    InMux I__10878 (
            .O(N__52615),
            .I(N__52607));
    Span12Mux_v I__10877 (
            .O(N__52610),
            .I(N__52604));
    LocalMux I__10876 (
            .O(N__52607),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv12 I__10875 (
            .O(N__52604),
            .I(\c0.FRAME_MATCHER_i_7 ));
    InMux I__10874 (
            .O(N__52599),
            .I(bfn_19_8_0_));
    SRMux I__10873 (
            .O(N__52596),
            .I(N__52593));
    LocalMux I__10872 (
            .O(N__52593),
            .I(N__52590));
    Span4Mux_v I__10871 (
            .O(N__52590),
            .I(N__52587));
    Span4Mux_v I__10870 (
            .O(N__52587),
            .I(N__52584));
    Span4Mux_v I__10869 (
            .O(N__52584),
            .I(N__52581));
    Span4Mux_h I__10868 (
            .O(N__52581),
            .I(N__52578));
    Odrv4 I__10867 (
            .O(N__52578),
            .I(\c0.n3_adj_4422 ));
    InMux I__10866 (
            .O(N__52575),
            .I(N__52572));
    LocalMux I__10865 (
            .O(N__52572),
            .I(N__52569));
    Span4Mux_v I__10864 (
            .O(N__52569),
            .I(N__52565));
    InMux I__10863 (
            .O(N__52568),
            .I(N__52562));
    Span4Mux_v I__10862 (
            .O(N__52565),
            .I(N__52556));
    LocalMux I__10861 (
            .O(N__52562),
            .I(N__52556));
    InMux I__10860 (
            .O(N__52561),
            .I(N__52553));
    Span4Mux_v I__10859 (
            .O(N__52556),
            .I(N__52549));
    LocalMux I__10858 (
            .O(N__52553),
            .I(N__52546));
    InMux I__10857 (
            .O(N__52552),
            .I(N__52543));
    Span4Mux_v I__10856 (
            .O(N__52549),
            .I(N__52540));
    Span4Mux_h I__10855 (
            .O(N__52546),
            .I(N__52537));
    LocalMux I__10854 (
            .O(N__52543),
            .I(N__52534));
    Span4Mux_v I__10853 (
            .O(N__52540),
            .I(N__52531));
    Sp12to4 I__10852 (
            .O(N__52537),
            .I(N__52526));
    Sp12to4 I__10851 (
            .O(N__52534),
            .I(N__52526));
    Span4Mux_h I__10850 (
            .O(N__52531),
            .I(N__52522));
    Span12Mux_v I__10849 (
            .O(N__52526),
            .I(N__52519));
    InMux I__10848 (
            .O(N__52525),
            .I(N__52516));
    Odrv4 I__10847 (
            .O(N__52522),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv12 I__10846 (
            .O(N__52519),
            .I(\c0.FRAME_MATCHER_i_6 ));
    LocalMux I__10845 (
            .O(N__52516),
            .I(\c0.FRAME_MATCHER_i_6 ));
    InMux I__10844 (
            .O(N__52509),
            .I(bfn_19_7_0_));
    SRMux I__10843 (
            .O(N__52506),
            .I(N__52503));
    LocalMux I__10842 (
            .O(N__52503),
            .I(N__52500));
    Span4Mux_v I__10841 (
            .O(N__52500),
            .I(N__52497));
    Span4Mux_v I__10840 (
            .O(N__52497),
            .I(N__52494));
    Sp12to4 I__10839 (
            .O(N__52494),
            .I(N__52491));
    Span12Mux_h I__10838 (
            .O(N__52491),
            .I(N__52488));
    Odrv12 I__10837 (
            .O(N__52488),
            .I(\c0.n3_adj_4424 ));
    InMux I__10836 (
            .O(N__52485),
            .I(N__52482));
    LocalMux I__10835 (
            .O(N__52482),
            .I(N__52477));
    InMux I__10834 (
            .O(N__52481),
            .I(N__52474));
    InMux I__10833 (
            .O(N__52480),
            .I(N__52471));
    Span4Mux_v I__10832 (
            .O(N__52477),
            .I(N__52468));
    LocalMux I__10831 (
            .O(N__52474),
            .I(N__52465));
    LocalMux I__10830 (
            .O(N__52471),
            .I(N__52462));
    Sp12to4 I__10829 (
            .O(N__52468),
            .I(N__52459));
    Span4Mux_h I__10828 (
            .O(N__52465),
            .I(N__52456));
    Span12Mux_h I__10827 (
            .O(N__52462),
            .I(N__52451));
    Span12Mux_h I__10826 (
            .O(N__52459),
            .I(N__52446));
    Sp12to4 I__10825 (
            .O(N__52456),
            .I(N__52446));
    InMux I__10824 (
            .O(N__52455),
            .I(N__52443));
    InMux I__10823 (
            .O(N__52454),
            .I(N__52440));
    Span12Mux_v I__10822 (
            .O(N__52451),
            .I(N__52437));
    Span12Mux_v I__10821 (
            .O(N__52446),
            .I(N__52434));
    LocalMux I__10820 (
            .O(N__52443),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__10819 (
            .O(N__52440),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv12 I__10818 (
            .O(N__52437),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv12 I__10817 (
            .O(N__52434),
            .I(\c0.FRAME_MATCHER_i_5 ));
    InMux I__10816 (
            .O(N__52425),
            .I(bfn_19_6_0_));
    SRMux I__10815 (
            .O(N__52422),
            .I(N__52419));
    LocalMux I__10814 (
            .O(N__52419),
            .I(N__52416));
    Span4Mux_v I__10813 (
            .O(N__52416),
            .I(N__52413));
    Odrv4 I__10812 (
            .O(N__52413),
            .I(\c0.n3_adj_4426 ));
    InMux I__10811 (
            .O(N__52410),
            .I(N__52404));
    InMux I__10810 (
            .O(N__52409),
            .I(N__52401));
    InMux I__10809 (
            .O(N__52408),
            .I(N__52398));
    InMux I__10808 (
            .O(N__52407),
            .I(N__52395));
    LocalMux I__10807 (
            .O(N__52404),
            .I(N__52392));
    LocalMux I__10806 (
            .O(N__52401),
            .I(N__52389));
    LocalMux I__10805 (
            .O(N__52398),
            .I(N__52384));
    LocalMux I__10804 (
            .O(N__52395),
            .I(N__52384));
    Span4Mux_h I__10803 (
            .O(N__52392),
            .I(N__52381));
    Span4Mux_h I__10802 (
            .O(N__52389),
            .I(N__52378));
    Span4Mux_h I__10801 (
            .O(N__52384),
            .I(N__52375));
    Span4Mux_v I__10800 (
            .O(N__52381),
            .I(N__52371));
    Sp12to4 I__10799 (
            .O(N__52378),
            .I(N__52366));
    Sp12to4 I__10798 (
            .O(N__52375),
            .I(N__52366));
    InMux I__10797 (
            .O(N__52374),
            .I(N__52363));
    Span4Mux_v I__10796 (
            .O(N__52371),
            .I(N__52359));
    Span12Mux_s7_v I__10795 (
            .O(N__52366),
            .I(N__52356));
    LocalMux I__10794 (
            .O(N__52363),
            .I(N__52353));
    InMux I__10793 (
            .O(N__52362),
            .I(N__52350));
    Span4Mux_v I__10792 (
            .O(N__52359),
            .I(N__52347));
    Span12Mux_v I__10791 (
            .O(N__52356),
            .I(N__52344));
    Odrv4 I__10790 (
            .O(N__52353),
            .I(\c0.FRAME_MATCHER_i_4 ));
    LocalMux I__10789 (
            .O(N__52350),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv4 I__10788 (
            .O(N__52347),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv12 I__10787 (
            .O(N__52344),
            .I(\c0.FRAME_MATCHER_i_4 ));
    InMux I__10786 (
            .O(N__52335),
            .I(bfn_19_5_0_));
    SRMux I__10785 (
            .O(N__52332),
            .I(N__52329));
    LocalMux I__10784 (
            .O(N__52329),
            .I(N__52326));
    Span4Mux_h I__10783 (
            .O(N__52326),
            .I(N__52323));
    Odrv4 I__10782 (
            .O(N__52323),
            .I(\c0.n3_adj_4428 ));
    InMux I__10781 (
            .O(N__52320),
            .I(bfn_19_4_0_));
    SRMux I__10780 (
            .O(N__52317),
            .I(N__52314));
    LocalMux I__10779 (
            .O(N__52314),
            .I(N__52311));
    Span4Mux_h I__10778 (
            .O(N__52311),
            .I(N__52308));
    Span4Mux_v I__10777 (
            .O(N__52308),
            .I(N__52305));
    Odrv4 I__10776 (
            .O(N__52305),
            .I(\c0.n3_adj_4434 ));
    InMux I__10775 (
            .O(N__52302),
            .I(bfn_19_3_0_));
    SRMux I__10774 (
            .O(N__52299),
            .I(N__52296));
    LocalMux I__10773 (
            .O(N__52296),
            .I(N__52293));
    Span4Mux_v I__10772 (
            .O(N__52293),
            .I(N__52290));
    Span4Mux_v I__10771 (
            .O(N__52290),
            .I(N__52287));
    Odrv4 I__10770 (
            .O(N__52287),
            .I(\c0.n3_adj_4432 ));
    CascadeMux I__10769 (
            .O(N__52284),
            .I(N__52281));
    InMux I__10768 (
            .O(N__52281),
            .I(N__52278));
    LocalMux I__10767 (
            .O(N__52278),
            .I(\c0.n161 ));
    InMux I__10766 (
            .O(N__52275),
            .I(bfn_19_2_0_));
    InMux I__10765 (
            .O(N__52272),
            .I(N__52269));
    LocalMux I__10764 (
            .O(N__52269),
            .I(\c0.n41_adj_4292 ));
    CascadeMux I__10763 (
            .O(N__52266),
            .I(\c0.n42_adj_4272_cascade_ ));
    InMux I__10762 (
            .O(N__52263),
            .I(N__52260));
    LocalMux I__10761 (
            .O(N__52260),
            .I(\c0.n44_adj_4270 ));
    InMux I__10760 (
            .O(N__52257),
            .I(N__52254));
    LocalMux I__10759 (
            .O(N__52254),
            .I(\c0.n50_adj_4296 ));
    InMux I__10758 (
            .O(N__52251),
            .I(N__52248));
    LocalMux I__10757 (
            .O(N__52248),
            .I(\c0.n43_adj_4275 ));
    CascadeMux I__10756 (
            .O(N__52245),
            .I(N__52242));
    InMux I__10755 (
            .O(N__52242),
            .I(N__52238));
    CascadeMux I__10754 (
            .O(N__52241),
            .I(N__52235));
    LocalMux I__10753 (
            .O(N__52238),
            .I(N__52232));
    InMux I__10752 (
            .O(N__52235),
            .I(N__52229));
    Span4Mux_v I__10751 (
            .O(N__52232),
            .I(N__52226));
    LocalMux I__10750 (
            .O(N__52229),
            .I(N__52223));
    Sp12to4 I__10749 (
            .O(N__52226),
            .I(N__52220));
    Odrv4 I__10748 (
            .O(N__52223),
            .I(\c0.data_in_frame_28_7 ));
    Odrv12 I__10747 (
            .O(N__52220),
            .I(\c0.data_in_frame_28_7 ));
    CascadeMux I__10746 (
            .O(N__52215),
            .I(N__52212));
    InMux I__10745 (
            .O(N__52212),
            .I(N__52209));
    LocalMux I__10744 (
            .O(N__52209),
            .I(\c0.n45_adj_4298 ));
    InMux I__10743 (
            .O(N__52206),
            .I(N__52201));
    InMux I__10742 (
            .O(N__52205),
            .I(N__52198));
    CascadeMux I__10741 (
            .O(N__52204),
            .I(N__52195));
    LocalMux I__10740 (
            .O(N__52201),
            .I(N__52192));
    LocalMux I__10739 (
            .O(N__52198),
            .I(N__52188));
    InMux I__10738 (
            .O(N__52195),
            .I(N__52185));
    Span4Mux_h I__10737 (
            .O(N__52192),
            .I(N__52182));
    InMux I__10736 (
            .O(N__52191),
            .I(N__52179));
    Span4Mux_v I__10735 (
            .O(N__52188),
            .I(N__52176));
    LocalMux I__10734 (
            .O(N__52185),
            .I(\c0.data_in_frame_25_3 ));
    Odrv4 I__10733 (
            .O(N__52182),
            .I(\c0.data_in_frame_25_3 ));
    LocalMux I__10732 (
            .O(N__52179),
            .I(\c0.data_in_frame_25_3 ));
    Odrv4 I__10731 (
            .O(N__52176),
            .I(\c0.data_in_frame_25_3 ));
    InMux I__10730 (
            .O(N__52167),
            .I(N__52162));
    InMux I__10729 (
            .O(N__52166),
            .I(N__52159));
    CascadeMux I__10728 (
            .O(N__52165),
            .I(N__52156));
    LocalMux I__10727 (
            .O(N__52162),
            .I(N__52150));
    LocalMux I__10726 (
            .O(N__52159),
            .I(N__52150));
    InMux I__10725 (
            .O(N__52156),
            .I(N__52145));
    InMux I__10724 (
            .O(N__52155),
            .I(N__52145));
    Odrv12 I__10723 (
            .O(N__52150),
            .I(\c0.data_in_frame_25_2 ));
    LocalMux I__10722 (
            .O(N__52145),
            .I(\c0.data_in_frame_25_2 ));
    InMux I__10721 (
            .O(N__52140),
            .I(N__52137));
    LocalMux I__10720 (
            .O(N__52137),
            .I(\c0.n40_adj_4294 ));
    InMux I__10719 (
            .O(N__52134),
            .I(N__52129));
    InMux I__10718 (
            .O(N__52133),
            .I(N__52124));
    InMux I__10717 (
            .O(N__52132),
            .I(N__52124));
    LocalMux I__10716 (
            .O(N__52129),
            .I(N__52121));
    LocalMux I__10715 (
            .O(N__52124),
            .I(N__52118));
    Odrv4 I__10714 (
            .O(N__52121),
            .I(\c0.n5_adj_4349 ));
    Odrv4 I__10713 (
            .O(N__52118),
            .I(\c0.n5_adj_4349 ));
    CascadeMux I__10712 (
            .O(N__52113),
            .I(\c0.n10_adj_4371_cascade_ ));
    InMux I__10711 (
            .O(N__52110),
            .I(N__52107));
    LocalMux I__10710 (
            .O(N__52107),
            .I(\c0.n12_adj_4372 ));
    CascadeMux I__10709 (
            .O(N__52104),
            .I(\c0.n12_adj_4671_cascade_ ));
    CascadeMux I__10708 (
            .O(N__52101),
            .I(N__52098));
    InMux I__10707 (
            .O(N__52098),
            .I(N__52094));
    CascadeMux I__10706 (
            .O(N__52097),
            .I(N__52091));
    LocalMux I__10705 (
            .O(N__52094),
            .I(N__52087));
    InMux I__10704 (
            .O(N__52091),
            .I(N__52084));
    InMux I__10703 (
            .O(N__52090),
            .I(N__52081));
    Span4Mux_v I__10702 (
            .O(N__52087),
            .I(N__52078));
    LocalMux I__10701 (
            .O(N__52084),
            .I(N__52075));
    LocalMux I__10700 (
            .O(N__52081),
            .I(N__52072));
    Sp12to4 I__10699 (
            .O(N__52078),
            .I(N__52068));
    Span4Mux_h I__10698 (
            .O(N__52075),
            .I(N__52065));
    Span4Mux_h I__10697 (
            .O(N__52072),
            .I(N__52062));
    CascadeMux I__10696 (
            .O(N__52071),
            .I(N__52059));
    Span12Mux_h I__10695 (
            .O(N__52068),
            .I(N__52056));
    Sp12to4 I__10694 (
            .O(N__52065),
            .I(N__52051));
    Sp12to4 I__10693 (
            .O(N__52062),
            .I(N__52051));
    InMux I__10692 (
            .O(N__52059),
            .I(N__52048));
    Span12Mux_v I__10691 (
            .O(N__52056),
            .I(N__52045));
    Span12Mux_v I__10690 (
            .O(N__52051),
            .I(N__52042));
    LocalMux I__10689 (
            .O(N__52048),
            .I(\c0.data_in_frame_24_7 ));
    Odrv12 I__10688 (
            .O(N__52045),
            .I(\c0.data_in_frame_24_7 ));
    Odrv12 I__10687 (
            .O(N__52042),
            .I(\c0.data_in_frame_24_7 ));
    InMux I__10686 (
            .O(N__52035),
            .I(N__52032));
    LocalMux I__10685 (
            .O(N__52032),
            .I(\c0.n25467 ));
    InMux I__10684 (
            .O(N__52029),
            .I(N__52025));
    InMux I__10683 (
            .O(N__52028),
            .I(N__52022));
    LocalMux I__10682 (
            .O(N__52025),
            .I(\c0.n24098 ));
    LocalMux I__10681 (
            .O(N__52022),
            .I(\c0.n24098 ));
    CascadeMux I__10680 (
            .O(N__52017),
            .I(N__52014));
    InMux I__10679 (
            .O(N__52014),
            .I(N__52010));
    InMux I__10678 (
            .O(N__52013),
            .I(N__52007));
    LocalMux I__10677 (
            .O(N__52010),
            .I(N__52004));
    LocalMux I__10676 (
            .O(N__52007),
            .I(\c0.data_in_frame_29_4 ));
    Odrv12 I__10675 (
            .O(N__52004),
            .I(\c0.data_in_frame_29_4 ));
    InMux I__10674 (
            .O(N__51999),
            .I(N__51995));
    InMux I__10673 (
            .O(N__51998),
            .I(N__51992));
    LocalMux I__10672 (
            .O(N__51995),
            .I(N__51987));
    LocalMux I__10671 (
            .O(N__51992),
            .I(N__51987));
    Odrv4 I__10670 (
            .O(N__51987),
            .I(\c0.n23533 ));
    CascadeMux I__10669 (
            .O(N__51984),
            .I(N__51981));
    InMux I__10668 (
            .O(N__51981),
            .I(N__51978));
    LocalMux I__10667 (
            .O(N__51978),
            .I(N__51975));
    Span4Mux_v I__10666 (
            .O(N__51975),
            .I(N__51972));
    Odrv4 I__10665 (
            .O(N__51972),
            .I(\c0.n5_adj_4370 ));
    InMux I__10664 (
            .O(N__51969),
            .I(N__51966));
    LocalMux I__10663 (
            .O(N__51966),
            .I(N__51963));
    Odrv4 I__10662 (
            .O(N__51963),
            .I(\c0.n10_adj_4371 ));
    CascadeMux I__10661 (
            .O(N__51960),
            .I(\c0.n10_adj_4439_cascade_ ));
    InMux I__10660 (
            .O(N__51957),
            .I(N__51954));
    LocalMux I__10659 (
            .O(N__51954),
            .I(\c0.n20_adj_4441 ));
    CascadeMux I__10658 (
            .O(N__51951),
            .I(\c0.n13_adj_4442_cascade_ ));
    CascadeMux I__10657 (
            .O(N__51948),
            .I(\c0.n24528_cascade_ ));
    InMux I__10656 (
            .O(N__51945),
            .I(N__51940));
    InMux I__10655 (
            .O(N__51944),
            .I(N__51937));
    InMux I__10654 (
            .O(N__51943),
            .I(N__51934));
    LocalMux I__10653 (
            .O(N__51940),
            .I(N__51931));
    LocalMux I__10652 (
            .O(N__51937),
            .I(\c0.n23718 ));
    LocalMux I__10651 (
            .O(N__51934),
            .I(\c0.n23718 ));
    Odrv4 I__10650 (
            .O(N__51931),
            .I(\c0.n23718 ));
    InMux I__10649 (
            .O(N__51924),
            .I(N__51921));
    LocalMux I__10648 (
            .O(N__51921),
            .I(N__51918));
    Odrv4 I__10647 (
            .O(N__51918),
            .I(\c0.n12_adj_4506 ));
    InMux I__10646 (
            .O(N__51915),
            .I(N__51912));
    LocalMux I__10645 (
            .O(N__51912),
            .I(\c0.n20_adj_4512 ));
    InMux I__10644 (
            .O(N__51909),
            .I(N__51906));
    LocalMux I__10643 (
            .O(N__51906),
            .I(\c0.n24_adj_4509 ));
    InMux I__10642 (
            .O(N__51903),
            .I(N__51900));
    LocalMux I__10641 (
            .O(N__51900),
            .I(\c0.n22_adj_4507 ));
    InMux I__10640 (
            .O(N__51897),
            .I(N__51894));
    LocalMux I__10639 (
            .O(N__51894),
            .I(\c0.n23627 ));
    CascadeMux I__10638 (
            .O(N__51891),
            .I(\c0.n23627_cascade_ ));
    InMux I__10637 (
            .O(N__51888),
            .I(N__51882));
    InMux I__10636 (
            .O(N__51887),
            .I(N__51882));
    LocalMux I__10635 (
            .O(N__51882),
            .I(N__51878));
    InMux I__10634 (
            .O(N__51881),
            .I(N__51875));
    Odrv4 I__10633 (
            .O(N__51878),
            .I(\c0.n24528 ));
    LocalMux I__10632 (
            .O(N__51875),
            .I(\c0.n24528 ));
    InMux I__10631 (
            .O(N__51870),
            .I(N__51867));
    LocalMux I__10630 (
            .O(N__51867),
            .I(\c0.n10_adj_4575 ));
    InMux I__10629 (
            .O(N__51864),
            .I(N__51861));
    LocalMux I__10628 (
            .O(N__51861),
            .I(\c0.n23_adj_4598 ));
    CascadeMux I__10627 (
            .O(N__51858),
            .I(N__51855));
    InMux I__10626 (
            .O(N__51855),
            .I(N__51852));
    LocalMux I__10625 (
            .O(N__51852),
            .I(N__51849));
    Span4Mux_v I__10624 (
            .O(N__51849),
            .I(N__51846));
    Odrv4 I__10623 (
            .O(N__51846),
            .I(\c0.n4_adj_4352 ));
    InMux I__10622 (
            .O(N__51843),
            .I(N__51840));
    LocalMux I__10621 (
            .O(N__51840),
            .I(\c0.n23_adj_4353 ));
    CascadeMux I__10620 (
            .O(N__51837),
            .I(\c0.n23_adj_4353_cascade_ ));
    InMux I__10619 (
            .O(N__51834),
            .I(N__51828));
    InMux I__10618 (
            .O(N__51833),
            .I(N__51828));
    LocalMux I__10617 (
            .O(N__51828),
            .I(\c0.n15_adj_4344 ));
    InMux I__10616 (
            .O(N__51825),
            .I(N__51822));
    LocalMux I__10615 (
            .O(N__51822),
            .I(\c0.n21428 ));
    CascadeMux I__10614 (
            .O(N__51819),
            .I(\c0.n11_adj_4438_cascade_ ));
    InMux I__10613 (
            .O(N__51816),
            .I(N__51813));
    LocalMux I__10612 (
            .O(N__51813),
            .I(\c0.n16_adj_4437 ));
    InMux I__10611 (
            .O(N__51810),
            .I(N__51804));
    InMux I__10610 (
            .O(N__51809),
            .I(N__51804));
    LocalMux I__10609 (
            .O(N__51804),
            .I(\c0.n22420 ));
    CascadeMux I__10608 (
            .O(N__51801),
            .I(N__51797));
    CascadeMux I__10607 (
            .O(N__51800),
            .I(N__51794));
    InMux I__10606 (
            .O(N__51797),
            .I(N__51791));
    InMux I__10605 (
            .O(N__51794),
            .I(N__51788));
    LocalMux I__10604 (
            .O(N__51791),
            .I(N__51785));
    LocalMux I__10603 (
            .O(N__51788),
            .I(\c0.data_in_frame_28_0 ));
    Odrv4 I__10602 (
            .O(N__51785),
            .I(\c0.data_in_frame_28_0 ));
    InMux I__10601 (
            .O(N__51780),
            .I(N__51774));
    InMux I__10600 (
            .O(N__51779),
            .I(N__51770));
    InMux I__10599 (
            .O(N__51778),
            .I(N__51767));
    InMux I__10598 (
            .O(N__51777),
            .I(N__51764));
    LocalMux I__10597 (
            .O(N__51774),
            .I(N__51761));
    InMux I__10596 (
            .O(N__51773),
            .I(N__51758));
    LocalMux I__10595 (
            .O(N__51770),
            .I(N__51751));
    LocalMux I__10594 (
            .O(N__51767),
            .I(N__51751));
    LocalMux I__10593 (
            .O(N__51764),
            .I(N__51751));
    Span4Mux_v I__10592 (
            .O(N__51761),
            .I(N__51748));
    LocalMux I__10591 (
            .O(N__51758),
            .I(\c0.n21491 ));
    Odrv12 I__10590 (
            .O(N__51751),
            .I(\c0.n21491 ));
    Odrv4 I__10589 (
            .O(N__51748),
            .I(\c0.n21491 ));
    CascadeMux I__10588 (
            .O(N__51741),
            .I(\c0.n23187_cascade_ ));
    CascadeMux I__10587 (
            .O(N__51738),
            .I(\c0.n10_adj_4591_cascade_ ));
    InMux I__10586 (
            .O(N__51735),
            .I(N__51732));
    LocalMux I__10585 (
            .O(N__51732),
            .I(\c0.n10_adj_4591 ));
    InMux I__10584 (
            .O(N__51729),
            .I(N__51724));
    InMux I__10583 (
            .O(N__51728),
            .I(N__51719));
    InMux I__10582 (
            .O(N__51727),
            .I(N__51719));
    LocalMux I__10581 (
            .O(N__51724),
            .I(data_in_frame_21_2));
    LocalMux I__10580 (
            .O(N__51719),
            .I(data_in_frame_21_2));
    CascadeMux I__10579 (
            .O(N__51714),
            .I(\c0.n12_adj_4606_cascade_ ));
    CascadeMux I__10578 (
            .O(N__51711),
            .I(\c0.n21325_cascade_ ));
    InMux I__10577 (
            .O(N__51708),
            .I(N__51705));
    LocalMux I__10576 (
            .O(N__51705),
            .I(N__51702));
    Span4Mux_h I__10575 (
            .O(N__51702),
            .I(N__51699));
    Span4Mux_v I__10574 (
            .O(N__51699),
            .I(N__51696));
    Odrv4 I__10573 (
            .O(N__51696),
            .I(\c0.n24384 ));
    CascadeMux I__10572 (
            .O(N__51693),
            .I(\c0.n4_adj_4464_cascade_ ));
    CascadeMux I__10571 (
            .O(N__51690),
            .I(\c0.n21428_cascade_ ));
    InMux I__10570 (
            .O(N__51687),
            .I(N__51684));
    LocalMux I__10569 (
            .O(N__51684),
            .I(\c0.n24_adj_4593 ));
    InMux I__10568 (
            .O(N__51681),
            .I(N__51678));
    LocalMux I__10567 (
            .O(N__51678),
            .I(\c0.n154 ));
    CascadeMux I__10566 (
            .O(N__51675),
            .I(N__51672));
    InMux I__10565 (
            .O(N__51672),
            .I(N__51668));
    InMux I__10564 (
            .O(N__51671),
            .I(N__51665));
    LocalMux I__10563 (
            .O(N__51668),
            .I(N__51662));
    LocalMux I__10562 (
            .O(N__51665),
            .I(\c0.n15_adj_4301 ));
    Odrv4 I__10561 (
            .O(N__51662),
            .I(\c0.n15_adj_4301 ));
    InMux I__10560 (
            .O(N__51657),
            .I(N__51654));
    LocalMux I__10559 (
            .O(N__51654),
            .I(\c0.n21_adj_4605 ));
    CascadeMux I__10558 (
            .O(N__51651),
            .I(N__51648));
    InMux I__10557 (
            .O(N__51648),
            .I(N__51645));
    LocalMux I__10556 (
            .O(N__51645),
            .I(\c0.n19_adj_4604 ));
    InMux I__10555 (
            .O(N__51642),
            .I(N__51639));
    LocalMux I__10554 (
            .O(N__51639),
            .I(N__51636));
    Odrv12 I__10553 (
            .O(N__51636),
            .I(\c0.n16_adj_4256 ));
    InMux I__10552 (
            .O(N__51633),
            .I(N__51630));
    LocalMux I__10551 (
            .O(N__51630),
            .I(\c0.n22 ));
    InMux I__10550 (
            .O(N__51627),
            .I(N__51623));
    InMux I__10549 (
            .O(N__51626),
            .I(N__51620));
    LocalMux I__10548 (
            .O(N__51623),
            .I(N__51617));
    LocalMux I__10547 (
            .O(N__51620),
            .I(N__51614));
    Span4Mux_v I__10546 (
            .O(N__51617),
            .I(N__51610));
    Sp12to4 I__10545 (
            .O(N__51614),
            .I(N__51607));
    InMux I__10544 (
            .O(N__51613),
            .I(N__51604));
    Odrv4 I__10543 (
            .O(N__51610),
            .I(\c0.n13280 ));
    Odrv12 I__10542 (
            .O(N__51607),
            .I(\c0.n13280 ));
    LocalMux I__10541 (
            .O(N__51604),
            .I(\c0.n13280 ));
    CascadeMux I__10540 (
            .O(N__51597),
            .I(\c0.n13_cascade_ ));
    InMux I__10539 (
            .O(N__51594),
            .I(N__51591));
    LocalMux I__10538 (
            .O(N__51591),
            .I(N__51588));
    Odrv12 I__10537 (
            .O(N__51588),
            .I(\c0.n20_adj_4222 ));
    InMux I__10536 (
            .O(N__51585),
            .I(N__51582));
    LocalMux I__10535 (
            .O(N__51582),
            .I(N__51578));
    InMux I__10534 (
            .O(N__51581),
            .I(N__51575));
    Span4Mux_v I__10533 (
            .O(N__51578),
            .I(N__51568));
    LocalMux I__10532 (
            .O(N__51575),
            .I(N__51568));
    InMux I__10531 (
            .O(N__51574),
            .I(N__51565));
    InMux I__10530 (
            .O(N__51573),
            .I(N__51559));
    Span4Mux_v I__10529 (
            .O(N__51568),
            .I(N__51556));
    LocalMux I__10528 (
            .O(N__51565),
            .I(N__51553));
    InMux I__10527 (
            .O(N__51564),
            .I(N__51550));
    InMux I__10526 (
            .O(N__51563),
            .I(N__51547));
    InMux I__10525 (
            .O(N__51562),
            .I(N__51544));
    LocalMux I__10524 (
            .O(N__51559),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__10523 (
            .O(N__51556),
            .I(\c0.data_in_frame_3_5 ));
    Odrv12 I__10522 (
            .O(N__51553),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__10521 (
            .O(N__51550),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__10520 (
            .O(N__51547),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__10519 (
            .O(N__51544),
            .I(\c0.data_in_frame_3_5 ));
    CascadeMux I__10518 (
            .O(N__51531),
            .I(\c0.n22_adj_4223_cascade_ ));
    CascadeMux I__10517 (
            .O(N__51528),
            .I(\c0.n21_adj_4225_cascade_ ));
    CascadeMux I__10516 (
            .O(N__51525),
            .I(\c0.n10_adj_4277_cascade_ ));
    CascadeMux I__10515 (
            .O(N__51522),
            .I(N__51518));
    InMux I__10514 (
            .O(N__51521),
            .I(N__51510));
    InMux I__10513 (
            .O(N__51518),
            .I(N__51510));
    InMux I__10512 (
            .O(N__51517),
            .I(N__51510));
    LocalMux I__10511 (
            .O(N__51510),
            .I(\c0.n23116 ));
    InMux I__10510 (
            .O(N__51507),
            .I(N__51504));
    LocalMux I__10509 (
            .O(N__51504),
            .I(N__51501));
    Span4Mux_h I__10508 (
            .O(N__51501),
            .I(N__51498));
    Span4Mux_v I__10507 (
            .O(N__51498),
            .I(N__51495));
    Odrv4 I__10506 (
            .O(N__51495),
            .I(\c0.n128 ));
    CascadeMux I__10505 (
            .O(N__51492),
            .I(\c0.n129_cascade_ ));
    InMux I__10504 (
            .O(N__51489),
            .I(N__51486));
    LocalMux I__10503 (
            .O(N__51486),
            .I(\c0.n11_adj_4614 ));
    CascadeMux I__10502 (
            .O(N__51483),
            .I(\c0.n16_adj_4613_cascade_ ));
    InMux I__10501 (
            .O(N__51480),
            .I(N__51477));
    LocalMux I__10500 (
            .O(N__51477),
            .I(N__51474));
    Span4Mux_v I__10499 (
            .O(N__51474),
            .I(N__51471));
    Span4Mux_v I__10498 (
            .O(N__51471),
            .I(N__51468));
    Span4Mux_h I__10497 (
            .O(N__51468),
            .I(N__51461));
    InMux I__10496 (
            .O(N__51467),
            .I(N__51455));
    InMux I__10495 (
            .O(N__51466),
            .I(N__51455));
    CascadeMux I__10494 (
            .O(N__51465),
            .I(N__51452));
    CascadeMux I__10493 (
            .O(N__51464),
            .I(N__51449));
    Span4Mux_v I__10492 (
            .O(N__51461),
            .I(N__51443));
    InMux I__10491 (
            .O(N__51460),
            .I(N__51440));
    LocalMux I__10490 (
            .O(N__51455),
            .I(N__51436));
    InMux I__10489 (
            .O(N__51452),
            .I(N__51433));
    InMux I__10488 (
            .O(N__51449),
            .I(N__51428));
    InMux I__10487 (
            .O(N__51448),
            .I(N__51428));
    CascadeMux I__10486 (
            .O(N__51447),
            .I(N__51425));
    CascadeMux I__10485 (
            .O(N__51446),
            .I(N__51421));
    Span4Mux_h I__10484 (
            .O(N__51443),
            .I(N__51415));
    LocalMux I__10483 (
            .O(N__51440),
            .I(N__51412));
    InMux I__10482 (
            .O(N__51439),
            .I(N__51409));
    Span4Mux_v I__10481 (
            .O(N__51436),
            .I(N__51402));
    LocalMux I__10480 (
            .O(N__51433),
            .I(N__51402));
    LocalMux I__10479 (
            .O(N__51428),
            .I(N__51402));
    InMux I__10478 (
            .O(N__51425),
            .I(N__51397));
    InMux I__10477 (
            .O(N__51424),
            .I(N__51397));
    InMux I__10476 (
            .O(N__51421),
            .I(N__51390));
    InMux I__10475 (
            .O(N__51420),
            .I(N__51390));
    InMux I__10474 (
            .O(N__51419),
            .I(N__51390));
    InMux I__10473 (
            .O(N__51418),
            .I(N__51387));
    Odrv4 I__10472 (
            .O(N__51415),
            .I(data_in_frame_1_3));
    Odrv4 I__10471 (
            .O(N__51412),
            .I(data_in_frame_1_3));
    LocalMux I__10470 (
            .O(N__51409),
            .I(data_in_frame_1_3));
    Odrv4 I__10469 (
            .O(N__51402),
            .I(data_in_frame_1_3));
    LocalMux I__10468 (
            .O(N__51397),
            .I(data_in_frame_1_3));
    LocalMux I__10467 (
            .O(N__51390),
            .I(data_in_frame_1_3));
    LocalMux I__10466 (
            .O(N__51387),
            .I(data_in_frame_1_3));
    InMux I__10465 (
            .O(N__51372),
            .I(N__51369));
    LocalMux I__10464 (
            .O(N__51369),
            .I(N__51366));
    Odrv12 I__10463 (
            .O(N__51366),
            .I(\c0.n126 ));
    InMux I__10462 (
            .O(N__51363),
            .I(N__51360));
    LocalMux I__10461 (
            .O(N__51360),
            .I(\c0.n123 ));
    CascadeMux I__10460 (
            .O(N__51357),
            .I(\c0.n144_cascade_ ));
    InMux I__10459 (
            .O(N__51354),
            .I(N__51351));
    LocalMux I__10458 (
            .O(N__51351),
            .I(N__51348));
    Odrv4 I__10457 (
            .O(N__51348),
            .I(\c0.n7_adj_4221 ));
    InMux I__10456 (
            .O(N__51345),
            .I(N__51342));
    LocalMux I__10455 (
            .O(N__51342),
            .I(\c0.n16_adj_4641 ));
    CascadeMux I__10454 (
            .O(N__51339),
            .I(\c0.n23116_cascade_ ));
    InMux I__10453 (
            .O(N__51336),
            .I(N__51332));
    InMux I__10452 (
            .O(N__51335),
            .I(N__51329));
    LocalMux I__10451 (
            .O(N__51332),
            .I(N__51323));
    LocalMux I__10450 (
            .O(N__51329),
            .I(N__51323));
    InMux I__10449 (
            .O(N__51328),
            .I(N__51320));
    Span4Mux_v I__10448 (
            .O(N__51323),
            .I(N__51317));
    LocalMux I__10447 (
            .O(N__51320),
            .I(\c0.n7_adj_4337 ));
    Odrv4 I__10446 (
            .O(N__51317),
            .I(\c0.n7_adj_4337 ));
    CascadeMux I__10445 (
            .O(N__51312),
            .I(\c0.n38_adj_4573_cascade_ ));
    InMux I__10444 (
            .O(N__51309),
            .I(N__51306));
    LocalMux I__10443 (
            .O(N__51306),
            .I(N__51303));
    Odrv4 I__10442 (
            .O(N__51303),
            .I(\c0.n44_adj_4744 ));
    CascadeMux I__10441 (
            .O(N__51300),
            .I(\c0.n43_adj_4574_cascade_ ));
    InMux I__10440 (
            .O(N__51297),
            .I(N__51294));
    LocalMux I__10439 (
            .O(N__51294),
            .I(\c0.n41_adj_4745 ));
    InMux I__10438 (
            .O(N__51291),
            .I(N__51288));
    LocalMux I__10437 (
            .O(N__51288),
            .I(N__51285));
    Odrv4 I__10436 (
            .O(N__51285),
            .I(\c0.n24048 ));
    CascadeMux I__10435 (
            .O(N__51282),
            .I(\c0.n24048_cascade_ ));
    InMux I__10434 (
            .O(N__51279),
            .I(N__51276));
    LocalMux I__10433 (
            .O(N__51276),
            .I(N__51272));
    InMux I__10432 (
            .O(N__51275),
            .I(N__51269));
    Odrv4 I__10431 (
            .O(N__51272),
            .I(\c0.n109 ));
    LocalMux I__10430 (
            .O(N__51269),
            .I(\c0.n109 ));
    CascadeMux I__10429 (
            .O(N__51264),
            .I(N__51261));
    InMux I__10428 (
            .O(N__51261),
            .I(N__51258));
    LocalMux I__10427 (
            .O(N__51258),
            .I(N__51255));
    Odrv4 I__10426 (
            .O(N__51255),
            .I(\c0.n23_adj_4590 ));
    InMux I__10425 (
            .O(N__51252),
            .I(N__51249));
    LocalMux I__10424 (
            .O(N__51249),
            .I(N__51246));
    Span4Mux_h I__10423 (
            .O(N__51246),
            .I(N__51243));
    Odrv4 I__10422 (
            .O(N__51243),
            .I(\c0.n29_adj_4734 ));
    CascadeMux I__10421 (
            .O(N__51240),
            .I(\c0.n20_adj_4290_cascade_ ));
    InMux I__10420 (
            .O(N__51237),
            .I(N__51234));
    LocalMux I__10419 (
            .O(N__51234),
            .I(N__51229));
    InMux I__10418 (
            .O(N__51233),
            .I(N__51224));
    InMux I__10417 (
            .O(N__51232),
            .I(N__51224));
    Span4Mux_v I__10416 (
            .O(N__51229),
            .I(N__51220));
    LocalMux I__10415 (
            .O(N__51224),
            .I(N__51213));
    InMux I__10414 (
            .O(N__51223),
            .I(N__51208));
    Sp12to4 I__10413 (
            .O(N__51220),
            .I(N__51203));
    InMux I__10412 (
            .O(N__51219),
            .I(N__51200));
    InMux I__10411 (
            .O(N__51218),
            .I(N__51197));
    InMux I__10410 (
            .O(N__51217),
            .I(N__51192));
    InMux I__10409 (
            .O(N__51216),
            .I(N__51192));
    Span4Mux_v I__10408 (
            .O(N__51213),
            .I(N__51189));
    InMux I__10407 (
            .O(N__51212),
            .I(N__51184));
    InMux I__10406 (
            .O(N__51211),
            .I(N__51184));
    LocalMux I__10405 (
            .O(N__51208),
            .I(N__51181));
    InMux I__10404 (
            .O(N__51207),
            .I(N__51176));
    InMux I__10403 (
            .O(N__51206),
            .I(N__51176));
    Odrv12 I__10402 (
            .O(N__51203),
            .I(data_in_frame_1_1));
    LocalMux I__10401 (
            .O(N__51200),
            .I(data_in_frame_1_1));
    LocalMux I__10400 (
            .O(N__51197),
            .I(data_in_frame_1_1));
    LocalMux I__10399 (
            .O(N__51192),
            .I(data_in_frame_1_1));
    Odrv4 I__10398 (
            .O(N__51189),
            .I(data_in_frame_1_1));
    LocalMux I__10397 (
            .O(N__51184),
            .I(data_in_frame_1_1));
    Odrv4 I__10396 (
            .O(N__51181),
            .I(data_in_frame_1_1));
    LocalMux I__10395 (
            .O(N__51176),
            .I(data_in_frame_1_1));
    InMux I__10394 (
            .O(N__51159),
            .I(N__51156));
    LocalMux I__10393 (
            .O(N__51156),
            .I(N__51153));
    Odrv12 I__10392 (
            .O(N__51153),
            .I(\c0.n51 ));
    InMux I__10391 (
            .O(N__51150),
            .I(N__51144));
    InMux I__10390 (
            .O(N__51149),
            .I(N__51144));
    LocalMux I__10389 (
            .O(N__51144),
            .I(\c0.n29 ));
    CascadeMux I__10388 (
            .O(N__51141),
            .I(\c0.n51_cascade_ ));
    InMux I__10387 (
            .O(N__51138),
            .I(N__51131));
    InMux I__10386 (
            .O(N__51137),
            .I(N__51131));
    InMux I__10385 (
            .O(N__51136),
            .I(N__51128));
    LocalMux I__10384 (
            .O(N__51131),
            .I(N__51125));
    LocalMux I__10383 (
            .O(N__51128),
            .I(\c0.n22_adj_4647 ));
    Odrv4 I__10382 (
            .O(N__51125),
            .I(\c0.n22_adj_4647 ));
    CascadeMux I__10381 (
            .O(N__51120),
            .I(\c0.n102_cascade_ ));
    InMux I__10380 (
            .O(N__51117),
            .I(N__51114));
    LocalMux I__10379 (
            .O(N__51114),
            .I(\c0.n32 ));
    CascadeMux I__10378 (
            .O(N__51111),
            .I(\c0.n16_adj_4256_cascade_ ));
    CascadeMux I__10377 (
            .O(N__51108),
            .I(N__51105));
    InMux I__10376 (
            .O(N__51105),
            .I(N__51102));
    LocalMux I__10375 (
            .O(N__51102),
            .I(\c0.n9_adj_4279 ));
    CascadeMux I__10374 (
            .O(N__51099),
            .I(N__51096));
    InMux I__10373 (
            .O(N__51096),
            .I(N__51093));
    LocalMux I__10372 (
            .O(N__51093),
            .I(N__51089));
    InMux I__10371 (
            .O(N__51092),
            .I(N__51086));
    Span4Mux_h I__10370 (
            .O(N__51089),
            .I(N__51082));
    LocalMux I__10369 (
            .O(N__51086),
            .I(N__51079));
    InMux I__10368 (
            .O(N__51085),
            .I(N__51076));
    Odrv4 I__10367 (
            .O(N__51082),
            .I(\c0.n13141 ));
    Odrv12 I__10366 (
            .O(N__51079),
            .I(\c0.n13141 ));
    LocalMux I__10365 (
            .O(N__51076),
            .I(\c0.n13141 ));
    CascadeMux I__10364 (
            .O(N__51069),
            .I(\c0.n9_adj_4279_cascade_ ));
    CascadeMux I__10363 (
            .O(N__51066),
            .I(\c0.n23574_cascade_ ));
    InMux I__10362 (
            .O(N__51063),
            .I(N__51060));
    LocalMux I__10361 (
            .O(N__51060),
            .I(\c0.n11_adj_4257 ));
    CascadeMux I__10360 (
            .O(N__51057),
            .I(\c0.n38_adj_4285_cascade_ ));
    InMux I__10359 (
            .O(N__51054),
            .I(N__51051));
    LocalMux I__10358 (
            .O(N__51051),
            .I(\c0.n26_adj_4289 ));
    CascadeMux I__10357 (
            .O(N__51048),
            .I(\c0.n26_adj_4289_cascade_ ));
    InMux I__10356 (
            .O(N__51045),
            .I(N__51041));
    InMux I__10355 (
            .O(N__51044),
            .I(N__51038));
    LocalMux I__10354 (
            .O(N__51041),
            .I(N__51035));
    LocalMux I__10353 (
            .O(N__51038),
            .I(\c0.data_out_frame_0__7__N_2626 ));
    Odrv4 I__10352 (
            .O(N__51035),
            .I(\c0.data_out_frame_0__7__N_2626 ));
    InMux I__10351 (
            .O(N__51030),
            .I(N__51024));
    InMux I__10350 (
            .O(N__51029),
            .I(N__51024));
    LocalMux I__10349 (
            .O(N__51024),
            .I(\c0.n20_adj_4290 ));
    InMux I__10348 (
            .O(N__51021),
            .I(N__51018));
    LocalMux I__10347 (
            .O(N__51018),
            .I(\c0.n12_adj_4657 ));
    CascadeMux I__10346 (
            .O(N__51015),
            .I(N__51012));
    InMux I__10345 (
            .O(N__51012),
            .I(N__51009));
    LocalMux I__10344 (
            .O(N__51009),
            .I(N__51006));
    Span4Mux_h I__10343 (
            .O(N__51006),
            .I(N__51003));
    Odrv4 I__10342 (
            .O(N__51003),
            .I(\c0.n23_adj_4648 ));
    InMux I__10341 (
            .O(N__51000),
            .I(N__50997));
    LocalMux I__10340 (
            .O(N__50997),
            .I(\c0.n39_adj_4737 ));
    InMux I__10339 (
            .O(N__50994),
            .I(N__50991));
    LocalMux I__10338 (
            .O(N__50991),
            .I(\c0.n38_adj_4736 ));
    CascadeMux I__10337 (
            .O(N__50988),
            .I(N__50985));
    InMux I__10336 (
            .O(N__50985),
            .I(N__50979));
    InMux I__10335 (
            .O(N__50984),
            .I(N__50979));
    LocalMux I__10334 (
            .O(N__50979),
            .I(\c0.n23562 ));
    CascadeMux I__10333 (
            .O(N__50976),
            .I(\c0.n23562_cascade_ ));
    InMux I__10332 (
            .O(N__50973),
            .I(N__50966));
    InMux I__10331 (
            .O(N__50972),
            .I(N__50961));
    InMux I__10330 (
            .O(N__50971),
            .I(N__50961));
    InMux I__10329 (
            .O(N__50970),
            .I(N__50956));
    InMux I__10328 (
            .O(N__50969),
            .I(N__50956));
    LocalMux I__10327 (
            .O(N__50966),
            .I(data_in_frame_5_5));
    LocalMux I__10326 (
            .O(N__50961),
            .I(data_in_frame_5_5));
    LocalMux I__10325 (
            .O(N__50956),
            .I(data_in_frame_5_5));
    CascadeMux I__10324 (
            .O(N__50949),
            .I(N__50946));
    InMux I__10323 (
            .O(N__50946),
            .I(N__50937));
    InMux I__10322 (
            .O(N__50945),
            .I(N__50932));
    InMux I__10321 (
            .O(N__50944),
            .I(N__50932));
    InMux I__10320 (
            .O(N__50943),
            .I(N__50927));
    InMux I__10319 (
            .O(N__50942),
            .I(N__50927));
    InMux I__10318 (
            .O(N__50941),
            .I(N__50922));
    InMux I__10317 (
            .O(N__50940),
            .I(N__50922));
    LocalMux I__10316 (
            .O(N__50937),
            .I(\c0.data_in_frame_3_4 ));
    LocalMux I__10315 (
            .O(N__50932),
            .I(\c0.data_in_frame_3_4 ));
    LocalMux I__10314 (
            .O(N__50927),
            .I(\c0.data_in_frame_3_4 ));
    LocalMux I__10313 (
            .O(N__50922),
            .I(\c0.data_in_frame_3_4 ));
    CascadeMux I__10312 (
            .O(N__50913),
            .I(N__50905));
    CascadeMux I__10311 (
            .O(N__50912),
            .I(N__50901));
    CascadeMux I__10310 (
            .O(N__50911),
            .I(N__50898));
    CascadeMux I__10309 (
            .O(N__50910),
            .I(N__50895));
    InMux I__10308 (
            .O(N__50909),
            .I(N__50892));
    CascadeMux I__10307 (
            .O(N__50908),
            .I(N__50889));
    InMux I__10306 (
            .O(N__50905),
            .I(N__50886));
    CascadeMux I__10305 (
            .O(N__50904),
            .I(N__50883));
    InMux I__10304 (
            .O(N__50901),
            .I(N__50880));
    InMux I__10303 (
            .O(N__50898),
            .I(N__50877));
    InMux I__10302 (
            .O(N__50895),
            .I(N__50874));
    LocalMux I__10301 (
            .O(N__50892),
            .I(N__50871));
    InMux I__10300 (
            .O(N__50889),
            .I(N__50868));
    LocalMux I__10299 (
            .O(N__50886),
            .I(N__50861));
    InMux I__10298 (
            .O(N__50883),
            .I(N__50858));
    LocalMux I__10297 (
            .O(N__50880),
            .I(N__50851));
    LocalMux I__10296 (
            .O(N__50877),
            .I(N__50851));
    LocalMux I__10295 (
            .O(N__50874),
            .I(N__50851));
    Span4Mux_s3_v I__10294 (
            .O(N__50871),
            .I(N__50848));
    LocalMux I__10293 (
            .O(N__50868),
            .I(N__50845));
    InMux I__10292 (
            .O(N__50867),
            .I(N__50842));
    InMux I__10291 (
            .O(N__50866),
            .I(N__50837));
    InMux I__10290 (
            .O(N__50865),
            .I(N__50837));
    CascadeMux I__10289 (
            .O(N__50864),
            .I(N__50834));
    Span4Mux_v I__10288 (
            .O(N__50861),
            .I(N__50829));
    LocalMux I__10287 (
            .O(N__50858),
            .I(N__50829));
    Span4Mux_h I__10286 (
            .O(N__50851),
            .I(N__50826));
    Span4Mux_h I__10285 (
            .O(N__50848),
            .I(N__50822));
    Span4Mux_v I__10284 (
            .O(N__50845),
            .I(N__50817));
    LocalMux I__10283 (
            .O(N__50842),
            .I(N__50817));
    LocalMux I__10282 (
            .O(N__50837),
            .I(N__50814));
    InMux I__10281 (
            .O(N__50834),
            .I(N__50811));
    Span4Mux_v I__10280 (
            .O(N__50829),
            .I(N__50808));
    Span4Mux_h I__10279 (
            .O(N__50826),
            .I(N__50805));
    InMux I__10278 (
            .O(N__50825),
            .I(N__50802));
    Sp12to4 I__10277 (
            .O(N__50822),
            .I(N__50799));
    Span4Mux_h I__10276 (
            .O(N__50817),
            .I(N__50796));
    Span4Mux_v I__10275 (
            .O(N__50814),
            .I(N__50793));
    LocalMux I__10274 (
            .O(N__50811),
            .I(N__50790));
    Span4Mux_h I__10273 (
            .O(N__50808),
            .I(N__50787));
    Span4Mux_h I__10272 (
            .O(N__50805),
            .I(N__50782));
    LocalMux I__10271 (
            .O(N__50802),
            .I(N__50782));
    Span12Mux_h I__10270 (
            .O(N__50799),
            .I(N__50779));
    Span4Mux_h I__10269 (
            .O(N__50796),
            .I(N__50776));
    Span4Mux_h I__10268 (
            .O(N__50793),
            .I(N__50773));
    Sp12to4 I__10267 (
            .O(N__50790),
            .I(N__50770));
    Span4Mux_h I__10266 (
            .O(N__50787),
            .I(N__50767));
    Sp12to4 I__10265 (
            .O(N__50782),
            .I(N__50760));
    Span12Mux_v I__10264 (
            .O(N__50779),
            .I(N__50760));
    Sp12to4 I__10263 (
            .O(N__50776),
            .I(N__50760));
    Span4Mux_h I__10262 (
            .O(N__50773),
            .I(N__50757));
    Span12Mux_h I__10261 (
            .O(N__50770),
            .I(N__50754));
    Span4Mux_h I__10260 (
            .O(N__50767),
            .I(N__50751));
    Span12Mux_v I__10259 (
            .O(N__50760),
            .I(N__50748));
    Span4Mux_v I__10258 (
            .O(N__50757),
            .I(N__50745));
    Odrv12 I__10257 (
            .O(N__50754),
            .I(r_Rx_Data));
    Odrv4 I__10256 (
            .O(N__50751),
            .I(r_Rx_Data));
    Odrv12 I__10255 (
            .O(N__50748),
            .I(r_Rx_Data));
    Odrv4 I__10254 (
            .O(N__50745),
            .I(r_Rx_Data));
    CascadeMux I__10253 (
            .O(N__50736),
            .I(n4_cascade_));
    InMux I__10252 (
            .O(N__50733),
            .I(N__50730));
    LocalMux I__10251 (
            .O(N__50730),
            .I(N__50727));
    Span4Mux_s2_v I__10250 (
            .O(N__50727),
            .I(N__50723));
    InMux I__10249 (
            .O(N__50726),
            .I(N__50720));
    Sp12to4 I__10248 (
            .O(N__50723),
            .I(N__50715));
    LocalMux I__10247 (
            .O(N__50720),
            .I(N__50712));
    InMux I__10246 (
            .O(N__50719),
            .I(N__50709));
    InMux I__10245 (
            .O(N__50718),
            .I(N__50706));
    Span12Mux_h I__10244 (
            .O(N__50715),
            .I(N__50703));
    Span4Mux_h I__10243 (
            .O(N__50712),
            .I(N__50698));
    LocalMux I__10242 (
            .O(N__50709),
            .I(N__50698));
    LocalMux I__10241 (
            .O(N__50706),
            .I(N__50695));
    Span12Mux_v I__10240 (
            .O(N__50703),
            .I(N__50692));
    Span4Mux_v I__10239 (
            .O(N__50698),
            .I(N__50689));
    Span4Mux_v I__10238 (
            .O(N__50695),
            .I(N__50686));
    Odrv12 I__10237 (
            .O(N__50692),
            .I(n12904));
    Odrv4 I__10236 (
            .O(N__50689),
            .I(n12904));
    Odrv4 I__10235 (
            .O(N__50686),
            .I(n12904));
    InMux I__10234 (
            .O(N__50679),
            .I(N__50676));
    LocalMux I__10233 (
            .O(N__50676),
            .I(N__50673));
    Span12Mux_s4_v I__10232 (
            .O(N__50673),
            .I(N__50670));
    Span12Mux_v I__10231 (
            .O(N__50670),
            .I(N__50667));
    Odrv12 I__10230 (
            .O(N__50667),
            .I(\c0.rx.n14277 ));
    InMux I__10229 (
            .O(N__50664),
            .I(N__50661));
    LocalMux I__10228 (
            .O(N__50661),
            .I(N__50658));
    Sp12to4 I__10227 (
            .O(N__50658),
            .I(N__50655));
    Span12Mux_s3_v I__10226 (
            .O(N__50655),
            .I(N__50652));
    Span12Mux_v I__10225 (
            .O(N__50652),
            .I(N__50647));
    InMux I__10224 (
            .O(N__50651),
            .I(N__50644));
    InMux I__10223 (
            .O(N__50650),
            .I(N__50641));
    Odrv12 I__10222 (
            .O(N__50647),
            .I(\c0.n12514 ));
    LocalMux I__10221 (
            .O(N__50644),
            .I(\c0.n12514 ));
    LocalMux I__10220 (
            .O(N__50641),
            .I(\c0.n12514 ));
    InMux I__10219 (
            .O(N__50634),
            .I(N__50631));
    LocalMux I__10218 (
            .O(N__50631),
            .I(N__50628));
    Span4Mux_h I__10217 (
            .O(N__50628),
            .I(N__50625));
    Span4Mux_v I__10216 (
            .O(N__50625),
            .I(N__50622));
    Span4Mux_v I__10215 (
            .O(N__50622),
            .I(N__50617));
    InMux I__10214 (
            .O(N__50621),
            .I(N__50614));
    InMux I__10213 (
            .O(N__50620),
            .I(N__50611));
    Span4Mux_v I__10212 (
            .O(N__50617),
            .I(N__50606));
    LocalMux I__10211 (
            .O(N__50614),
            .I(N__50606));
    LocalMux I__10210 (
            .O(N__50611),
            .I(N__50601));
    Span4Mux_h I__10209 (
            .O(N__50606),
            .I(N__50601));
    Odrv4 I__10208 (
            .O(N__50601),
            .I(\c0.n20641 ));
    CascadeMux I__10207 (
            .O(N__50598),
            .I(N__50595));
    InMux I__10206 (
            .O(N__50595),
            .I(N__50592));
    LocalMux I__10205 (
            .O(N__50592),
            .I(N__50589));
    Span4Mux_s3_v I__10204 (
            .O(N__50589),
            .I(N__50585));
    InMux I__10203 (
            .O(N__50588),
            .I(N__50581));
    Span4Mux_h I__10202 (
            .O(N__50585),
            .I(N__50578));
    InMux I__10201 (
            .O(N__50584),
            .I(N__50575));
    LocalMux I__10200 (
            .O(N__50581),
            .I(N__50571));
    Span4Mux_h I__10199 (
            .O(N__50578),
            .I(N__50568));
    LocalMux I__10198 (
            .O(N__50575),
            .I(N__50565));
    InMux I__10197 (
            .O(N__50574),
            .I(N__50562));
    Span4Mux_h I__10196 (
            .O(N__50571),
            .I(N__50559));
    Sp12to4 I__10195 (
            .O(N__50568),
            .I(N__50556));
    Span4Mux_h I__10194 (
            .O(N__50565),
            .I(N__50553));
    LocalMux I__10193 (
            .O(N__50562),
            .I(N__50550));
    Odrv4 I__10192 (
            .O(N__50559),
            .I(\c0.n21391 ));
    Odrv12 I__10191 (
            .O(N__50556),
            .I(\c0.n21391 ));
    Odrv4 I__10190 (
            .O(N__50553),
            .I(\c0.n21391 ));
    Odrv4 I__10189 (
            .O(N__50550),
            .I(\c0.n21391 ));
    InMux I__10188 (
            .O(N__50541),
            .I(N__50538));
    LocalMux I__10187 (
            .O(N__50538),
            .I(N__50535));
    Span4Mux_h I__10186 (
            .O(N__50535),
            .I(N__50532));
    Sp12to4 I__10185 (
            .O(N__50532),
            .I(N__50529));
    Span12Mux_v I__10184 (
            .O(N__50529),
            .I(N__50523));
    InMux I__10183 (
            .O(N__50528),
            .I(N__50520));
    InMux I__10182 (
            .O(N__50527),
            .I(N__50517));
    InMux I__10181 (
            .O(N__50526),
            .I(N__50514));
    Odrv12 I__10180 (
            .O(N__50523),
            .I(\c0.n21360 ));
    LocalMux I__10179 (
            .O(N__50520),
            .I(\c0.n21360 ));
    LocalMux I__10178 (
            .O(N__50517),
            .I(\c0.n21360 ));
    LocalMux I__10177 (
            .O(N__50514),
            .I(\c0.n21360 ));
    InMux I__10176 (
            .O(N__50505),
            .I(N__50502));
    LocalMux I__10175 (
            .O(N__50502),
            .I(N__50499));
    Span4Mux_h I__10174 (
            .O(N__50499),
            .I(N__50496));
    Span4Mux_h I__10173 (
            .O(N__50496),
            .I(N__50493));
    Sp12to4 I__10172 (
            .O(N__50493),
            .I(N__50490));
    Span12Mux_v I__10171 (
            .O(N__50490),
            .I(N__50487));
    Odrv12 I__10170 (
            .O(N__50487),
            .I(\c0.n21_adj_4719 ));
    InMux I__10169 (
            .O(N__50484),
            .I(N__50477));
    InMux I__10168 (
            .O(N__50483),
            .I(N__50474));
    InMux I__10167 (
            .O(N__50482),
            .I(N__50467));
    InMux I__10166 (
            .O(N__50481),
            .I(N__50467));
    InMux I__10165 (
            .O(N__50480),
            .I(N__50455));
    LocalMux I__10164 (
            .O(N__50477),
            .I(N__50448));
    LocalMux I__10163 (
            .O(N__50474),
            .I(N__50448));
    InMux I__10162 (
            .O(N__50473),
            .I(N__50445));
    InMux I__10161 (
            .O(N__50472),
            .I(N__50442));
    LocalMux I__10160 (
            .O(N__50467),
            .I(N__50439));
    InMux I__10159 (
            .O(N__50466),
            .I(N__50433));
    CascadeMux I__10158 (
            .O(N__50465),
            .I(N__50430));
    InMux I__10157 (
            .O(N__50464),
            .I(N__50420));
    InMux I__10156 (
            .O(N__50463),
            .I(N__50417));
    InMux I__10155 (
            .O(N__50462),
            .I(N__50410));
    InMux I__10154 (
            .O(N__50461),
            .I(N__50410));
    InMux I__10153 (
            .O(N__50460),
            .I(N__50410));
    InMux I__10152 (
            .O(N__50459),
            .I(N__50405));
    InMux I__10151 (
            .O(N__50458),
            .I(N__50405));
    LocalMux I__10150 (
            .O(N__50455),
            .I(N__50398));
    InMux I__10149 (
            .O(N__50454),
            .I(N__50395));
    InMux I__10148 (
            .O(N__50453),
            .I(N__50392));
    Span4Mux_h I__10147 (
            .O(N__50448),
            .I(N__50386));
    LocalMux I__10146 (
            .O(N__50445),
            .I(N__50386));
    LocalMux I__10145 (
            .O(N__50442),
            .I(N__50381));
    Span4Mux_v I__10144 (
            .O(N__50439),
            .I(N__50381));
    InMux I__10143 (
            .O(N__50438),
            .I(N__50378));
    InMux I__10142 (
            .O(N__50437),
            .I(N__50375));
    InMux I__10141 (
            .O(N__50436),
            .I(N__50372));
    LocalMux I__10140 (
            .O(N__50433),
            .I(N__50369));
    InMux I__10139 (
            .O(N__50430),
            .I(N__50362));
    InMux I__10138 (
            .O(N__50429),
            .I(N__50362));
    InMux I__10137 (
            .O(N__50428),
            .I(N__50362));
    InMux I__10136 (
            .O(N__50427),
            .I(N__50359));
    InMux I__10135 (
            .O(N__50426),
            .I(N__50356));
    InMux I__10134 (
            .O(N__50425),
            .I(N__50353));
    InMux I__10133 (
            .O(N__50424),
            .I(N__50348));
    InMux I__10132 (
            .O(N__50423),
            .I(N__50348));
    LocalMux I__10131 (
            .O(N__50420),
            .I(N__50339));
    LocalMux I__10130 (
            .O(N__50417),
            .I(N__50339));
    LocalMux I__10129 (
            .O(N__50410),
            .I(N__50339));
    LocalMux I__10128 (
            .O(N__50405),
            .I(N__50339));
    InMux I__10127 (
            .O(N__50404),
            .I(N__50334));
    InMux I__10126 (
            .O(N__50403),
            .I(N__50334));
    InMux I__10125 (
            .O(N__50402),
            .I(N__50329));
    InMux I__10124 (
            .O(N__50401),
            .I(N__50329));
    Span4Mux_v I__10123 (
            .O(N__50398),
            .I(N__50326));
    LocalMux I__10122 (
            .O(N__50395),
            .I(N__50323));
    LocalMux I__10121 (
            .O(N__50392),
            .I(N__50320));
    InMux I__10120 (
            .O(N__50391),
            .I(N__50317));
    Span4Mux_v I__10119 (
            .O(N__50386),
            .I(N__50314));
    Span4Mux_v I__10118 (
            .O(N__50381),
            .I(N__50311));
    LocalMux I__10117 (
            .O(N__50378),
            .I(N__50306));
    LocalMux I__10116 (
            .O(N__50375),
            .I(N__50306));
    LocalMux I__10115 (
            .O(N__50372),
            .I(N__50301));
    Span4Mux_v I__10114 (
            .O(N__50369),
            .I(N__50301));
    LocalMux I__10113 (
            .O(N__50362),
            .I(N__50286));
    LocalMux I__10112 (
            .O(N__50359),
            .I(N__50286));
    LocalMux I__10111 (
            .O(N__50356),
            .I(N__50286));
    LocalMux I__10110 (
            .O(N__50353),
            .I(N__50286));
    LocalMux I__10109 (
            .O(N__50348),
            .I(N__50286));
    Span4Mux_v I__10108 (
            .O(N__50339),
            .I(N__50286));
    LocalMux I__10107 (
            .O(N__50334),
            .I(N__50286));
    LocalMux I__10106 (
            .O(N__50329),
            .I(N__50283));
    Span4Mux_h I__10105 (
            .O(N__50326),
            .I(N__50278));
    Span4Mux_v I__10104 (
            .O(N__50323),
            .I(N__50278));
    Span4Mux_v I__10103 (
            .O(N__50320),
            .I(N__50273));
    LocalMux I__10102 (
            .O(N__50317),
            .I(N__50273));
    Span4Mux_v I__10101 (
            .O(N__50314),
            .I(N__50268));
    Span4Mux_v I__10100 (
            .O(N__50311),
            .I(N__50268));
    Span4Mux_v I__10099 (
            .O(N__50306),
            .I(N__50261));
    Span4Mux_v I__10098 (
            .O(N__50301),
            .I(N__50261));
    Span4Mux_v I__10097 (
            .O(N__50286),
            .I(N__50261));
    Span4Mux_h I__10096 (
            .O(N__50283),
            .I(N__50256));
    Span4Mux_v I__10095 (
            .O(N__50278),
            .I(N__50256));
    Sp12to4 I__10094 (
            .O(N__50273),
            .I(N__50253));
    Span4Mux_h I__10093 (
            .O(N__50268),
            .I(N__50250));
    Sp12to4 I__10092 (
            .O(N__50261),
            .I(N__50247));
    Span4Mux_v I__10091 (
            .O(N__50256),
            .I(N__50244));
    Span12Mux_v I__10090 (
            .O(N__50253),
            .I(N__50241));
    Sp12to4 I__10089 (
            .O(N__50250),
            .I(N__50236));
    Span12Mux_h I__10088 (
            .O(N__50247),
            .I(N__50236));
    Span4Mux_v I__10087 (
            .O(N__50244),
            .I(N__50230));
    Span12Mux_v I__10086 (
            .O(N__50241),
            .I(N__50227));
    Span12Mux_v I__10085 (
            .O(N__50236),
            .I(N__50224));
    InMux I__10084 (
            .O(N__50235),
            .I(N__50217));
    InMux I__10083 (
            .O(N__50234),
            .I(N__50217));
    InMux I__10082 (
            .O(N__50233),
            .I(N__50217));
    Odrv4 I__10081 (
            .O(N__50230),
            .I(rx_data_ready));
    Odrv12 I__10080 (
            .O(N__50227),
            .I(rx_data_ready));
    Odrv12 I__10079 (
            .O(N__50224),
            .I(rx_data_ready));
    LocalMux I__10078 (
            .O(N__50217),
            .I(rx_data_ready));
    InMux I__10077 (
            .O(N__50208),
            .I(N__50205));
    LocalMux I__10076 (
            .O(N__50205),
            .I(N__50202));
    Sp12to4 I__10075 (
            .O(N__50202),
            .I(N__50199));
    Span12Mux_h I__10074 (
            .O(N__50199),
            .I(N__50195));
    InMux I__10073 (
            .O(N__50198),
            .I(N__50192));
    Span12Mux_v I__10072 (
            .O(N__50195),
            .I(N__50189));
    LocalMux I__10071 (
            .O(N__50192),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    Odrv12 I__10070 (
            .O(N__50189),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    CascadeMux I__10069 (
            .O(N__50184),
            .I(N__50180));
    CascadeMux I__10068 (
            .O(N__50183),
            .I(N__50174));
    InMux I__10067 (
            .O(N__50180),
            .I(N__50169));
    InMux I__10066 (
            .O(N__50179),
            .I(N__50169));
    CascadeMux I__10065 (
            .O(N__50178),
            .I(N__50166));
    CascadeMux I__10064 (
            .O(N__50177),
            .I(N__50163));
    InMux I__10063 (
            .O(N__50174),
            .I(N__50158));
    LocalMux I__10062 (
            .O(N__50169),
            .I(N__50154));
    InMux I__10061 (
            .O(N__50166),
            .I(N__50150));
    InMux I__10060 (
            .O(N__50163),
            .I(N__50147));
    CascadeMux I__10059 (
            .O(N__50162),
            .I(N__50144));
    InMux I__10058 (
            .O(N__50161),
            .I(N__50141));
    LocalMux I__10057 (
            .O(N__50158),
            .I(N__50138));
    CascadeMux I__10056 (
            .O(N__50157),
            .I(N__50135));
    Span12Mux_h I__10055 (
            .O(N__50154),
            .I(N__50132));
    InMux I__10054 (
            .O(N__50153),
            .I(N__50129));
    LocalMux I__10053 (
            .O(N__50150),
            .I(N__50126));
    LocalMux I__10052 (
            .O(N__50147),
            .I(N__50123));
    InMux I__10051 (
            .O(N__50144),
            .I(N__50120));
    LocalMux I__10050 (
            .O(N__50141),
            .I(N__50117));
    Span4Mux_v I__10049 (
            .O(N__50138),
            .I(N__50114));
    InMux I__10048 (
            .O(N__50135),
            .I(N__50111));
    Span12Mux_v I__10047 (
            .O(N__50132),
            .I(N__50108));
    LocalMux I__10046 (
            .O(N__50129),
            .I(N__50103));
    Span4Mux_h I__10045 (
            .O(N__50126),
            .I(N__50100));
    Span4Mux_h I__10044 (
            .O(N__50123),
            .I(N__50095));
    LocalMux I__10043 (
            .O(N__50120),
            .I(N__50095));
    Span4Mux_v I__10042 (
            .O(N__50117),
            .I(N__50090));
    Span4Mux_v I__10041 (
            .O(N__50114),
            .I(N__50090));
    LocalMux I__10040 (
            .O(N__50111),
            .I(N__50087));
    Span12Mux_v I__10039 (
            .O(N__50108),
            .I(N__50084));
    InMux I__10038 (
            .O(N__50107),
            .I(N__50079));
    InMux I__10037 (
            .O(N__50106),
            .I(N__50079));
    Span12Mux_h I__10036 (
            .O(N__50103),
            .I(N__50076));
    Span4Mux_v I__10035 (
            .O(N__50100),
            .I(N__50071));
    Span4Mux_h I__10034 (
            .O(N__50095),
            .I(N__50071));
    Span4Mux_h I__10033 (
            .O(N__50090),
            .I(N__50066));
    Span4Mux_v I__10032 (
            .O(N__50087),
            .I(N__50066));
    Odrv12 I__10031 (
            .O(N__50084),
            .I(r_SM_Main_1));
    LocalMux I__10030 (
            .O(N__50079),
            .I(r_SM_Main_1));
    Odrv12 I__10029 (
            .O(N__50076),
            .I(r_SM_Main_1));
    Odrv4 I__10028 (
            .O(N__50071),
            .I(r_SM_Main_1));
    Odrv4 I__10027 (
            .O(N__50066),
            .I(r_SM_Main_1));
    InMux I__10026 (
            .O(N__50055),
            .I(N__50052));
    LocalMux I__10025 (
            .O(N__50052),
            .I(N__50049));
    Span4Mux_s0_v I__10024 (
            .O(N__50049),
            .I(N__50045));
    InMux I__10023 (
            .O(N__50048),
            .I(N__50039));
    Sp12to4 I__10022 (
            .O(N__50045),
            .I(N__50036));
    InMux I__10021 (
            .O(N__50044),
            .I(N__50031));
    InMux I__10020 (
            .O(N__50043),
            .I(N__50026));
    InMux I__10019 (
            .O(N__50042),
            .I(N__50026));
    LocalMux I__10018 (
            .O(N__50039),
            .I(N__50022));
    Span12Mux_s4_v I__10017 (
            .O(N__50036),
            .I(N__50019));
    InMux I__10016 (
            .O(N__50035),
            .I(N__50016));
    InMux I__10015 (
            .O(N__50034),
            .I(N__50013));
    LocalMux I__10014 (
            .O(N__50031),
            .I(N__50010));
    LocalMux I__10013 (
            .O(N__50026),
            .I(N__50007));
    InMux I__10012 (
            .O(N__50025),
            .I(N__50004));
    Span4Mux_v I__10011 (
            .O(N__50022),
            .I(N__50001));
    Span12Mux_h I__10010 (
            .O(N__50019),
            .I(N__49997));
    LocalMux I__10009 (
            .O(N__50016),
            .I(N__49992));
    LocalMux I__10008 (
            .O(N__50013),
            .I(N__49992));
    Span4Mux_h I__10007 (
            .O(N__50010),
            .I(N__49985));
    Span4Mux_v I__10006 (
            .O(N__50007),
            .I(N__49985));
    LocalMux I__10005 (
            .O(N__50004),
            .I(N__49985));
    Span4Mux_h I__10004 (
            .O(N__50001),
            .I(N__49982));
    InMux I__10003 (
            .O(N__50000),
            .I(N__49979));
    Span12Mux_v I__10002 (
            .O(N__49997),
            .I(N__49974));
    Span12Mux_h I__10001 (
            .O(N__49992),
            .I(N__49974));
    Span4Mux_h I__10000 (
            .O(N__49985),
            .I(N__49971));
    Odrv4 I__9999 (
            .O(N__49982),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__9998 (
            .O(N__49979),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv12 I__9997 (
            .O(N__49974),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__9996 (
            .O(N__49971),
            .I(\c0.rx.r_SM_Main_0 ));
    InMux I__9995 (
            .O(N__49962),
            .I(N__49959));
    LocalMux I__9994 (
            .O(N__49959),
            .I(N__49953));
    InMux I__9993 (
            .O(N__49958),
            .I(N__49948));
    InMux I__9992 (
            .O(N__49957),
            .I(N__49948));
    InMux I__9991 (
            .O(N__49956),
            .I(N__49945));
    Span4Mux_h I__9990 (
            .O(N__49953),
            .I(N__49935));
    LocalMux I__9989 (
            .O(N__49948),
            .I(N__49935));
    LocalMux I__9988 (
            .O(N__49945),
            .I(N__49932));
    InMux I__9987 (
            .O(N__49944),
            .I(N__49929));
    InMux I__9986 (
            .O(N__49943),
            .I(N__49924));
    InMux I__9985 (
            .O(N__49942),
            .I(N__49924));
    InMux I__9984 (
            .O(N__49941),
            .I(N__49921));
    InMux I__9983 (
            .O(N__49940),
            .I(N__49918));
    Span4Mux_h I__9982 (
            .O(N__49935),
            .I(N__49915));
    Span4Mux_h I__9981 (
            .O(N__49932),
            .I(N__49910));
    LocalMux I__9980 (
            .O(N__49929),
            .I(N__49910));
    LocalMux I__9979 (
            .O(N__49924),
            .I(N__49907));
    LocalMux I__9978 (
            .O(N__49921),
            .I(N__49904));
    LocalMux I__9977 (
            .O(N__49918),
            .I(N__49901));
    Sp12to4 I__9976 (
            .O(N__49915),
            .I(N__49896));
    Sp12to4 I__9975 (
            .O(N__49910),
            .I(N__49896));
    Span12Mux_s8_v I__9974 (
            .O(N__49907),
            .I(N__49893));
    Span12Mux_s9_h I__9973 (
            .O(N__49904),
            .I(N__49886));
    Span12Mux_h I__9972 (
            .O(N__49901),
            .I(N__49886));
    Span12Mux_v I__9971 (
            .O(N__49896),
            .I(N__49886));
    Odrv12 I__9970 (
            .O(N__49893),
            .I(r_SM_Main_2));
    Odrv12 I__9969 (
            .O(N__49886),
            .I(r_SM_Main_2));
    SRMux I__9968 (
            .O(N__49881),
            .I(N__49878));
    LocalMux I__9967 (
            .O(N__49878),
            .I(N__49875));
    Span4Mux_h I__9966 (
            .O(N__49875),
            .I(N__49872));
    Sp12to4 I__9965 (
            .O(N__49872),
            .I(N__49869));
    Span12Mux_v I__9964 (
            .O(N__49869),
            .I(N__49866));
    Odrv12 I__9963 (
            .O(N__49866),
            .I(\c0.rx.n22094 ));
    InMux I__9962 (
            .O(N__49863),
            .I(N__49860));
    LocalMux I__9961 (
            .O(N__49860),
            .I(\c0.n46_adj_4739 ));
    InMux I__9960 (
            .O(N__49857),
            .I(N__49854));
    LocalMux I__9959 (
            .O(N__49854),
            .I(N__49851));
    Span4Mux_v I__9958 (
            .O(N__49851),
            .I(N__49848));
    Odrv4 I__9957 (
            .O(N__49848),
            .I(\c0.n39_adj_4295 ));
    InMux I__9956 (
            .O(N__49845),
            .I(N__49841));
    InMux I__9955 (
            .O(N__49844),
            .I(N__49838));
    LocalMux I__9954 (
            .O(N__49841),
            .I(N__49833));
    LocalMux I__9953 (
            .O(N__49838),
            .I(N__49833));
    Odrv4 I__9952 (
            .O(N__49833),
            .I(\c0.n13043 ));
    InMux I__9951 (
            .O(N__49830),
            .I(N__49824));
    InMux I__9950 (
            .O(N__49829),
            .I(N__49821));
    InMux I__9949 (
            .O(N__49828),
            .I(N__49818));
    InMux I__9948 (
            .O(N__49827),
            .I(N__49815));
    LocalMux I__9947 (
            .O(N__49824),
            .I(N__49812));
    LocalMux I__9946 (
            .O(N__49821),
            .I(N__49809));
    LocalMux I__9945 (
            .O(N__49818),
            .I(N__49806));
    LocalMux I__9944 (
            .O(N__49815),
            .I(N__49799));
    Span4Mux_v I__9943 (
            .O(N__49812),
            .I(N__49799));
    Span4Mux_v I__9942 (
            .O(N__49809),
            .I(N__49799));
    Odrv4 I__9941 (
            .O(N__49806),
            .I(\c0.n23912 ));
    Odrv4 I__9940 (
            .O(N__49799),
            .I(\c0.n23912 ));
    InMux I__9939 (
            .O(N__49794),
            .I(N__49788));
    InMux I__9938 (
            .O(N__49793),
            .I(N__49788));
    LocalMux I__9937 (
            .O(N__49788),
            .I(N__49783));
    InMux I__9936 (
            .O(N__49787),
            .I(N__49780));
    InMux I__9935 (
            .O(N__49786),
            .I(N__49777));
    Span4Mux_v I__9934 (
            .O(N__49783),
            .I(N__49774));
    LocalMux I__9933 (
            .O(N__49780),
            .I(N__49771));
    LocalMux I__9932 (
            .O(N__49777),
            .I(N__49768));
    Span4Mux_h I__9931 (
            .O(N__49774),
            .I(N__49765));
    Span4Mux_v I__9930 (
            .O(N__49771),
            .I(N__49762));
    Odrv4 I__9929 (
            .O(N__49768),
            .I(\c0.n35 ));
    Odrv4 I__9928 (
            .O(N__49765),
            .I(\c0.n35 ));
    Odrv4 I__9927 (
            .O(N__49762),
            .I(\c0.n35 ));
    CascadeMux I__9926 (
            .O(N__49755),
            .I(N__49752));
    InMux I__9925 (
            .O(N__49752),
            .I(N__49749));
    LocalMux I__9924 (
            .O(N__49749),
            .I(N__49746));
    Span4Mux_h I__9923 (
            .O(N__49746),
            .I(N__49743));
    Odrv4 I__9922 (
            .O(N__49743),
            .I(\c0.n22885 ));
    InMux I__9921 (
            .O(N__49740),
            .I(N__49737));
    LocalMux I__9920 (
            .O(N__49737),
            .I(N__49734));
    Span4Mux_s1_v I__9919 (
            .O(N__49734),
            .I(N__49731));
    Span4Mux_v I__9918 (
            .O(N__49731),
            .I(N__49727));
    CascadeMux I__9917 (
            .O(N__49730),
            .I(N__49724));
    Span4Mux_v I__9916 (
            .O(N__49727),
            .I(N__49719));
    InMux I__9915 (
            .O(N__49724),
            .I(N__49713));
    InMux I__9914 (
            .O(N__49723),
            .I(N__49713));
    InMux I__9913 (
            .O(N__49722),
            .I(N__49710));
    Span4Mux_v I__9912 (
            .O(N__49719),
            .I(N__49707));
    InMux I__9911 (
            .O(N__49718),
            .I(N__49704));
    LocalMux I__9910 (
            .O(N__49713),
            .I(N__49701));
    LocalMux I__9909 (
            .O(N__49710),
            .I(N__49698));
    Span4Mux_v I__9908 (
            .O(N__49707),
            .I(N__49693));
    LocalMux I__9907 (
            .O(N__49704),
            .I(N__49693));
    Span4Mux_v I__9906 (
            .O(N__49701),
            .I(N__49686));
    Span4Mux_v I__9905 (
            .O(N__49698),
            .I(N__49686));
    Span4Mux_h I__9904 (
            .O(N__49693),
            .I(N__49686));
    Span4Mux_h I__9903 (
            .O(N__49686),
            .I(N__49681));
    InMux I__9902 (
            .O(N__49685),
            .I(N__49678));
    InMux I__9901 (
            .O(N__49684),
            .I(N__49675));
    Span4Mux_h I__9900 (
            .O(N__49681),
            .I(N__49672));
    LocalMux I__9899 (
            .O(N__49678),
            .I(N__49669));
    LocalMux I__9898 (
            .O(N__49675),
            .I(r_Bit_Index_2));
    Odrv4 I__9897 (
            .O(N__49672),
            .I(r_Bit_Index_2));
    Odrv4 I__9896 (
            .O(N__49669),
            .I(r_Bit_Index_2));
    InMux I__9895 (
            .O(N__49662),
            .I(N__49659));
    LocalMux I__9894 (
            .O(N__49659),
            .I(N__49653));
    InMux I__9893 (
            .O(N__49658),
            .I(N__49650));
    InMux I__9892 (
            .O(N__49657),
            .I(N__49645));
    InMux I__9891 (
            .O(N__49656),
            .I(N__49642));
    Span4Mux_s1_v I__9890 (
            .O(N__49653),
            .I(N__49639));
    LocalMux I__9889 (
            .O(N__49650),
            .I(N__49635));
    InMux I__9888 (
            .O(N__49649),
            .I(N__49629));
    InMux I__9887 (
            .O(N__49648),
            .I(N__49629));
    LocalMux I__9886 (
            .O(N__49645),
            .I(N__49626));
    LocalMux I__9885 (
            .O(N__49642),
            .I(N__49623));
    Sp12to4 I__9884 (
            .O(N__49639),
            .I(N__49620));
    CascadeMux I__9883 (
            .O(N__49638),
            .I(N__49617));
    Span4Mux_v I__9882 (
            .O(N__49635),
            .I(N__49614));
    InMux I__9881 (
            .O(N__49634),
            .I(N__49611));
    LocalMux I__9880 (
            .O(N__49629),
            .I(N__49608));
    Span4Mux_h I__9879 (
            .O(N__49626),
            .I(N__49603));
    Span4Mux_h I__9878 (
            .O(N__49623),
            .I(N__49603));
    Span12Mux_h I__9877 (
            .O(N__49620),
            .I(N__49600));
    InMux I__9876 (
            .O(N__49617),
            .I(N__49597));
    Span4Mux_h I__9875 (
            .O(N__49614),
            .I(N__49592));
    LocalMux I__9874 (
            .O(N__49611),
            .I(N__49592));
    Span4Mux_h I__9873 (
            .O(N__49608),
            .I(N__49589));
    Span4Mux_h I__9872 (
            .O(N__49603),
            .I(N__49586));
    Span12Mux_v I__9871 (
            .O(N__49600),
            .I(N__49583));
    LocalMux I__9870 (
            .O(N__49597),
            .I(r_Bit_Index_1));
    Odrv4 I__9869 (
            .O(N__49592),
            .I(r_Bit_Index_1));
    Odrv4 I__9868 (
            .O(N__49589),
            .I(r_Bit_Index_1));
    Odrv4 I__9867 (
            .O(N__49586),
            .I(r_Bit_Index_1));
    Odrv12 I__9866 (
            .O(N__49583),
            .I(r_Bit_Index_1));
    InMux I__9865 (
            .O(N__49572),
            .I(N__49569));
    LocalMux I__9864 (
            .O(N__49569),
            .I(N__49566));
    Span12Mux_h I__9863 (
            .O(N__49566),
            .I(N__49563));
    Span12Mux_v I__9862 (
            .O(N__49563),
            .I(N__49560));
    Odrv12 I__9861 (
            .O(N__49560),
            .I(n4));
    CascadeMux I__9860 (
            .O(N__49557),
            .I(\c0.n20793_cascade_ ));
    InMux I__9859 (
            .O(N__49554),
            .I(N__49545));
    InMux I__9858 (
            .O(N__49553),
            .I(N__49545));
    InMux I__9857 (
            .O(N__49552),
            .I(N__49545));
    LocalMux I__9856 (
            .O(N__49545),
            .I(N__49542));
    Odrv4 I__9855 (
            .O(N__49542),
            .I(\c0.n12927 ));
    CascadeMux I__9854 (
            .O(N__49539),
            .I(\c0.n52_cascade_ ));
    CascadeMux I__9853 (
            .O(N__49536),
            .I(\c0.n47_adj_4537_cascade_ ));
    InMux I__9852 (
            .O(N__49533),
            .I(N__49530));
    LocalMux I__9851 (
            .O(N__49530),
            .I(N__49527));
    Odrv4 I__9850 (
            .O(N__49527),
            .I(\c0.n24581 ));
    CascadeMux I__9849 (
            .O(N__49524),
            .I(N__49520));
    CascadeMux I__9848 (
            .O(N__49523),
            .I(N__49517));
    InMux I__9847 (
            .O(N__49520),
            .I(N__49512));
    InMux I__9846 (
            .O(N__49517),
            .I(N__49512));
    LocalMux I__9845 (
            .O(N__49512),
            .I(\c0.data_in_frame_29_1 ));
    InMux I__9844 (
            .O(N__49509),
            .I(N__49503));
    InMux I__9843 (
            .O(N__49508),
            .I(N__49503));
    LocalMux I__9842 (
            .O(N__49503),
            .I(\c0.data_in_frame_29_6 ));
    InMux I__9841 (
            .O(N__49500),
            .I(N__49497));
    LocalMux I__9840 (
            .O(N__49497),
            .I(\c0.n20793 ));
    CascadeMux I__9839 (
            .O(N__49494),
            .I(N__49491));
    InMux I__9838 (
            .O(N__49491),
            .I(N__49488));
    LocalMux I__9837 (
            .O(N__49488),
            .I(N__49485));
    Span4Mux_h I__9836 (
            .O(N__49485),
            .I(N__49482));
    Sp12to4 I__9835 (
            .O(N__49482),
            .I(N__49479));
    Odrv12 I__9834 (
            .O(N__49479),
            .I(\c0.n5_adj_4302 ));
    CascadeMux I__9833 (
            .O(N__49476),
            .I(\c0.n12_adj_4348_cascade_ ));
    InMux I__9832 (
            .O(N__49473),
            .I(N__49470));
    LocalMux I__9831 (
            .O(N__49470),
            .I(\c0.n8_adj_4526 ));
    CascadeMux I__9830 (
            .O(N__49467),
            .I(\c0.n8_adj_4526_cascade_ ));
    InMux I__9829 (
            .O(N__49464),
            .I(N__49461));
    LocalMux I__9828 (
            .O(N__49461),
            .I(\c0.n9_adj_4536 ));
    InMux I__9827 (
            .O(N__49458),
            .I(N__49455));
    LocalMux I__9826 (
            .O(N__49455),
            .I(\c0.n14_adj_4528 ));
    InMux I__9825 (
            .O(N__49452),
            .I(N__49449));
    LocalMux I__9824 (
            .O(N__49449),
            .I(\c0.n14_adj_4576 ));
    InMux I__9823 (
            .O(N__49446),
            .I(N__49442));
    InMux I__9822 (
            .O(N__49445),
            .I(N__49439));
    LocalMux I__9821 (
            .O(N__49442),
            .I(\c0.data_in_frame_29_5 ));
    LocalMux I__9820 (
            .O(N__49439),
            .I(\c0.data_in_frame_29_5 ));
    CascadeMux I__9819 (
            .O(N__49434),
            .I(\c0.n24098_cascade_ ));
    InMux I__9818 (
            .O(N__49431),
            .I(N__49428));
    LocalMux I__9817 (
            .O(N__49428),
            .I(\c0.n10_adj_4484 ));
    InMux I__9816 (
            .O(N__49425),
            .I(N__49419));
    InMux I__9815 (
            .O(N__49424),
            .I(N__49416));
    InMux I__9814 (
            .O(N__49423),
            .I(N__49413));
    InMux I__9813 (
            .O(N__49422),
            .I(N__49410));
    LocalMux I__9812 (
            .O(N__49419),
            .I(N__49407));
    LocalMux I__9811 (
            .O(N__49416),
            .I(N__49402));
    LocalMux I__9810 (
            .O(N__49413),
            .I(N__49402));
    LocalMux I__9809 (
            .O(N__49410),
            .I(N__49397));
    Span4Mux_h I__9808 (
            .O(N__49407),
            .I(N__49397));
    Span4Mux_v I__9807 (
            .O(N__49402),
            .I(N__49394));
    Odrv4 I__9806 (
            .O(N__49397),
            .I(data_in_3_0));
    Odrv4 I__9805 (
            .O(N__49394),
            .I(data_in_3_0));
    InMux I__9804 (
            .O(N__49389),
            .I(N__49386));
    LocalMux I__9803 (
            .O(N__49386),
            .I(N__49382));
    InMux I__9802 (
            .O(N__49385),
            .I(N__49379));
    Span4Mux_v I__9801 (
            .O(N__49382),
            .I(N__49373));
    LocalMux I__9800 (
            .O(N__49379),
            .I(N__49373));
    InMux I__9799 (
            .O(N__49378),
            .I(N__49370));
    Span4Mux_v I__9798 (
            .O(N__49373),
            .I(N__49366));
    LocalMux I__9797 (
            .O(N__49370),
            .I(N__49363));
    InMux I__9796 (
            .O(N__49369),
            .I(N__49360));
    Span4Mux_v I__9795 (
            .O(N__49366),
            .I(N__49353));
    Span4Mux_h I__9794 (
            .O(N__49363),
            .I(N__49353));
    LocalMux I__9793 (
            .O(N__49360),
            .I(N__49353));
    Odrv4 I__9792 (
            .O(N__49353),
            .I(n12981));
    InMux I__9791 (
            .O(N__49350),
            .I(N__49344));
    InMux I__9790 (
            .O(N__49349),
            .I(N__49344));
    LocalMux I__9789 (
            .O(N__49344),
            .I(N__49341));
    Span4Mux_h I__9788 (
            .O(N__49341),
            .I(N__49338));
    Span4Mux_h I__9787 (
            .O(N__49338),
            .I(N__49335));
    Odrv4 I__9786 (
            .O(N__49335),
            .I(n4_adj_4762));
    InMux I__9785 (
            .O(N__49332),
            .I(N__49329));
    LocalMux I__9784 (
            .O(N__49329),
            .I(N__49326));
    Odrv4 I__9783 (
            .O(N__49326),
            .I(\c0.n22716 ));
    CascadeMux I__9782 (
            .O(N__49323),
            .I(\c0.n22716_cascade_ ));
    InMux I__9781 (
            .O(N__49320),
            .I(N__49317));
    LocalMux I__9780 (
            .O(N__49317),
            .I(\c0.n8_adj_4248 ));
    CascadeMux I__9779 (
            .O(N__49314),
            .I(N__49311));
    InMux I__9778 (
            .O(N__49311),
            .I(N__49307));
    InMux I__9777 (
            .O(N__49310),
            .I(N__49304));
    LocalMux I__9776 (
            .O(N__49307),
            .I(N__49299));
    LocalMux I__9775 (
            .O(N__49304),
            .I(N__49296));
    InMux I__9774 (
            .O(N__49303),
            .I(N__49293));
    InMux I__9773 (
            .O(N__49302),
            .I(N__49290));
    Span4Mux_h I__9772 (
            .O(N__49299),
            .I(N__49287));
    Span4Mux_h I__9771 (
            .O(N__49296),
            .I(N__49284));
    LocalMux I__9770 (
            .O(N__49293),
            .I(N__49281));
    LocalMux I__9769 (
            .O(N__49290),
            .I(data_in_3_1));
    Odrv4 I__9768 (
            .O(N__49287),
            .I(data_in_3_1));
    Odrv4 I__9767 (
            .O(N__49284),
            .I(data_in_3_1));
    Odrv12 I__9766 (
            .O(N__49281),
            .I(data_in_3_1));
    InMux I__9765 (
            .O(N__49272),
            .I(N__49269));
    LocalMux I__9764 (
            .O(N__49269),
            .I(N__49265));
    CascadeMux I__9763 (
            .O(N__49268),
            .I(N__49261));
    Span4Mux_v I__9762 (
            .O(N__49265),
            .I(N__49257));
    InMux I__9761 (
            .O(N__49264),
            .I(N__49254));
    InMux I__9760 (
            .O(N__49261),
            .I(N__49249));
    InMux I__9759 (
            .O(N__49260),
            .I(N__49249));
    Odrv4 I__9758 (
            .O(N__49257),
            .I(data_in_1_2));
    LocalMux I__9757 (
            .O(N__49254),
            .I(data_in_1_2));
    LocalMux I__9756 (
            .O(N__49249),
            .I(data_in_1_2));
    InMux I__9755 (
            .O(N__49242),
            .I(N__49239));
    LocalMux I__9754 (
            .O(N__49239),
            .I(N__49234));
    InMux I__9753 (
            .O(N__49238),
            .I(N__49231));
    InMux I__9752 (
            .O(N__49237),
            .I(N__49228));
    Span4Mux_h I__9751 (
            .O(N__49234),
            .I(N__49225));
    LocalMux I__9750 (
            .O(N__49231),
            .I(N__49222));
    LocalMux I__9749 (
            .O(N__49228),
            .I(data_in_0_2));
    Odrv4 I__9748 (
            .O(N__49225),
            .I(data_in_0_2));
    Odrv12 I__9747 (
            .O(N__49222),
            .I(data_in_0_2));
    CascadeMux I__9746 (
            .O(N__49215),
            .I(N__49212));
    InMux I__9745 (
            .O(N__49212),
            .I(N__49209));
    LocalMux I__9744 (
            .O(N__49209),
            .I(\c0.n10_adj_4732 ));
    CascadeMux I__9743 (
            .O(N__49206),
            .I(\c0.n26_adj_4733_cascade_ ));
    CascadeMux I__9742 (
            .O(N__49203),
            .I(\c0.n20409_cascade_ ));
    InMux I__9741 (
            .O(N__49200),
            .I(N__49197));
    LocalMux I__9740 (
            .O(N__49197),
            .I(N__49193));
    InMux I__9739 (
            .O(N__49196),
            .I(N__49190));
    Span4Mux_h I__9738 (
            .O(N__49193),
            .I(N__49187));
    LocalMux I__9737 (
            .O(N__49190),
            .I(N__49181));
    Span4Mux_h I__9736 (
            .O(N__49187),
            .I(N__49181));
    InMux I__9735 (
            .O(N__49186),
            .I(N__49178));
    Span4Mux_v I__9734 (
            .O(N__49181),
            .I(N__49175));
    LocalMux I__9733 (
            .O(N__49178),
            .I(\c0.FRAME_MATCHER_state_7 ));
    Odrv4 I__9732 (
            .O(N__49175),
            .I(\c0.FRAME_MATCHER_state_7 ));
    SRMux I__9731 (
            .O(N__49170),
            .I(N__49167));
    LocalMux I__9730 (
            .O(N__49167),
            .I(N__49164));
    Span4Mux_h I__9729 (
            .O(N__49164),
            .I(N__49161));
    Span4Mux_v I__9728 (
            .O(N__49161),
            .I(N__49158));
    Odrv4 I__9727 (
            .O(N__49158),
            .I(\c0.n21629 ));
    InMux I__9726 (
            .O(N__49155),
            .I(N__49152));
    LocalMux I__9725 (
            .O(N__49152),
            .I(N__49149));
    Span4Mux_h I__9724 (
            .O(N__49149),
            .I(N__49146));
    Odrv4 I__9723 (
            .O(N__49146),
            .I(\c0.n25_adj_4723 ));
    InMux I__9722 (
            .O(N__49143),
            .I(N__49140));
    LocalMux I__9721 (
            .O(N__49140),
            .I(N__49136));
    CascadeMux I__9720 (
            .O(N__49139),
            .I(N__49133));
    Span4Mux_v I__9719 (
            .O(N__49136),
            .I(N__49130));
    InMux I__9718 (
            .O(N__49133),
            .I(N__49126));
    Span4Mux_h I__9717 (
            .O(N__49130),
            .I(N__49123));
    InMux I__9716 (
            .O(N__49129),
            .I(N__49120));
    LocalMux I__9715 (
            .O(N__49126),
            .I(N__49117));
    Sp12to4 I__9714 (
            .O(N__49123),
            .I(N__49114));
    LocalMux I__9713 (
            .O(N__49120),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv4 I__9712 (
            .O(N__49117),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv12 I__9711 (
            .O(N__49114),
            .I(\c0.FRAME_MATCHER_state_19 ));
    InMux I__9710 (
            .O(N__49107),
            .I(N__49104));
    LocalMux I__9709 (
            .O(N__49104),
            .I(N__49099));
    InMux I__9708 (
            .O(N__49103),
            .I(N__49096));
    InMux I__9707 (
            .O(N__49102),
            .I(N__49093));
    Span12Mux_h I__9706 (
            .O(N__49099),
            .I(N__49090));
    LocalMux I__9705 (
            .O(N__49096),
            .I(\c0.FRAME_MATCHER_state_23 ));
    LocalMux I__9704 (
            .O(N__49093),
            .I(\c0.FRAME_MATCHER_state_23 ));
    Odrv12 I__9703 (
            .O(N__49090),
            .I(\c0.FRAME_MATCHER_state_23 ));
    CascadeMux I__9702 (
            .O(N__49083),
            .I(N__49080));
    InMux I__9701 (
            .O(N__49080),
            .I(N__49077));
    LocalMux I__9700 (
            .O(N__49077),
            .I(N__49074));
    Span4Mux_v I__9699 (
            .O(N__49074),
            .I(N__49070));
    InMux I__9698 (
            .O(N__49073),
            .I(N__49066));
    Span4Mux_h I__9697 (
            .O(N__49070),
            .I(N__49063));
    InMux I__9696 (
            .O(N__49069),
            .I(N__49060));
    LocalMux I__9695 (
            .O(N__49066),
            .I(N__49057));
    Sp12to4 I__9694 (
            .O(N__49063),
            .I(N__49054));
    LocalMux I__9693 (
            .O(N__49060),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv4 I__9692 (
            .O(N__49057),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv12 I__9691 (
            .O(N__49054),
            .I(\c0.FRAME_MATCHER_state_21 ));
    InMux I__9690 (
            .O(N__49047),
            .I(N__49044));
    LocalMux I__9689 (
            .O(N__49044),
            .I(N__49040));
    InMux I__9688 (
            .O(N__49043),
            .I(N__49037));
    Span4Mux_v I__9687 (
            .O(N__49040),
            .I(N__49033));
    LocalMux I__9686 (
            .O(N__49037),
            .I(N__49030));
    InMux I__9685 (
            .O(N__49036),
            .I(N__49027));
    Span4Mux_v I__9684 (
            .O(N__49033),
            .I(N__49024));
    Sp12to4 I__9683 (
            .O(N__49030),
            .I(N__49019));
    LocalMux I__9682 (
            .O(N__49027),
            .I(N__49019));
    Sp12to4 I__9681 (
            .O(N__49024),
            .I(N__49014));
    Span12Mux_v I__9680 (
            .O(N__49019),
            .I(N__49014));
    Odrv12 I__9679 (
            .O(N__49014),
            .I(\c0.n22049 ));
    InMux I__9678 (
            .O(N__49011),
            .I(N__49008));
    LocalMux I__9677 (
            .O(N__49008),
            .I(N__49004));
    InMux I__9676 (
            .O(N__49007),
            .I(N__49000));
    Span4Mux_h I__9675 (
            .O(N__49004),
            .I(N__48996));
    InMux I__9674 (
            .O(N__49003),
            .I(N__48993));
    LocalMux I__9673 (
            .O(N__49000),
            .I(N__48981));
    InMux I__9672 (
            .O(N__48999),
            .I(N__48975));
    Span4Mux_v I__9671 (
            .O(N__48996),
            .I(N__48970));
    LocalMux I__9670 (
            .O(N__48993),
            .I(N__48970));
    InMux I__9669 (
            .O(N__48992),
            .I(N__48966));
    InMux I__9668 (
            .O(N__48991),
            .I(N__48963));
    InMux I__9667 (
            .O(N__48990),
            .I(N__48957));
    InMux I__9666 (
            .O(N__48989),
            .I(N__48954));
    InMux I__9665 (
            .O(N__48988),
            .I(N__48951));
    InMux I__9664 (
            .O(N__48987),
            .I(N__48948));
    InMux I__9663 (
            .O(N__48986),
            .I(N__48945));
    InMux I__9662 (
            .O(N__48985),
            .I(N__48942));
    InMux I__9661 (
            .O(N__48984),
            .I(N__48938));
    Span4Mux_v I__9660 (
            .O(N__48981),
            .I(N__48935));
    InMux I__9659 (
            .O(N__48980),
            .I(N__48932));
    InMux I__9658 (
            .O(N__48979),
            .I(N__48929));
    InMux I__9657 (
            .O(N__48978),
            .I(N__48925));
    LocalMux I__9656 (
            .O(N__48975),
            .I(N__48922));
    Span4Mux_v I__9655 (
            .O(N__48970),
            .I(N__48919));
    InMux I__9654 (
            .O(N__48969),
            .I(N__48916));
    LocalMux I__9653 (
            .O(N__48966),
            .I(N__48911));
    LocalMux I__9652 (
            .O(N__48963),
            .I(N__48911));
    InMux I__9651 (
            .O(N__48962),
            .I(N__48908));
    InMux I__9650 (
            .O(N__48961),
            .I(N__48905));
    InMux I__9649 (
            .O(N__48960),
            .I(N__48902));
    LocalMux I__9648 (
            .O(N__48957),
            .I(N__48889));
    LocalMux I__9647 (
            .O(N__48954),
            .I(N__48889));
    LocalMux I__9646 (
            .O(N__48951),
            .I(N__48889));
    LocalMux I__9645 (
            .O(N__48948),
            .I(N__48889));
    LocalMux I__9644 (
            .O(N__48945),
            .I(N__48889));
    LocalMux I__9643 (
            .O(N__48942),
            .I(N__48889));
    InMux I__9642 (
            .O(N__48941),
            .I(N__48886));
    LocalMux I__9641 (
            .O(N__48938),
            .I(N__48883));
    Span4Mux_h I__9640 (
            .O(N__48935),
            .I(N__48879));
    LocalMux I__9639 (
            .O(N__48932),
            .I(N__48874));
    LocalMux I__9638 (
            .O(N__48929),
            .I(N__48874));
    InMux I__9637 (
            .O(N__48928),
            .I(N__48871));
    LocalMux I__9636 (
            .O(N__48925),
            .I(N__48867));
    Span4Mux_h I__9635 (
            .O(N__48922),
            .I(N__48860));
    Span4Mux_h I__9634 (
            .O(N__48919),
            .I(N__48860));
    LocalMux I__9633 (
            .O(N__48916),
            .I(N__48860));
    Span4Mux_h I__9632 (
            .O(N__48911),
            .I(N__48853));
    LocalMux I__9631 (
            .O(N__48908),
            .I(N__48853));
    LocalMux I__9630 (
            .O(N__48905),
            .I(N__48853));
    LocalMux I__9629 (
            .O(N__48902),
            .I(N__48850));
    Span4Mux_v I__9628 (
            .O(N__48889),
            .I(N__48845));
    LocalMux I__9627 (
            .O(N__48886),
            .I(N__48845));
    Span12Mux_h I__9626 (
            .O(N__48883),
            .I(N__48842));
    InMux I__9625 (
            .O(N__48882),
            .I(N__48839));
    Span4Mux_h I__9624 (
            .O(N__48879),
            .I(N__48834));
    Span4Mux_h I__9623 (
            .O(N__48874),
            .I(N__48829));
    LocalMux I__9622 (
            .O(N__48871),
            .I(N__48829));
    InMux I__9621 (
            .O(N__48870),
            .I(N__48826));
    Span12Mux_v I__9620 (
            .O(N__48867),
            .I(N__48821));
    Span4Mux_v I__9619 (
            .O(N__48860),
            .I(N__48814));
    Span4Mux_v I__9618 (
            .O(N__48853),
            .I(N__48814));
    Span4Mux_v I__9617 (
            .O(N__48850),
            .I(N__48814));
    Span4Mux_h I__9616 (
            .O(N__48845),
            .I(N__48811));
    Span12Mux_v I__9615 (
            .O(N__48842),
            .I(N__48806));
    LocalMux I__9614 (
            .O(N__48839),
            .I(N__48806));
    InMux I__9613 (
            .O(N__48838),
            .I(N__48803));
    InMux I__9612 (
            .O(N__48837),
            .I(N__48800));
    Span4Mux_v I__9611 (
            .O(N__48834),
            .I(N__48793));
    Span4Mux_h I__9610 (
            .O(N__48829),
            .I(N__48793));
    LocalMux I__9609 (
            .O(N__48826),
            .I(N__48793));
    InMux I__9608 (
            .O(N__48825),
            .I(N__48790));
    InMux I__9607 (
            .O(N__48824),
            .I(N__48787));
    Odrv12 I__9606 (
            .O(N__48821),
            .I(\c0.n5 ));
    Odrv4 I__9605 (
            .O(N__48814),
            .I(\c0.n5 ));
    Odrv4 I__9604 (
            .O(N__48811),
            .I(\c0.n5 ));
    Odrv12 I__9603 (
            .O(N__48806),
            .I(\c0.n5 ));
    LocalMux I__9602 (
            .O(N__48803),
            .I(\c0.n5 ));
    LocalMux I__9601 (
            .O(N__48800),
            .I(\c0.n5 ));
    Odrv4 I__9600 (
            .O(N__48793),
            .I(\c0.n5 ));
    LocalMux I__9599 (
            .O(N__48790),
            .I(\c0.n5 ));
    LocalMux I__9598 (
            .O(N__48787),
            .I(\c0.n5 ));
    InMux I__9597 (
            .O(N__48768),
            .I(N__48763));
    InMux I__9596 (
            .O(N__48767),
            .I(N__48758));
    InMux I__9595 (
            .O(N__48766),
            .I(N__48758));
    LocalMux I__9594 (
            .O(N__48763),
            .I(\c0.FRAME_MATCHER_state_27 ));
    LocalMux I__9593 (
            .O(N__48758),
            .I(\c0.FRAME_MATCHER_state_27 ));
    SRMux I__9592 (
            .O(N__48753),
            .I(N__48750));
    LocalMux I__9591 (
            .O(N__48750),
            .I(N__48747));
    Odrv4 I__9590 (
            .O(N__48747),
            .I(\c0.n21647 ));
    InMux I__9589 (
            .O(N__48744),
            .I(N__48740));
    InMux I__9588 (
            .O(N__48743),
            .I(N__48736));
    LocalMux I__9587 (
            .O(N__48740),
            .I(N__48733));
    InMux I__9586 (
            .O(N__48739),
            .I(N__48728));
    LocalMux I__9585 (
            .O(N__48736),
            .I(N__48723));
    Span4Mux_v I__9584 (
            .O(N__48733),
            .I(N__48723));
    InMux I__9583 (
            .O(N__48732),
            .I(N__48718));
    InMux I__9582 (
            .O(N__48731),
            .I(N__48718));
    LocalMux I__9581 (
            .O(N__48728),
            .I(data_in_frame_5_6));
    Odrv4 I__9580 (
            .O(N__48723),
            .I(data_in_frame_5_6));
    LocalMux I__9579 (
            .O(N__48718),
            .I(data_in_frame_5_6));
    CascadeMux I__9578 (
            .O(N__48711),
            .I(N__48707));
    InMux I__9577 (
            .O(N__48710),
            .I(N__48704));
    InMux I__9576 (
            .O(N__48707),
            .I(N__48701));
    LocalMux I__9575 (
            .O(N__48704),
            .I(N__48698));
    LocalMux I__9574 (
            .O(N__48701),
            .I(N__48692));
    Span4Mux_v I__9573 (
            .O(N__48698),
            .I(N__48692));
    InMux I__9572 (
            .O(N__48697),
            .I(N__48689));
    Odrv4 I__9571 (
            .O(N__48692),
            .I(\c0.data_in_frame_7_7 ));
    LocalMux I__9570 (
            .O(N__48689),
            .I(\c0.data_in_frame_7_7 ));
    CascadeMux I__9569 (
            .O(N__48684),
            .I(N__48681));
    InMux I__9568 (
            .O(N__48681),
            .I(N__48676));
    InMux I__9567 (
            .O(N__48680),
            .I(N__48673));
    InMux I__9566 (
            .O(N__48679),
            .I(N__48670));
    LocalMux I__9565 (
            .O(N__48676),
            .I(N__48667));
    LocalMux I__9564 (
            .O(N__48673),
            .I(N__48663));
    LocalMux I__9563 (
            .O(N__48670),
            .I(N__48660));
    Span4Mux_v I__9562 (
            .O(N__48667),
            .I(N__48657));
    InMux I__9561 (
            .O(N__48666),
            .I(N__48654));
    Span12Mux_h I__9560 (
            .O(N__48663),
            .I(N__48651));
    Span4Mux_v I__9559 (
            .O(N__48660),
            .I(N__48648));
    Span4Mux_h I__9558 (
            .O(N__48657),
            .I(N__48645));
    LocalMux I__9557 (
            .O(N__48654),
            .I(data_in_3_3));
    Odrv12 I__9556 (
            .O(N__48651),
            .I(data_in_3_3));
    Odrv4 I__9555 (
            .O(N__48648),
            .I(data_in_3_3));
    Odrv4 I__9554 (
            .O(N__48645),
            .I(data_in_3_3));
    InMux I__9553 (
            .O(N__48636),
            .I(N__48633));
    LocalMux I__9552 (
            .O(N__48633),
            .I(N__48629));
    InMux I__9551 (
            .O(N__48632),
            .I(N__48625));
    Span4Mux_v I__9550 (
            .O(N__48629),
            .I(N__48622));
    InMux I__9549 (
            .O(N__48628),
            .I(N__48619));
    LocalMux I__9548 (
            .O(N__48625),
            .I(N__48616));
    Span4Mux_h I__9547 (
            .O(N__48622),
            .I(N__48613));
    LocalMux I__9546 (
            .O(N__48619),
            .I(data_in_0_7));
    Odrv4 I__9545 (
            .O(N__48616),
            .I(data_in_0_7));
    Odrv4 I__9544 (
            .O(N__48613),
            .I(data_in_0_7));
    InMux I__9543 (
            .O(N__48606),
            .I(N__48603));
    LocalMux I__9542 (
            .O(N__48603),
            .I(N__48600));
    Span4Mux_v I__9541 (
            .O(N__48600),
            .I(N__48597));
    Odrv4 I__9540 (
            .O(N__48597),
            .I(\c0.n14 ));
    InMux I__9539 (
            .O(N__48594),
            .I(N__48591));
    LocalMux I__9538 (
            .O(N__48591),
            .I(\c0.n20_adj_4729 ));
    CascadeMux I__9537 (
            .O(N__48588),
            .I(N__48585));
    InMux I__9536 (
            .O(N__48585),
            .I(N__48582));
    LocalMux I__9535 (
            .O(N__48582),
            .I(\c0.n6_adj_4704 ));
    CascadeMux I__9534 (
            .O(N__48579),
            .I(\c0.n14016_cascade_ ));
    CascadeMux I__9533 (
            .O(N__48576),
            .I(\c0.n20_cascade_ ));
    CascadeMux I__9532 (
            .O(N__48573),
            .I(\c0.n6_adj_4254_cascade_ ));
    InMux I__9531 (
            .O(N__48570),
            .I(N__48567));
    LocalMux I__9530 (
            .O(N__48567),
            .I(N__48564));
    Span4Mux_h I__9529 (
            .O(N__48564),
            .I(N__48561));
    Odrv4 I__9528 (
            .O(N__48561),
            .I(\c0.n28_adj_4731 ));
    CascadeMux I__9527 (
            .O(N__48558),
            .I(\c0.n14_adj_4607_cascade_ ));
    InMux I__9526 (
            .O(N__48555),
            .I(N__48549));
    InMux I__9525 (
            .O(N__48554),
            .I(N__48549));
    LocalMux I__9524 (
            .O(N__48549),
            .I(\c0.n22626 ));
    CascadeMux I__9523 (
            .O(N__48546),
            .I(\c0.data_out_frame_0__7__N_2626_cascade_ ));
    InMux I__9522 (
            .O(N__48543),
            .I(N__48537));
    InMux I__9521 (
            .O(N__48542),
            .I(N__48537));
    LocalMux I__9520 (
            .O(N__48537),
            .I(\c0.n30_adj_4585 ));
    InMux I__9519 (
            .O(N__48534),
            .I(N__48531));
    LocalMux I__9518 (
            .O(N__48531),
            .I(\c0.n20_adj_4642 ));
    CascadeMux I__9517 (
            .O(N__48528),
            .I(N__48525));
    InMux I__9516 (
            .O(N__48525),
            .I(N__48522));
    LocalMux I__9515 (
            .O(N__48522),
            .I(\c0.n4_adj_4266 ));
    CascadeMux I__9514 (
            .O(N__48519),
            .I(N__48516));
    InMux I__9513 (
            .O(N__48516),
            .I(N__48512));
    CascadeMux I__9512 (
            .O(N__48515),
            .I(N__48507));
    LocalMux I__9511 (
            .O(N__48512),
            .I(N__48504));
    InMux I__9510 (
            .O(N__48511),
            .I(N__48501));
    InMux I__9509 (
            .O(N__48510),
            .I(N__48496));
    InMux I__9508 (
            .O(N__48507),
            .I(N__48496));
    Span4Mux_v I__9507 (
            .O(N__48504),
            .I(N__48493));
    LocalMux I__9506 (
            .O(N__48501),
            .I(N__48486));
    LocalMux I__9505 (
            .O(N__48496),
            .I(N__48486));
    Sp12to4 I__9504 (
            .O(N__48493),
            .I(N__48486));
    Odrv12 I__9503 (
            .O(N__48486),
            .I(\c0.n5024 ));
    InMux I__9502 (
            .O(N__48483),
            .I(N__48479));
    InMux I__9501 (
            .O(N__48482),
            .I(N__48476));
    LocalMux I__9500 (
            .O(N__48479),
            .I(N__48472));
    LocalMux I__9499 (
            .O(N__48476),
            .I(N__48469));
    InMux I__9498 (
            .O(N__48475),
            .I(N__48466));
    Span4Mux_v I__9497 (
            .O(N__48472),
            .I(N__48463));
    Span4Mux_h I__9496 (
            .O(N__48469),
            .I(N__48460));
    LocalMux I__9495 (
            .O(N__48466),
            .I(N__48457));
    Odrv4 I__9494 (
            .O(N__48463),
            .I(\c0.n12992 ));
    Odrv4 I__9493 (
            .O(N__48460),
            .I(\c0.n12992 ));
    Odrv12 I__9492 (
            .O(N__48457),
            .I(\c0.n12992 ));
    InMux I__9491 (
            .O(N__48450),
            .I(N__48447));
    LocalMux I__9490 (
            .O(N__48447),
            .I(N__48444));
    Span4Mux_h I__9489 (
            .O(N__48444),
            .I(N__48440));
    InMux I__9488 (
            .O(N__48443),
            .I(N__48437));
    Odrv4 I__9487 (
            .O(N__48440),
            .I(\c0.n13052 ));
    LocalMux I__9486 (
            .O(N__48437),
            .I(\c0.n13052 ));
    CascadeMux I__9485 (
            .O(N__48432),
            .I(N__48429));
    InMux I__9484 (
            .O(N__48429),
            .I(N__48426));
    LocalMux I__9483 (
            .O(N__48426),
            .I(N__48423));
    Odrv4 I__9482 (
            .O(N__48423),
            .I(\c0.n24736 ));
    InMux I__9481 (
            .O(N__48420),
            .I(N__48417));
    LocalMux I__9480 (
            .O(N__48417),
            .I(N__48413));
    InMux I__9479 (
            .O(N__48416),
            .I(N__48409));
    Span4Mux_v I__9478 (
            .O(N__48413),
            .I(N__48406));
    InMux I__9477 (
            .O(N__48412),
            .I(N__48403));
    LocalMux I__9476 (
            .O(N__48409),
            .I(N__48400));
    Span4Mux_h I__9475 (
            .O(N__48406),
            .I(N__48397));
    LocalMux I__9474 (
            .O(N__48403),
            .I(\c0.FRAME_MATCHER_state_31 ));
    Odrv4 I__9473 (
            .O(N__48400),
            .I(\c0.FRAME_MATCHER_state_31 ));
    Odrv4 I__9472 (
            .O(N__48397),
            .I(\c0.FRAME_MATCHER_state_31 ));
    SRMux I__9471 (
            .O(N__48390),
            .I(N__48387));
    LocalMux I__9470 (
            .O(N__48387),
            .I(N__48384));
    Odrv4 I__9469 (
            .O(N__48384),
            .I(\c0.n21651 ));
    CascadeMux I__9468 (
            .O(N__48381),
            .I(N__48369));
    CascadeMux I__9467 (
            .O(N__48380),
            .I(N__48366));
    InMux I__9466 (
            .O(N__48379),
            .I(N__48359));
    CascadeMux I__9465 (
            .O(N__48378),
            .I(N__48356));
    CascadeMux I__9464 (
            .O(N__48377),
            .I(N__48353));
    InMux I__9463 (
            .O(N__48376),
            .I(N__48350));
    InMux I__9462 (
            .O(N__48375),
            .I(N__48338));
    InMux I__9461 (
            .O(N__48374),
            .I(N__48338));
    InMux I__9460 (
            .O(N__48373),
            .I(N__48338));
    InMux I__9459 (
            .O(N__48372),
            .I(N__48335));
    InMux I__9458 (
            .O(N__48369),
            .I(N__48330));
    InMux I__9457 (
            .O(N__48366),
            .I(N__48330));
    InMux I__9456 (
            .O(N__48365),
            .I(N__48325));
    InMux I__9455 (
            .O(N__48364),
            .I(N__48325));
    InMux I__9454 (
            .O(N__48363),
            .I(N__48316));
    InMux I__9453 (
            .O(N__48362),
            .I(N__48313));
    LocalMux I__9452 (
            .O(N__48359),
            .I(N__48310));
    InMux I__9451 (
            .O(N__48356),
            .I(N__48305));
    InMux I__9450 (
            .O(N__48353),
            .I(N__48305));
    LocalMux I__9449 (
            .O(N__48350),
            .I(N__48302));
    InMux I__9448 (
            .O(N__48349),
            .I(N__48295));
    InMux I__9447 (
            .O(N__48348),
            .I(N__48295));
    InMux I__9446 (
            .O(N__48347),
            .I(N__48295));
    InMux I__9445 (
            .O(N__48346),
            .I(N__48288));
    InMux I__9444 (
            .O(N__48345),
            .I(N__48288));
    LocalMux I__9443 (
            .O(N__48338),
            .I(N__48283));
    LocalMux I__9442 (
            .O(N__48335),
            .I(N__48283));
    LocalMux I__9441 (
            .O(N__48330),
            .I(N__48278));
    LocalMux I__9440 (
            .O(N__48325),
            .I(N__48278));
    CascadeMux I__9439 (
            .O(N__48324),
            .I(N__48275));
    CascadeMux I__9438 (
            .O(N__48323),
            .I(N__48272));
    InMux I__9437 (
            .O(N__48322),
            .I(N__48260));
    InMux I__9436 (
            .O(N__48321),
            .I(N__48260));
    InMux I__9435 (
            .O(N__48320),
            .I(N__48260));
    InMux I__9434 (
            .O(N__48319),
            .I(N__48260));
    LocalMux I__9433 (
            .O(N__48316),
            .I(N__48257));
    LocalMux I__9432 (
            .O(N__48313),
            .I(N__48227));
    Span4Mux_h I__9431 (
            .O(N__48310),
            .I(N__48227));
    LocalMux I__9430 (
            .O(N__48305),
            .I(N__48227));
    Span4Mux_v I__9429 (
            .O(N__48302),
            .I(N__48227));
    LocalMux I__9428 (
            .O(N__48295),
            .I(N__48227));
    InMux I__9427 (
            .O(N__48294),
            .I(N__48222));
    InMux I__9426 (
            .O(N__48293),
            .I(N__48222));
    LocalMux I__9425 (
            .O(N__48288),
            .I(N__48215));
    Span4Mux_v I__9424 (
            .O(N__48283),
            .I(N__48215));
    Span4Mux_v I__9423 (
            .O(N__48278),
            .I(N__48215));
    InMux I__9422 (
            .O(N__48275),
            .I(N__48210));
    InMux I__9421 (
            .O(N__48272),
            .I(N__48210));
    InMux I__9420 (
            .O(N__48271),
            .I(N__48197));
    InMux I__9419 (
            .O(N__48270),
            .I(N__48194));
    CascadeMux I__9418 (
            .O(N__48269),
            .I(N__48191));
    LocalMux I__9417 (
            .O(N__48260),
            .I(N__48182));
    Span4Mux_v I__9416 (
            .O(N__48257),
            .I(N__48179));
    InMux I__9415 (
            .O(N__48256),
            .I(N__48176));
    InMux I__9414 (
            .O(N__48255),
            .I(N__48169));
    InMux I__9413 (
            .O(N__48254),
            .I(N__48169));
    InMux I__9412 (
            .O(N__48253),
            .I(N__48169));
    InMux I__9411 (
            .O(N__48252),
            .I(N__48162));
    InMux I__9410 (
            .O(N__48251),
            .I(N__48162));
    InMux I__9409 (
            .O(N__48250),
            .I(N__48162));
    InMux I__9408 (
            .O(N__48249),
            .I(N__48159));
    InMux I__9407 (
            .O(N__48248),
            .I(N__48154));
    InMux I__9406 (
            .O(N__48247),
            .I(N__48154));
    InMux I__9405 (
            .O(N__48246),
            .I(N__48143));
    InMux I__9404 (
            .O(N__48245),
            .I(N__48143));
    InMux I__9403 (
            .O(N__48244),
            .I(N__48143));
    InMux I__9402 (
            .O(N__48243),
            .I(N__48143));
    InMux I__9401 (
            .O(N__48242),
            .I(N__48143));
    CascadeMux I__9400 (
            .O(N__48241),
            .I(N__48138));
    CascadeMux I__9399 (
            .O(N__48240),
            .I(N__48135));
    InMux I__9398 (
            .O(N__48239),
            .I(N__48126));
    InMux I__9397 (
            .O(N__48238),
            .I(N__48126));
    Span4Mux_v I__9396 (
            .O(N__48227),
            .I(N__48117));
    LocalMux I__9395 (
            .O(N__48222),
            .I(N__48117));
    Span4Mux_h I__9394 (
            .O(N__48215),
            .I(N__48117));
    LocalMux I__9393 (
            .O(N__48210),
            .I(N__48117));
    InMux I__9392 (
            .O(N__48209),
            .I(N__48108));
    InMux I__9391 (
            .O(N__48208),
            .I(N__48108));
    InMux I__9390 (
            .O(N__48207),
            .I(N__48108));
    InMux I__9389 (
            .O(N__48206),
            .I(N__48108));
    InMux I__9388 (
            .O(N__48205),
            .I(N__48099));
    InMux I__9387 (
            .O(N__48204),
            .I(N__48099));
    InMux I__9386 (
            .O(N__48203),
            .I(N__48099));
    InMux I__9385 (
            .O(N__48202),
            .I(N__48099));
    InMux I__9384 (
            .O(N__48201),
            .I(N__48094));
    InMux I__9383 (
            .O(N__48200),
            .I(N__48094));
    LocalMux I__9382 (
            .O(N__48197),
            .I(N__48091));
    LocalMux I__9381 (
            .O(N__48194),
            .I(N__48088));
    InMux I__9380 (
            .O(N__48191),
            .I(N__48078));
    InMux I__9379 (
            .O(N__48190),
            .I(N__48078));
    InMux I__9378 (
            .O(N__48189),
            .I(N__48078));
    InMux I__9377 (
            .O(N__48188),
            .I(N__48072));
    InMux I__9376 (
            .O(N__48187),
            .I(N__48072));
    InMux I__9375 (
            .O(N__48186),
            .I(N__48069));
    InMux I__9374 (
            .O(N__48185),
            .I(N__48064));
    Span4Mux_v I__9373 (
            .O(N__48182),
            .I(N__48047));
    Span4Mux_h I__9372 (
            .O(N__48179),
            .I(N__48047));
    LocalMux I__9371 (
            .O(N__48176),
            .I(N__48047));
    LocalMux I__9370 (
            .O(N__48169),
            .I(N__48047));
    LocalMux I__9369 (
            .O(N__48162),
            .I(N__48047));
    LocalMux I__9368 (
            .O(N__48159),
            .I(N__48047));
    LocalMux I__9367 (
            .O(N__48154),
            .I(N__48047));
    LocalMux I__9366 (
            .O(N__48143),
            .I(N__48047));
    InMux I__9365 (
            .O(N__48142),
            .I(N__48036));
    InMux I__9364 (
            .O(N__48141),
            .I(N__48036));
    InMux I__9363 (
            .O(N__48138),
            .I(N__48036));
    InMux I__9362 (
            .O(N__48135),
            .I(N__48036));
    InMux I__9361 (
            .O(N__48134),
            .I(N__48036));
    InMux I__9360 (
            .O(N__48133),
            .I(N__48029));
    InMux I__9359 (
            .O(N__48132),
            .I(N__48029));
    InMux I__9358 (
            .O(N__48131),
            .I(N__48029));
    LocalMux I__9357 (
            .O(N__48126),
            .I(N__48024));
    Span4Mux_v I__9356 (
            .O(N__48117),
            .I(N__48024));
    LocalMux I__9355 (
            .O(N__48108),
            .I(N__48013));
    LocalMux I__9354 (
            .O(N__48099),
            .I(N__48013));
    LocalMux I__9353 (
            .O(N__48094),
            .I(N__48013));
    Span4Mux_h I__9352 (
            .O(N__48091),
            .I(N__48013));
    Span4Mux_v I__9351 (
            .O(N__48088),
            .I(N__48013));
    InMux I__9350 (
            .O(N__48087),
            .I(N__48006));
    InMux I__9349 (
            .O(N__48086),
            .I(N__48006));
    InMux I__9348 (
            .O(N__48085),
            .I(N__48006));
    LocalMux I__9347 (
            .O(N__48078),
            .I(N__48003));
    InMux I__9346 (
            .O(N__48077),
            .I(N__48000));
    LocalMux I__9345 (
            .O(N__48072),
            .I(N__47995));
    LocalMux I__9344 (
            .O(N__48069),
            .I(N__47995));
    InMux I__9343 (
            .O(N__48068),
            .I(N__47991));
    InMux I__9342 (
            .O(N__48067),
            .I(N__47988));
    LocalMux I__9341 (
            .O(N__48064),
            .I(N__47983));
    Span4Mux_v I__9340 (
            .O(N__48047),
            .I(N__47983));
    LocalMux I__9339 (
            .O(N__48036),
            .I(N__47974));
    LocalMux I__9338 (
            .O(N__48029),
            .I(N__47974));
    Span4Mux_h I__9337 (
            .O(N__48024),
            .I(N__47974));
    Span4Mux_v I__9336 (
            .O(N__48013),
            .I(N__47974));
    LocalMux I__9335 (
            .O(N__48006),
            .I(N__47969));
    Span4Mux_h I__9334 (
            .O(N__48003),
            .I(N__47969));
    LocalMux I__9333 (
            .O(N__48000),
            .I(N__47964));
    Span4Mux_v I__9332 (
            .O(N__47995),
            .I(N__47964));
    InMux I__9331 (
            .O(N__47994),
            .I(N__47961));
    LocalMux I__9330 (
            .O(N__47991),
            .I(N__47956));
    LocalMux I__9329 (
            .O(N__47988),
            .I(N__47956));
    Sp12to4 I__9328 (
            .O(N__47983),
            .I(N__47953));
    Span4Mux_v I__9327 (
            .O(N__47974),
            .I(N__47950));
    Span4Mux_h I__9326 (
            .O(N__47969),
            .I(N__47947));
    Sp12to4 I__9325 (
            .O(N__47964),
            .I(N__47944));
    LocalMux I__9324 (
            .O(N__47961),
            .I(N__47939));
    Span12Mux_v I__9323 (
            .O(N__47956),
            .I(N__47939));
    Span12Mux_h I__9322 (
            .O(N__47953),
            .I(N__47936));
    Span4Mux_v I__9321 (
            .O(N__47950),
            .I(N__47933));
    Span4Mux_v I__9320 (
            .O(N__47947),
            .I(N__47930));
    Span12Mux_h I__9319 (
            .O(N__47944),
            .I(N__47927));
    Span12Mux_v I__9318 (
            .O(N__47939),
            .I(N__47922));
    Span12Mux_v I__9317 (
            .O(N__47936),
            .I(N__47922));
    Span4Mux_v I__9316 (
            .O(N__47933),
            .I(N__47919));
    Odrv4 I__9315 (
            .O(N__47930),
            .I(FRAME_MATCHER_state_31_N_2975_2));
    Odrv12 I__9314 (
            .O(N__47927),
            .I(FRAME_MATCHER_state_31_N_2975_2));
    Odrv12 I__9313 (
            .O(N__47922),
            .I(FRAME_MATCHER_state_31_N_2975_2));
    Odrv4 I__9312 (
            .O(N__47919),
            .I(FRAME_MATCHER_state_31_N_2975_2));
    CascadeMux I__9311 (
            .O(N__47910),
            .I(\c0.n22_adj_4643_cascade_ ));
    CascadeMux I__9310 (
            .O(N__47907),
            .I(\c0.n10_adj_4639_cascade_ ));
    InMux I__9309 (
            .O(N__47904),
            .I(N__47901));
    LocalMux I__9308 (
            .O(N__47901),
            .I(\c0.n13_adj_4640 ));
    CascadeMux I__9307 (
            .O(N__47898),
            .I(\c0.n22134_cascade_ ));
    CascadeMux I__9306 (
            .O(N__47895),
            .I(N__47890));
    InMux I__9305 (
            .O(N__47894),
            .I(N__47887));
    InMux I__9304 (
            .O(N__47893),
            .I(N__47884));
    InMux I__9303 (
            .O(N__47890),
            .I(N__47880));
    LocalMux I__9302 (
            .O(N__47887),
            .I(N__47873));
    LocalMux I__9301 (
            .O(N__47884),
            .I(N__47873));
    InMux I__9300 (
            .O(N__47883),
            .I(N__47870));
    LocalMux I__9299 (
            .O(N__47880),
            .I(N__47867));
    InMux I__9298 (
            .O(N__47879),
            .I(N__47862));
    InMux I__9297 (
            .O(N__47878),
            .I(N__47862));
    Span4Mux_h I__9296 (
            .O(N__47873),
            .I(N__47859));
    LocalMux I__9295 (
            .O(N__47870),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv12 I__9294 (
            .O(N__47867),
            .I(\c0.FRAME_MATCHER_state_11 ));
    LocalMux I__9293 (
            .O(N__47862),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv4 I__9292 (
            .O(N__47859),
            .I(\c0.FRAME_MATCHER_state_11 ));
    SRMux I__9291 (
            .O(N__47850),
            .I(N__47847));
    LocalMux I__9290 (
            .O(N__47847),
            .I(N__47844));
    Odrv4 I__9289 (
            .O(N__47844),
            .I(\c0.n21633 ));
    InMux I__9288 (
            .O(N__47841),
            .I(N__47838));
    LocalMux I__9287 (
            .O(N__47838),
            .I(N__47833));
    InMux I__9286 (
            .O(N__47837),
            .I(N__47830));
    InMux I__9285 (
            .O(N__47836),
            .I(N__47824));
    Span4Mux_v I__9284 (
            .O(N__47833),
            .I(N__47819));
    LocalMux I__9283 (
            .O(N__47830),
            .I(N__47819));
    InMux I__9282 (
            .O(N__47829),
            .I(N__47809));
    InMux I__9281 (
            .O(N__47828),
            .I(N__47809));
    InMux I__9280 (
            .O(N__47827),
            .I(N__47806));
    LocalMux I__9279 (
            .O(N__47824),
            .I(N__47803));
    Span4Mux_h I__9278 (
            .O(N__47819),
            .I(N__47800));
    InMux I__9277 (
            .O(N__47818),
            .I(N__47791));
    InMux I__9276 (
            .O(N__47817),
            .I(N__47791));
    InMux I__9275 (
            .O(N__47816),
            .I(N__47791));
    InMux I__9274 (
            .O(N__47815),
            .I(N__47791));
    InMux I__9273 (
            .O(N__47814),
            .I(N__47784));
    LocalMux I__9272 (
            .O(N__47809),
            .I(N__47781));
    LocalMux I__9271 (
            .O(N__47806),
            .I(N__47778));
    Span12Mux_v I__9270 (
            .O(N__47803),
            .I(N__47775));
    Span4Mux_v I__9269 (
            .O(N__47800),
            .I(N__47770));
    LocalMux I__9268 (
            .O(N__47791),
            .I(N__47770));
    InMux I__9267 (
            .O(N__47790),
            .I(N__47763));
    InMux I__9266 (
            .O(N__47789),
            .I(N__47763));
    InMux I__9265 (
            .O(N__47788),
            .I(N__47763));
    InMux I__9264 (
            .O(N__47787),
            .I(N__47760));
    LocalMux I__9263 (
            .O(N__47784),
            .I(N__47757));
    Span4Mux_h I__9262 (
            .O(N__47781),
            .I(N__47752));
    Span4Mux_v I__9261 (
            .O(N__47778),
            .I(N__47752));
    Odrv12 I__9260 (
            .O(N__47775),
            .I(\c0.n6 ));
    Odrv4 I__9259 (
            .O(N__47770),
            .I(\c0.n6 ));
    LocalMux I__9258 (
            .O(N__47763),
            .I(\c0.n6 ));
    LocalMux I__9257 (
            .O(N__47760),
            .I(\c0.n6 ));
    Odrv4 I__9256 (
            .O(N__47757),
            .I(\c0.n6 ));
    Odrv4 I__9255 (
            .O(N__47752),
            .I(\c0.n6 ));
    InMux I__9254 (
            .O(N__47739),
            .I(N__47736));
    LocalMux I__9253 (
            .O(N__47736),
            .I(\c0.n18_adj_4485 ));
    CascadeMux I__9252 (
            .O(N__47733),
            .I(N__47717));
    InMux I__9251 (
            .O(N__47732),
            .I(N__47712));
    InMux I__9250 (
            .O(N__47731),
            .I(N__47700));
    InMux I__9249 (
            .O(N__47730),
            .I(N__47700));
    InMux I__9248 (
            .O(N__47729),
            .I(N__47700));
    InMux I__9247 (
            .O(N__47728),
            .I(N__47700));
    InMux I__9246 (
            .O(N__47727),
            .I(N__47700));
    InMux I__9245 (
            .O(N__47726),
            .I(N__47697));
    InMux I__9244 (
            .O(N__47725),
            .I(N__47691));
    InMux I__9243 (
            .O(N__47724),
            .I(N__47691));
    InMux I__9242 (
            .O(N__47723),
            .I(N__47688));
    InMux I__9241 (
            .O(N__47722),
            .I(N__47683));
    InMux I__9240 (
            .O(N__47721),
            .I(N__47683));
    InMux I__9239 (
            .O(N__47720),
            .I(N__47680));
    InMux I__9238 (
            .O(N__47717),
            .I(N__47673));
    InMux I__9237 (
            .O(N__47716),
            .I(N__47673));
    InMux I__9236 (
            .O(N__47715),
            .I(N__47673));
    LocalMux I__9235 (
            .O(N__47712),
            .I(N__47670));
    InMux I__9234 (
            .O(N__47711),
            .I(N__47667));
    LocalMux I__9233 (
            .O(N__47700),
            .I(N__47662));
    LocalMux I__9232 (
            .O(N__47697),
            .I(N__47662));
    InMux I__9231 (
            .O(N__47696),
            .I(N__47659));
    LocalMux I__9230 (
            .O(N__47691),
            .I(N__47649));
    LocalMux I__9229 (
            .O(N__47688),
            .I(N__47642));
    LocalMux I__9228 (
            .O(N__47683),
            .I(N__47642));
    LocalMux I__9227 (
            .O(N__47680),
            .I(N__47637));
    LocalMux I__9226 (
            .O(N__47673),
            .I(N__47637));
    Span4Mux_v I__9225 (
            .O(N__47670),
            .I(N__47628));
    LocalMux I__9224 (
            .O(N__47667),
            .I(N__47628));
    Span4Mux_v I__9223 (
            .O(N__47662),
            .I(N__47628));
    LocalMux I__9222 (
            .O(N__47659),
            .I(N__47628));
    InMux I__9221 (
            .O(N__47658),
            .I(N__47623));
    InMux I__9220 (
            .O(N__47657),
            .I(N__47623));
    InMux I__9219 (
            .O(N__47656),
            .I(N__47616));
    InMux I__9218 (
            .O(N__47655),
            .I(N__47616));
    InMux I__9217 (
            .O(N__47654),
            .I(N__47616));
    InMux I__9216 (
            .O(N__47653),
            .I(N__47613));
    CascadeMux I__9215 (
            .O(N__47652),
            .I(N__47607));
    Span4Mux_v I__9214 (
            .O(N__47649),
            .I(N__47604));
    InMux I__9213 (
            .O(N__47648),
            .I(N__47599));
    InMux I__9212 (
            .O(N__47647),
            .I(N__47599));
    Span4Mux_v I__9211 (
            .O(N__47642),
            .I(N__47594));
    Span4Mux_h I__9210 (
            .O(N__47637),
            .I(N__47585));
    Span4Mux_v I__9209 (
            .O(N__47628),
            .I(N__47585));
    LocalMux I__9208 (
            .O(N__47623),
            .I(N__47585));
    LocalMux I__9207 (
            .O(N__47616),
            .I(N__47585));
    LocalMux I__9206 (
            .O(N__47613),
            .I(N__47582));
    InMux I__9205 (
            .O(N__47612),
            .I(N__47579));
    InMux I__9204 (
            .O(N__47611),
            .I(N__47576));
    InMux I__9203 (
            .O(N__47610),
            .I(N__47571));
    InMux I__9202 (
            .O(N__47607),
            .I(N__47571));
    Span4Mux_h I__9201 (
            .O(N__47604),
            .I(N__47566));
    LocalMux I__9200 (
            .O(N__47599),
            .I(N__47566));
    InMux I__9199 (
            .O(N__47598),
            .I(N__47563));
    InMux I__9198 (
            .O(N__47597),
            .I(N__47560));
    Sp12to4 I__9197 (
            .O(N__47594),
            .I(N__47557));
    Span4Mux_h I__9196 (
            .O(N__47585),
            .I(N__47554));
    Span12Mux_v I__9195 (
            .O(N__47582),
            .I(N__47545));
    LocalMux I__9194 (
            .O(N__47579),
            .I(N__47545));
    LocalMux I__9193 (
            .O(N__47576),
            .I(N__47545));
    LocalMux I__9192 (
            .O(N__47571),
            .I(N__47545));
    Sp12to4 I__9191 (
            .O(N__47566),
            .I(N__47538));
    LocalMux I__9190 (
            .O(N__47563),
            .I(N__47538));
    LocalMux I__9189 (
            .O(N__47560),
            .I(N__47538));
    Span12Mux_h I__9188 (
            .O(N__47557),
            .I(N__47535));
    Span4Mux_h I__9187 (
            .O(N__47554),
            .I(N__47532));
    Span12Mux_h I__9186 (
            .O(N__47545),
            .I(N__47527));
    Span12Mux_s11_v I__9185 (
            .O(N__47538),
            .I(N__47527));
    Odrv12 I__9184 (
            .O(N__47535),
            .I(count_enable));
    Odrv4 I__9183 (
            .O(N__47532),
            .I(count_enable));
    Odrv12 I__9182 (
            .O(N__47527),
            .I(count_enable));
    InMux I__9181 (
            .O(N__47520),
            .I(N__47517));
    LocalMux I__9180 (
            .O(N__47517),
            .I(N__47514));
    Span4Mux_h I__9179 (
            .O(N__47514),
            .I(N__47511));
    Span4Mux_v I__9178 (
            .O(N__47511),
            .I(N__47508));
    Span4Mux_v I__9177 (
            .O(N__47508),
            .I(N__47505));
    Odrv4 I__9176 (
            .O(N__47505),
            .I(n2343));
    CascadeMux I__9175 (
            .O(N__47502),
            .I(N__47498));
    CascadeMux I__9174 (
            .O(N__47501),
            .I(N__47494));
    InMux I__9173 (
            .O(N__47498),
            .I(N__47489));
    InMux I__9172 (
            .O(N__47497),
            .I(N__47489));
    InMux I__9171 (
            .O(N__47494),
            .I(N__47486));
    LocalMux I__9170 (
            .O(N__47489),
            .I(N__47481));
    LocalMux I__9169 (
            .O(N__47486),
            .I(N__47478));
    InMux I__9168 (
            .O(N__47485),
            .I(N__47475));
    InMux I__9167 (
            .O(N__47484),
            .I(N__47472));
    Span4Mux_h I__9166 (
            .O(N__47481),
            .I(N__47469));
    Sp12to4 I__9165 (
            .O(N__47478),
            .I(N__47465));
    LocalMux I__9164 (
            .O(N__47475),
            .I(N__47462));
    LocalMux I__9163 (
            .O(N__47472),
            .I(N__47457));
    Span4Mux_v I__9162 (
            .O(N__47469),
            .I(N__47457));
    InMux I__9161 (
            .O(N__47468),
            .I(N__47453));
    Span12Mux_v I__9160 (
            .O(N__47465),
            .I(N__47450));
    Span12Mux_h I__9159 (
            .O(N__47462),
            .I(N__47447));
    Span4Mux_v I__9158 (
            .O(N__47457),
            .I(N__47444));
    InMux I__9157 (
            .O(N__47456),
            .I(N__47441));
    LocalMux I__9156 (
            .O(N__47453),
            .I(encoder0_position_14));
    Odrv12 I__9155 (
            .O(N__47450),
            .I(encoder0_position_14));
    Odrv12 I__9154 (
            .O(N__47447),
            .I(encoder0_position_14));
    Odrv4 I__9153 (
            .O(N__47444),
            .I(encoder0_position_14));
    LocalMux I__9152 (
            .O(N__47441),
            .I(encoder0_position_14));
    InMux I__9151 (
            .O(N__47430),
            .I(N__47426));
    InMux I__9150 (
            .O(N__47429),
            .I(N__47423));
    LocalMux I__9149 (
            .O(N__47426),
            .I(N__47420));
    LocalMux I__9148 (
            .O(N__47423),
            .I(N__47415));
    Span4Mux_v I__9147 (
            .O(N__47420),
            .I(N__47415));
    Span4Mux_h I__9146 (
            .O(N__47415),
            .I(N__47412));
    Odrv4 I__9145 (
            .O(N__47412),
            .I(n4_adj_4761));
    CascadeMux I__9144 (
            .O(N__47409),
            .I(N__47405));
    CascadeMux I__9143 (
            .O(N__47408),
            .I(N__47402));
    InMux I__9142 (
            .O(N__47405),
            .I(N__47399));
    InMux I__9141 (
            .O(N__47402),
            .I(N__47396));
    LocalMux I__9140 (
            .O(N__47399),
            .I(N__47393));
    LocalMux I__9139 (
            .O(N__47396),
            .I(\c0.data_in_frame_29_3 ));
    Odrv4 I__9138 (
            .O(N__47393),
            .I(\c0.data_in_frame_29_3 ));
    InMux I__9137 (
            .O(N__47388),
            .I(N__47385));
    LocalMux I__9136 (
            .O(N__47385),
            .I(N__47382));
    Span4Mux_v I__9135 (
            .O(N__47382),
            .I(N__47379));
    Odrv4 I__9134 (
            .O(N__47379),
            .I(\c0.n17_adj_4483 ));
    CascadeMux I__9133 (
            .O(N__47376),
            .I(\c0.n26_adj_4480_cascade_ ));
    InMux I__9132 (
            .O(N__47373),
            .I(N__47370));
    LocalMux I__9131 (
            .O(N__47370),
            .I(N__47367));
    Span4Mux_h I__9130 (
            .O(N__47367),
            .I(N__47363));
    InMux I__9129 (
            .O(N__47366),
            .I(N__47360));
    Odrv4 I__9128 (
            .O(N__47363),
            .I(\c0.n63_adj_4249 ));
    LocalMux I__9127 (
            .O(N__47360),
            .I(\c0.n63_adj_4249 ));
    CascadeMux I__9126 (
            .O(N__47355),
            .I(\c0.n34_adj_4546_cascade_ ));
    CascadeMux I__9125 (
            .O(N__47352),
            .I(N__47344));
    InMux I__9124 (
            .O(N__47351),
            .I(N__47336));
    InMux I__9123 (
            .O(N__47350),
            .I(N__47336));
    InMux I__9122 (
            .O(N__47349),
            .I(N__47336));
    InMux I__9121 (
            .O(N__47348),
            .I(N__47333));
    InMux I__9120 (
            .O(N__47347),
            .I(N__47326));
    InMux I__9119 (
            .O(N__47344),
            .I(N__47326));
    InMux I__9118 (
            .O(N__47343),
            .I(N__47326));
    LocalMux I__9117 (
            .O(N__47336),
            .I(n24622));
    LocalMux I__9116 (
            .O(N__47333),
            .I(n24622));
    LocalMux I__9115 (
            .O(N__47326),
            .I(n24622));
    CascadeMux I__9114 (
            .O(N__47319),
            .I(n24622_cascade_));
    CascadeMux I__9113 (
            .O(N__47316),
            .I(N__47313));
    InMux I__9112 (
            .O(N__47313),
            .I(N__47309));
    InMux I__9111 (
            .O(N__47312),
            .I(N__47306));
    LocalMux I__9110 (
            .O(N__47309),
            .I(N__47302));
    LocalMux I__9109 (
            .O(N__47306),
            .I(N__47299));
    CascadeMux I__9108 (
            .O(N__47305),
            .I(N__47295));
    Span4Mux_h I__9107 (
            .O(N__47302),
            .I(N__47290));
    Span4Mux_h I__9106 (
            .O(N__47299),
            .I(N__47287));
    InMux I__9105 (
            .O(N__47298),
            .I(N__47278));
    InMux I__9104 (
            .O(N__47295),
            .I(N__47278));
    InMux I__9103 (
            .O(N__47294),
            .I(N__47278));
    InMux I__9102 (
            .O(N__47293),
            .I(N__47278));
    Span4Mux_h I__9101 (
            .O(N__47290),
            .I(N__47271));
    Span4Mux_v I__9100 (
            .O(N__47287),
            .I(N__47271));
    LocalMux I__9099 (
            .O(N__47278),
            .I(N__47268));
    InMux I__9098 (
            .O(N__47277),
            .I(N__47265));
    InMux I__9097 (
            .O(N__47276),
            .I(N__47262));
    Span4Mux_v I__9096 (
            .O(N__47271),
            .I(N__47259));
    Span12Mux_s11_v I__9095 (
            .O(N__47268),
            .I(N__47256));
    LocalMux I__9094 (
            .O(N__47265),
            .I(control_mode_2));
    LocalMux I__9093 (
            .O(N__47262),
            .I(control_mode_2));
    Odrv4 I__9092 (
            .O(N__47259),
            .I(control_mode_2));
    Odrv12 I__9091 (
            .O(N__47256),
            .I(control_mode_2));
    InMux I__9090 (
            .O(N__47247),
            .I(N__47244));
    LocalMux I__9089 (
            .O(N__47244),
            .I(\c0.n24539 ));
    InMux I__9088 (
            .O(N__47241),
            .I(N__47238));
    LocalMux I__9087 (
            .O(N__47238),
            .I(\c0.n24733 ));
    InMux I__9086 (
            .O(N__47235),
            .I(N__47228));
    InMux I__9085 (
            .O(N__47234),
            .I(N__47224));
    InMux I__9084 (
            .O(N__47233),
            .I(N__47221));
    CascadeMux I__9083 (
            .O(N__47232),
            .I(N__47218));
    InMux I__9082 (
            .O(N__47231),
            .I(N__47215));
    LocalMux I__9081 (
            .O(N__47228),
            .I(N__47212));
    InMux I__9080 (
            .O(N__47227),
            .I(N__47209));
    LocalMux I__9079 (
            .O(N__47224),
            .I(N__47206));
    LocalMux I__9078 (
            .O(N__47221),
            .I(N__47203));
    InMux I__9077 (
            .O(N__47218),
            .I(N__47200));
    LocalMux I__9076 (
            .O(N__47215),
            .I(N__47197));
    Span4Mux_v I__9075 (
            .O(N__47212),
            .I(N__47194));
    LocalMux I__9074 (
            .O(N__47209),
            .I(N__47191));
    Span4Mux_v I__9073 (
            .O(N__47206),
            .I(N__47188));
    Span4Mux_v I__9072 (
            .O(N__47203),
            .I(N__47183));
    LocalMux I__9071 (
            .O(N__47200),
            .I(N__47183));
    Span4Mux_v I__9070 (
            .O(N__47197),
            .I(N__47180));
    Span4Mux_v I__9069 (
            .O(N__47194),
            .I(N__47174));
    Span4Mux_v I__9068 (
            .O(N__47191),
            .I(N__47174));
    Span4Mux_h I__9067 (
            .O(N__47188),
            .I(N__47167));
    Span4Mux_v I__9066 (
            .O(N__47183),
            .I(N__47167));
    Span4Mux_h I__9065 (
            .O(N__47180),
            .I(N__47167));
    InMux I__9064 (
            .O(N__47179),
            .I(N__47164));
    Sp12to4 I__9063 (
            .O(N__47174),
            .I(N__47159));
    Sp12to4 I__9062 (
            .O(N__47167),
            .I(N__47159));
    LocalMux I__9061 (
            .O(N__47164),
            .I(r_Bit_Index_0));
    Odrv12 I__9060 (
            .O(N__47159),
            .I(r_Bit_Index_0));
    CascadeMux I__9059 (
            .O(N__47154),
            .I(\c0.rx.n17834_cascade_ ));
    InMux I__9058 (
            .O(N__47151),
            .I(N__47146));
    InMux I__9057 (
            .O(N__47150),
            .I(N__47143));
    InMux I__9056 (
            .O(N__47149),
            .I(N__47139));
    LocalMux I__9055 (
            .O(N__47146),
            .I(N__47136));
    LocalMux I__9054 (
            .O(N__47143),
            .I(N__47133));
    InMux I__9053 (
            .O(N__47142),
            .I(N__47130));
    LocalMux I__9052 (
            .O(N__47139),
            .I(N__47127));
    Span4Mux_h I__9051 (
            .O(N__47136),
            .I(N__47124));
    Span4Mux_h I__9050 (
            .O(N__47133),
            .I(N__47121));
    LocalMux I__9049 (
            .O(N__47130),
            .I(N__47118));
    Span4Mux_v I__9048 (
            .O(N__47127),
            .I(N__47115));
    Span4Mux_h I__9047 (
            .O(N__47124),
            .I(N__47112));
    Odrv4 I__9046 (
            .O(N__47121),
            .I(n14484));
    Odrv4 I__9045 (
            .O(N__47118),
            .I(n14484));
    Odrv4 I__9044 (
            .O(N__47115),
            .I(n14484));
    Odrv4 I__9043 (
            .O(N__47112),
            .I(n14484));
    InMux I__9042 (
            .O(N__47103),
            .I(N__47099));
    InMux I__9041 (
            .O(N__47102),
            .I(N__47095));
    LocalMux I__9040 (
            .O(N__47099),
            .I(N__47092));
    InMux I__9039 (
            .O(N__47098),
            .I(N__47089));
    LocalMux I__9038 (
            .O(N__47095),
            .I(N__47086));
    Span4Mux_v I__9037 (
            .O(N__47092),
            .I(N__47083));
    LocalMux I__9036 (
            .O(N__47089),
            .I(N__47080));
    Span4Mux_h I__9035 (
            .O(N__47086),
            .I(N__47077));
    Span4Mux_h I__9034 (
            .O(N__47083),
            .I(N__47072));
    Span4Mux_v I__9033 (
            .O(N__47080),
            .I(N__47072));
    Span4Mux_v I__9032 (
            .O(N__47077),
            .I(N__47067));
    Span4Mux_h I__9031 (
            .O(N__47072),
            .I(N__47067));
    Odrv4 I__9030 (
            .O(N__47067),
            .I(n14988));
    InMux I__9029 (
            .O(N__47064),
            .I(N__47061));
    LocalMux I__9028 (
            .O(N__47061),
            .I(N__47058));
    Span4Mux_h I__9027 (
            .O(N__47058),
            .I(N__47054));
    InMux I__9026 (
            .O(N__47057),
            .I(N__47048));
    Span4Mux_h I__9025 (
            .O(N__47054),
            .I(N__47045));
    InMux I__9024 (
            .O(N__47053),
            .I(N__47040));
    InMux I__9023 (
            .O(N__47052),
            .I(N__47040));
    InMux I__9022 (
            .O(N__47051),
            .I(N__47037));
    LocalMux I__9021 (
            .O(N__47048),
            .I(control_mode_5));
    Odrv4 I__9020 (
            .O(N__47045),
            .I(control_mode_5));
    LocalMux I__9019 (
            .O(N__47040),
            .I(control_mode_5));
    LocalMux I__9018 (
            .O(N__47037),
            .I(control_mode_5));
    InMux I__9017 (
            .O(N__47028),
            .I(N__47024));
    CascadeMux I__9016 (
            .O(N__47027),
            .I(N__47021));
    LocalMux I__9015 (
            .O(N__47024),
            .I(N__47018));
    InMux I__9014 (
            .O(N__47021),
            .I(N__47015));
    Span4Mux_h I__9013 (
            .O(N__47018),
            .I(N__47008));
    LocalMux I__9012 (
            .O(N__47015),
            .I(N__47004));
    InMux I__9011 (
            .O(N__47014),
            .I(N__47001));
    InMux I__9010 (
            .O(N__47013),
            .I(N__46994));
    InMux I__9009 (
            .O(N__47012),
            .I(N__46994));
    InMux I__9008 (
            .O(N__47011),
            .I(N__46994));
    Span4Mux_v I__9007 (
            .O(N__47008),
            .I(N__46991));
    InMux I__9006 (
            .O(N__47007),
            .I(N__46988));
    Span4Mux_h I__9005 (
            .O(N__47004),
            .I(N__46985));
    LocalMux I__9004 (
            .O(N__47001),
            .I(N__46982));
    LocalMux I__9003 (
            .O(N__46994),
            .I(N__46979));
    Span4Mux_v I__9002 (
            .O(N__46991),
            .I(N__46976));
    LocalMux I__9001 (
            .O(N__46988),
            .I(N__46969));
    Span4Mux_h I__9000 (
            .O(N__46985),
            .I(N__46969));
    Span4Mux_v I__8999 (
            .O(N__46982),
            .I(N__46969));
    Odrv12 I__8998 (
            .O(N__46979),
            .I(control_mode_1));
    Odrv4 I__8997 (
            .O(N__46976),
            .I(control_mode_1));
    Odrv4 I__8996 (
            .O(N__46969),
            .I(control_mode_1));
    CascadeMux I__8995 (
            .O(N__46962),
            .I(N__46959));
    InMux I__8994 (
            .O(N__46959),
            .I(N__46956));
    LocalMux I__8993 (
            .O(N__46956),
            .I(N__46950));
    InMux I__8992 (
            .O(N__46955),
            .I(N__46946));
    InMux I__8991 (
            .O(N__46954),
            .I(N__46943));
    InMux I__8990 (
            .O(N__46953),
            .I(N__46940));
    Span12Mux_h I__8989 (
            .O(N__46950),
            .I(N__46937));
    InMux I__8988 (
            .O(N__46949),
            .I(N__46934));
    LocalMux I__8987 (
            .O(N__46946),
            .I(N__46929));
    LocalMux I__8986 (
            .O(N__46943),
            .I(N__46929));
    LocalMux I__8985 (
            .O(N__46940),
            .I(control_mode_3));
    Odrv12 I__8984 (
            .O(N__46937),
            .I(control_mode_3));
    LocalMux I__8983 (
            .O(N__46934),
            .I(control_mode_3));
    Odrv12 I__8982 (
            .O(N__46929),
            .I(control_mode_3));
    InMux I__8981 (
            .O(N__46920),
            .I(N__46915));
    InMux I__8980 (
            .O(N__46919),
            .I(N__46910));
    InMux I__8979 (
            .O(N__46918),
            .I(N__46910));
    LocalMux I__8978 (
            .O(N__46915),
            .I(N__46907));
    LocalMux I__8977 (
            .O(N__46910),
            .I(N__46903));
    Span4Mux_h I__8976 (
            .O(N__46907),
            .I(N__46900));
    InMux I__8975 (
            .O(N__46906),
            .I(N__46897));
    Span4Mux_h I__8974 (
            .O(N__46903),
            .I(N__46894));
    Odrv4 I__8973 (
            .O(N__46900),
            .I(data_in_2_3));
    LocalMux I__8972 (
            .O(N__46897),
            .I(data_in_2_3));
    Odrv4 I__8971 (
            .O(N__46894),
            .I(data_in_2_3));
    CascadeMux I__8970 (
            .O(N__46887),
            .I(\c0.n82_cascade_ ));
    InMux I__8969 (
            .O(N__46884),
            .I(N__46880));
    InMux I__8968 (
            .O(N__46883),
            .I(N__46874));
    LocalMux I__8967 (
            .O(N__46880),
            .I(N__46870));
    InMux I__8966 (
            .O(N__46879),
            .I(N__46867));
    InMux I__8965 (
            .O(N__46878),
            .I(N__46864));
    InMux I__8964 (
            .O(N__46877),
            .I(N__46861));
    LocalMux I__8963 (
            .O(N__46874),
            .I(N__46858));
    CascadeMux I__8962 (
            .O(N__46873),
            .I(N__46855));
    Span4Mux_v I__8961 (
            .O(N__46870),
            .I(N__46851));
    LocalMux I__8960 (
            .O(N__46867),
            .I(N__46846));
    LocalMux I__8959 (
            .O(N__46864),
            .I(N__46846));
    LocalMux I__8958 (
            .O(N__46861),
            .I(N__46841));
    Span4Mux_v I__8957 (
            .O(N__46858),
            .I(N__46841));
    InMux I__8956 (
            .O(N__46855),
            .I(N__46836));
    InMux I__8955 (
            .O(N__46854),
            .I(N__46836));
    Odrv4 I__8954 (
            .O(N__46851),
            .I(\c0.n10467 ));
    Odrv4 I__8953 (
            .O(N__46846),
            .I(\c0.n10467 ));
    Odrv4 I__8952 (
            .O(N__46841),
            .I(\c0.n10467 ));
    LocalMux I__8951 (
            .O(N__46836),
            .I(\c0.n10467 ));
    CascadeMux I__8950 (
            .O(N__46827),
            .I(N__46819));
    CascadeMux I__8949 (
            .O(N__46826),
            .I(N__46816));
    InMux I__8948 (
            .O(N__46825),
            .I(N__46808));
    InMux I__8947 (
            .O(N__46824),
            .I(N__46808));
    InMux I__8946 (
            .O(N__46823),
            .I(N__46808));
    InMux I__8945 (
            .O(N__46822),
            .I(N__46801));
    InMux I__8944 (
            .O(N__46819),
            .I(N__46801));
    InMux I__8943 (
            .O(N__46816),
            .I(N__46801));
    InMux I__8942 (
            .O(N__46815),
            .I(N__46797));
    LocalMux I__8941 (
            .O(N__46808),
            .I(N__46792));
    LocalMux I__8940 (
            .O(N__46801),
            .I(N__46792));
    InMux I__8939 (
            .O(N__46800),
            .I(N__46786));
    LocalMux I__8938 (
            .O(N__46797),
            .I(N__46783));
    Span4Mux_v I__8937 (
            .O(N__46792),
            .I(N__46780));
    InMux I__8936 (
            .O(N__46791),
            .I(N__46773));
    InMux I__8935 (
            .O(N__46790),
            .I(N__46773));
    InMux I__8934 (
            .O(N__46789),
            .I(N__46773));
    LocalMux I__8933 (
            .O(N__46786),
            .I(N__46770));
    Span4Mux_h I__8932 (
            .O(N__46783),
            .I(N__46767));
    Span4Mux_h I__8931 (
            .O(N__46780),
            .I(N__46762));
    LocalMux I__8930 (
            .O(N__46773),
            .I(N__46762));
    Span4Mux_v I__8929 (
            .O(N__46770),
            .I(N__46759));
    Odrv4 I__8928 (
            .O(N__46767),
            .I(\c0.n10500 ));
    Odrv4 I__8927 (
            .O(N__46762),
            .I(\c0.n10500 ));
    Odrv4 I__8926 (
            .O(N__46759),
            .I(\c0.n10500 ));
    InMux I__8925 (
            .O(N__46752),
            .I(N__46749));
    LocalMux I__8924 (
            .O(N__46749),
            .I(N__46746));
    Span4Mux_h I__8923 (
            .O(N__46746),
            .I(N__46737));
    InMux I__8922 (
            .O(N__46745),
            .I(N__46732));
    InMux I__8921 (
            .O(N__46744),
            .I(N__46732));
    InMux I__8920 (
            .O(N__46743),
            .I(N__46723));
    InMux I__8919 (
            .O(N__46742),
            .I(N__46723));
    InMux I__8918 (
            .O(N__46741),
            .I(N__46723));
    InMux I__8917 (
            .O(N__46740),
            .I(N__46723));
    Odrv4 I__8916 (
            .O(N__46737),
            .I(\c0.n21349 ));
    LocalMux I__8915 (
            .O(N__46732),
            .I(\c0.n21349 ));
    LocalMux I__8914 (
            .O(N__46723),
            .I(\c0.n21349 ));
    InMux I__8913 (
            .O(N__46716),
            .I(N__46713));
    LocalMux I__8912 (
            .O(N__46713),
            .I(\c0.n4_adj_4271 ));
    InMux I__8911 (
            .O(N__46710),
            .I(N__46707));
    LocalMux I__8910 (
            .O(N__46707),
            .I(\c0.data_out_frame_29__6__N_1538 ));
    InMux I__8909 (
            .O(N__46704),
            .I(N__46700));
    InMux I__8908 (
            .O(N__46703),
            .I(N__46697));
    LocalMux I__8907 (
            .O(N__46700),
            .I(N__46691));
    LocalMux I__8906 (
            .O(N__46697),
            .I(N__46691));
    InMux I__8905 (
            .O(N__46696),
            .I(N__46688));
    Span4Mux_v I__8904 (
            .O(N__46691),
            .I(N__46683));
    LocalMux I__8903 (
            .O(N__46688),
            .I(N__46683));
    Odrv4 I__8902 (
            .O(N__46683),
            .I(\c0.n21327 ));
    CascadeMux I__8901 (
            .O(N__46680),
            .I(\c0.n4_adj_4271_cascade_ ));
    InMux I__8900 (
            .O(N__46677),
            .I(N__46674));
    LocalMux I__8899 (
            .O(N__46674),
            .I(\c0.data_out_frame_29__3__N_1730 ));
    InMux I__8898 (
            .O(N__46671),
            .I(N__46667));
    InMux I__8897 (
            .O(N__46670),
            .I(N__46664));
    LocalMux I__8896 (
            .O(N__46667),
            .I(N__46661));
    LocalMux I__8895 (
            .O(N__46664),
            .I(data_out_frame_29__3__N_1661));
    Odrv4 I__8894 (
            .O(N__46661),
            .I(data_out_frame_29__3__N_1661));
    InMux I__8893 (
            .O(N__46656),
            .I(N__46653));
    LocalMux I__8892 (
            .O(N__46653),
            .I(N__46649));
    InMux I__8891 (
            .O(N__46652),
            .I(N__46646));
    Span4Mux_v I__8890 (
            .O(N__46649),
            .I(N__46643));
    LocalMux I__8889 (
            .O(N__46646),
            .I(N__46640));
    Odrv4 I__8888 (
            .O(N__46643),
            .I(\c0.rx.n12909 ));
    Odrv4 I__8887 (
            .O(N__46640),
            .I(\c0.rx.n12909 ));
    CascadeMux I__8886 (
            .O(N__46635),
            .I(\c0.n22112_cascade_ ));
    InMux I__8885 (
            .O(N__46632),
            .I(N__46628));
    InMux I__8884 (
            .O(N__46631),
            .I(N__46625));
    LocalMux I__8883 (
            .O(N__46628),
            .I(N__46620));
    LocalMux I__8882 (
            .O(N__46625),
            .I(N__46620));
    Span4Mux_v I__8881 (
            .O(N__46620),
            .I(N__46617));
    Odrv4 I__8880 (
            .O(N__46617),
            .I(\c0.n21355 ));
    InMux I__8879 (
            .O(N__46614),
            .I(N__46611));
    LocalMux I__8878 (
            .O(N__46611),
            .I(N__46603));
    InMux I__8877 (
            .O(N__46610),
            .I(N__46600));
    InMux I__8876 (
            .O(N__46609),
            .I(N__46594));
    InMux I__8875 (
            .O(N__46608),
            .I(N__46594));
    InMux I__8874 (
            .O(N__46607),
            .I(N__46591));
    InMux I__8873 (
            .O(N__46606),
            .I(N__46587));
    Sp12to4 I__8872 (
            .O(N__46603),
            .I(N__46582));
    LocalMux I__8871 (
            .O(N__46600),
            .I(N__46582));
    InMux I__8870 (
            .O(N__46599),
            .I(N__46579));
    LocalMux I__8869 (
            .O(N__46594),
            .I(N__46576));
    LocalMux I__8868 (
            .O(N__46591),
            .I(N__46573));
    InMux I__8867 (
            .O(N__46590),
            .I(N__46570));
    LocalMux I__8866 (
            .O(N__46587),
            .I(\c0.n12604 ));
    Odrv12 I__8865 (
            .O(N__46582),
            .I(\c0.n12604 ));
    LocalMux I__8864 (
            .O(N__46579),
            .I(\c0.n12604 ));
    Odrv4 I__8863 (
            .O(N__46576),
            .I(\c0.n12604 ));
    Odrv4 I__8862 (
            .O(N__46573),
            .I(\c0.n12604 ));
    LocalMux I__8861 (
            .O(N__46570),
            .I(\c0.n12604 ));
    InMux I__8860 (
            .O(N__46557),
            .I(N__46554));
    LocalMux I__8859 (
            .O(N__46554),
            .I(N__46550));
    InMux I__8858 (
            .O(N__46553),
            .I(N__46547));
    Odrv12 I__8857 (
            .O(N__46550),
            .I(\c0.n20786 ));
    LocalMux I__8856 (
            .O(N__46547),
            .I(\c0.n20786 ));
    CascadeMux I__8855 (
            .O(N__46542),
            .I(\c0.n20786_cascade_ ));
    InMux I__8854 (
            .O(N__46539),
            .I(N__46536));
    LocalMux I__8853 (
            .O(N__46536),
            .I(\c0.n9_adj_4494 ));
    InMux I__8852 (
            .O(N__46533),
            .I(N__46529));
    InMux I__8851 (
            .O(N__46532),
            .I(N__46526));
    LocalMux I__8850 (
            .O(N__46529),
            .I(N__46523));
    LocalMux I__8849 (
            .O(N__46526),
            .I(N__46519));
    Span4Mux_h I__8848 (
            .O(N__46523),
            .I(N__46516));
    InMux I__8847 (
            .O(N__46522),
            .I(N__46513));
    Span4Mux_h I__8846 (
            .O(N__46519),
            .I(N__46510));
    Span4Mux_h I__8845 (
            .O(N__46516),
            .I(N__46505));
    LocalMux I__8844 (
            .O(N__46513),
            .I(N__46505));
    Odrv4 I__8843 (
            .O(N__46510),
            .I(\c0.n10497 ));
    Odrv4 I__8842 (
            .O(N__46505),
            .I(\c0.n10497 ));
    InMux I__8841 (
            .O(N__46500),
            .I(N__46493));
    InMux I__8840 (
            .O(N__46499),
            .I(N__46493));
    InMux I__8839 (
            .O(N__46498),
            .I(N__46490));
    LocalMux I__8838 (
            .O(N__46493),
            .I(\c0.n21433 ));
    LocalMux I__8837 (
            .O(N__46490),
            .I(\c0.n21433 ));
    CascadeMux I__8836 (
            .O(N__46485),
            .I(N__46479));
    InMux I__8835 (
            .O(N__46484),
            .I(N__46475));
    InMux I__8834 (
            .O(N__46483),
            .I(N__46466));
    InMux I__8833 (
            .O(N__46482),
            .I(N__46466));
    InMux I__8832 (
            .O(N__46479),
            .I(N__46466));
    InMux I__8831 (
            .O(N__46478),
            .I(N__46466));
    LocalMux I__8830 (
            .O(N__46475),
            .I(\c0.n21311 ));
    LocalMux I__8829 (
            .O(N__46466),
            .I(\c0.n21311 ));
    InMux I__8828 (
            .O(N__46461),
            .I(N__46457));
    InMux I__8827 (
            .O(N__46460),
            .I(N__46454));
    LocalMux I__8826 (
            .O(N__46457),
            .I(\c0.n12590 ));
    LocalMux I__8825 (
            .O(N__46454),
            .I(\c0.n12590 ));
    InMux I__8824 (
            .O(N__46449),
            .I(N__46445));
    CascadeMux I__8823 (
            .O(N__46448),
            .I(N__46441));
    LocalMux I__8822 (
            .O(N__46445),
            .I(N__46437));
    InMux I__8821 (
            .O(N__46444),
            .I(N__46434));
    InMux I__8820 (
            .O(N__46441),
            .I(N__46431));
    InMux I__8819 (
            .O(N__46440),
            .I(N__46428));
    Span4Mux_h I__8818 (
            .O(N__46437),
            .I(N__46425));
    LocalMux I__8817 (
            .O(N__46434),
            .I(N__46422));
    LocalMux I__8816 (
            .O(N__46431),
            .I(N__46417));
    LocalMux I__8815 (
            .O(N__46428),
            .I(N__46417));
    Span4Mux_h I__8814 (
            .O(N__46425),
            .I(N__46414));
    Span4Mux_v I__8813 (
            .O(N__46422),
            .I(N__46411));
    Span4Mux_v I__8812 (
            .O(N__46417),
            .I(N__46408));
    Span4Mux_v I__8811 (
            .O(N__46414),
            .I(N__46405));
    Span4Mux_h I__8810 (
            .O(N__46411),
            .I(N__46402));
    Odrv4 I__8809 (
            .O(N__46408),
            .I(\c0.n21399 ));
    Odrv4 I__8808 (
            .O(N__46405),
            .I(\c0.n21399 ));
    Odrv4 I__8807 (
            .O(N__46402),
            .I(\c0.n21399 ));
    CascadeMux I__8806 (
            .O(N__46395),
            .I(N__46392));
    InMux I__8805 (
            .O(N__46392),
            .I(N__46388));
    InMux I__8804 (
            .O(N__46391),
            .I(N__46385));
    LocalMux I__8803 (
            .O(N__46388),
            .I(N__46382));
    LocalMux I__8802 (
            .O(N__46385),
            .I(N__46379));
    Span4Mux_v I__8801 (
            .O(N__46382),
            .I(N__46373));
    Span4Mux_v I__8800 (
            .O(N__46379),
            .I(N__46373));
    InMux I__8799 (
            .O(N__46378),
            .I(N__46370));
    Span4Mux_h I__8798 (
            .O(N__46373),
            .I(N__46365));
    LocalMux I__8797 (
            .O(N__46370),
            .I(N__46365));
    Odrv4 I__8796 (
            .O(N__46365),
            .I(\c0.n22553 ));
    CascadeMux I__8795 (
            .O(N__46362),
            .I(N__46358));
    CascadeMux I__8794 (
            .O(N__46361),
            .I(N__46353));
    InMux I__8793 (
            .O(N__46358),
            .I(N__46350));
    InMux I__8792 (
            .O(N__46357),
            .I(N__46345));
    InMux I__8791 (
            .O(N__46356),
            .I(N__46342));
    InMux I__8790 (
            .O(N__46353),
            .I(N__46339));
    LocalMux I__8789 (
            .O(N__46350),
            .I(N__46336));
    InMux I__8788 (
            .O(N__46349),
            .I(N__46333));
    InMux I__8787 (
            .O(N__46348),
            .I(N__46330));
    LocalMux I__8786 (
            .O(N__46345),
            .I(N__46326));
    LocalMux I__8785 (
            .O(N__46342),
            .I(N__46323));
    LocalMux I__8784 (
            .O(N__46339),
            .I(N__46320));
    Span4Mux_v I__8783 (
            .O(N__46336),
            .I(N__46315));
    LocalMux I__8782 (
            .O(N__46333),
            .I(N__46315));
    LocalMux I__8781 (
            .O(N__46330),
            .I(N__46311));
    InMux I__8780 (
            .O(N__46329),
            .I(N__46308));
    Span4Mux_v I__8779 (
            .O(N__46326),
            .I(N__46305));
    Span4Mux_h I__8778 (
            .O(N__46323),
            .I(N__46302));
    Span4Mux_v I__8777 (
            .O(N__46320),
            .I(N__46297));
    Span4Mux_h I__8776 (
            .O(N__46315),
            .I(N__46297));
    InMux I__8775 (
            .O(N__46314),
            .I(N__46294));
    Span4Mux_v I__8774 (
            .O(N__46311),
            .I(N__46289));
    LocalMux I__8773 (
            .O(N__46308),
            .I(N__46289));
    Span4Mux_v I__8772 (
            .O(N__46305),
            .I(N__46286));
    Span4Mux_v I__8771 (
            .O(N__46302),
            .I(N__46281));
    Span4Mux_h I__8770 (
            .O(N__46297),
            .I(N__46281));
    LocalMux I__8769 (
            .O(N__46294),
            .I(encoder1_position_2));
    Odrv4 I__8768 (
            .O(N__46289),
            .I(encoder1_position_2));
    Odrv4 I__8767 (
            .O(N__46286),
            .I(encoder1_position_2));
    Odrv4 I__8766 (
            .O(N__46281),
            .I(encoder1_position_2));
    InMux I__8765 (
            .O(N__46272),
            .I(N__46265));
    InMux I__8764 (
            .O(N__46271),
            .I(N__46265));
    InMux I__8763 (
            .O(N__46270),
            .I(N__46261));
    LocalMux I__8762 (
            .O(N__46265),
            .I(N__46258));
    CascadeMux I__8761 (
            .O(N__46264),
            .I(N__46255));
    LocalMux I__8760 (
            .O(N__46261),
            .I(N__46251));
    Span4Mux_h I__8759 (
            .O(N__46258),
            .I(N__46248));
    InMux I__8758 (
            .O(N__46255),
            .I(N__46244));
    InMux I__8757 (
            .O(N__46254),
            .I(N__46241));
    Span4Mux_h I__8756 (
            .O(N__46251),
            .I(N__46236));
    Span4Mux_h I__8755 (
            .O(N__46248),
            .I(N__46236));
    InMux I__8754 (
            .O(N__46247),
            .I(N__46233));
    LocalMux I__8753 (
            .O(N__46244),
            .I(N__46228));
    LocalMux I__8752 (
            .O(N__46241),
            .I(N__46228));
    Odrv4 I__8751 (
            .O(N__46236),
            .I(\c0.n21416 ));
    LocalMux I__8750 (
            .O(N__46233),
            .I(\c0.n21416 ));
    Odrv4 I__8749 (
            .O(N__46228),
            .I(\c0.n21416 ));
    InMux I__8748 (
            .O(N__46221),
            .I(N__46217));
    InMux I__8747 (
            .O(N__46220),
            .I(N__46214));
    LocalMux I__8746 (
            .O(N__46217),
            .I(N__46210));
    LocalMux I__8745 (
            .O(N__46214),
            .I(N__46207));
    InMux I__8744 (
            .O(N__46213),
            .I(N__46204));
    Span4Mux_h I__8743 (
            .O(N__46210),
            .I(N__46199));
    Span4Mux_v I__8742 (
            .O(N__46207),
            .I(N__46199));
    LocalMux I__8741 (
            .O(N__46204),
            .I(N__46196));
    Sp12to4 I__8740 (
            .O(N__46199),
            .I(N__46191));
    Span12Mux_s11_h I__8739 (
            .O(N__46196),
            .I(N__46191));
    Odrv12 I__8738 (
            .O(N__46191),
            .I(\c0.n10531 ));
    InMux I__8737 (
            .O(N__46188),
            .I(N__46185));
    LocalMux I__8736 (
            .O(N__46185),
            .I(N__46180));
    InMux I__8735 (
            .O(N__46184),
            .I(N__46174));
    InMux I__8734 (
            .O(N__46183),
            .I(N__46174));
    Span4Mux_h I__8733 (
            .O(N__46180),
            .I(N__46171));
    InMux I__8732 (
            .O(N__46179),
            .I(N__46168));
    LocalMux I__8731 (
            .O(N__46174),
            .I(N__46165));
    Odrv4 I__8730 (
            .O(N__46171),
            .I(\c0.n20511 ));
    LocalMux I__8729 (
            .O(N__46168),
            .I(\c0.n20511 ));
    Odrv12 I__8728 (
            .O(N__46165),
            .I(\c0.n20511 ));
    CascadeMux I__8727 (
            .O(N__46158),
            .I(\c0.n10531_cascade_ ));
    InMux I__8726 (
            .O(N__46155),
            .I(N__46152));
    LocalMux I__8725 (
            .O(N__46152),
            .I(N__46148));
    InMux I__8724 (
            .O(N__46151),
            .I(N__46145));
    Odrv4 I__8723 (
            .O(N__46148),
            .I(\c0.n21451 ));
    LocalMux I__8722 (
            .O(N__46145),
            .I(\c0.n21451 ));
    CascadeMux I__8721 (
            .O(N__46140),
            .I(N__46136));
    InMux I__8720 (
            .O(N__46139),
            .I(N__46129));
    InMux I__8719 (
            .O(N__46136),
            .I(N__46122));
    InMux I__8718 (
            .O(N__46135),
            .I(N__46122));
    InMux I__8717 (
            .O(N__46134),
            .I(N__46122));
    InMux I__8716 (
            .O(N__46133),
            .I(N__46119));
    InMux I__8715 (
            .O(N__46132),
            .I(N__46116));
    LocalMux I__8714 (
            .O(N__46129),
            .I(N__46113));
    LocalMux I__8713 (
            .O(N__46122),
            .I(N__46106));
    LocalMux I__8712 (
            .O(N__46119),
            .I(N__46106));
    LocalMux I__8711 (
            .O(N__46116),
            .I(N__46106));
    Odrv4 I__8710 (
            .O(N__46113),
            .I(\c0.n21437 ));
    Odrv12 I__8709 (
            .O(N__46106),
            .I(\c0.n21437 ));
    CascadeMux I__8708 (
            .O(N__46101),
            .I(\c0.n21451_cascade_ ));
    InMux I__8707 (
            .O(N__46098),
            .I(N__46080));
    InMux I__8706 (
            .O(N__46097),
            .I(N__46071));
    InMux I__8705 (
            .O(N__46096),
            .I(N__46071));
    InMux I__8704 (
            .O(N__46095),
            .I(N__46071));
    InMux I__8703 (
            .O(N__46094),
            .I(N__46064));
    InMux I__8702 (
            .O(N__46093),
            .I(N__46064));
    InMux I__8701 (
            .O(N__46092),
            .I(N__46064));
    InMux I__8700 (
            .O(N__46091),
            .I(N__46052));
    InMux I__8699 (
            .O(N__46090),
            .I(N__46044));
    InMux I__8698 (
            .O(N__46089),
            .I(N__46041));
    InMux I__8697 (
            .O(N__46088),
            .I(N__46032));
    InMux I__8696 (
            .O(N__46087),
            .I(N__46032));
    InMux I__8695 (
            .O(N__46086),
            .I(N__46032));
    InMux I__8694 (
            .O(N__46085),
            .I(N__46032));
    InMux I__8693 (
            .O(N__46084),
            .I(N__46027));
    InMux I__8692 (
            .O(N__46083),
            .I(N__46015));
    LocalMux I__8691 (
            .O(N__46080),
            .I(N__46012));
    InMux I__8690 (
            .O(N__46079),
            .I(N__46005));
    InMux I__8689 (
            .O(N__46078),
            .I(N__46005));
    LocalMux I__8688 (
            .O(N__46071),
            .I(N__46002));
    LocalMux I__8687 (
            .O(N__46064),
            .I(N__45999));
    InMux I__8686 (
            .O(N__46063),
            .I(N__45972));
    InMux I__8685 (
            .O(N__46062),
            .I(N__45972));
    InMux I__8684 (
            .O(N__46061),
            .I(N__45972));
    InMux I__8683 (
            .O(N__46060),
            .I(N__45972));
    InMux I__8682 (
            .O(N__46059),
            .I(N__45972));
    InMux I__8681 (
            .O(N__46058),
            .I(N__45963));
    InMux I__8680 (
            .O(N__46057),
            .I(N__45963));
    InMux I__8679 (
            .O(N__46056),
            .I(N__45963));
    InMux I__8678 (
            .O(N__46055),
            .I(N__45963));
    LocalMux I__8677 (
            .O(N__46052),
            .I(N__45960));
    InMux I__8676 (
            .O(N__46051),
            .I(N__45949));
    InMux I__8675 (
            .O(N__46050),
            .I(N__45949));
    InMux I__8674 (
            .O(N__46049),
            .I(N__45949));
    InMux I__8673 (
            .O(N__46048),
            .I(N__45949));
    InMux I__8672 (
            .O(N__46047),
            .I(N__45949));
    LocalMux I__8671 (
            .O(N__46044),
            .I(N__45946));
    LocalMux I__8670 (
            .O(N__46041),
            .I(N__45940));
    LocalMux I__8669 (
            .O(N__46032),
            .I(N__45940));
    InMux I__8668 (
            .O(N__46031),
            .I(N__45937));
    InMux I__8667 (
            .O(N__46030),
            .I(N__45933));
    LocalMux I__8666 (
            .O(N__46027),
            .I(N__45930));
    InMux I__8665 (
            .O(N__46026),
            .I(N__45927));
    InMux I__8664 (
            .O(N__46025),
            .I(N__45922));
    InMux I__8663 (
            .O(N__46024),
            .I(N__45922));
    InMux I__8662 (
            .O(N__46023),
            .I(N__45919));
    InMux I__8661 (
            .O(N__46022),
            .I(N__45914));
    InMux I__8660 (
            .O(N__46021),
            .I(N__45914));
    InMux I__8659 (
            .O(N__46020),
            .I(N__45907));
    InMux I__8658 (
            .O(N__46019),
            .I(N__45907));
    InMux I__8657 (
            .O(N__46018),
            .I(N__45907));
    LocalMux I__8656 (
            .O(N__46015),
            .I(N__45902));
    Span4Mux_h I__8655 (
            .O(N__46012),
            .I(N__45902));
    InMux I__8654 (
            .O(N__46011),
            .I(N__45897));
    InMux I__8653 (
            .O(N__46010),
            .I(N__45897));
    LocalMux I__8652 (
            .O(N__46005),
            .I(N__45890));
    Span4Mux_h I__8651 (
            .O(N__46002),
            .I(N__45890));
    Span4Mux_h I__8650 (
            .O(N__45999),
            .I(N__45890));
    CascadeMux I__8649 (
            .O(N__45998),
            .I(N__45886));
    CascadeMux I__8648 (
            .O(N__45997),
            .I(N__45883));
    InMux I__8647 (
            .O(N__45996),
            .I(N__45864));
    InMux I__8646 (
            .O(N__45995),
            .I(N__45864));
    InMux I__8645 (
            .O(N__45994),
            .I(N__45864));
    InMux I__8644 (
            .O(N__45993),
            .I(N__45859));
    InMux I__8643 (
            .O(N__45992),
            .I(N__45859));
    InMux I__8642 (
            .O(N__45991),
            .I(N__45852));
    InMux I__8641 (
            .O(N__45990),
            .I(N__45852));
    InMux I__8640 (
            .O(N__45989),
            .I(N__45852));
    InMux I__8639 (
            .O(N__45988),
            .I(N__45839));
    InMux I__8638 (
            .O(N__45987),
            .I(N__45839));
    InMux I__8637 (
            .O(N__45986),
            .I(N__45839));
    InMux I__8636 (
            .O(N__45985),
            .I(N__45839));
    InMux I__8635 (
            .O(N__45984),
            .I(N__45839));
    InMux I__8634 (
            .O(N__45983),
            .I(N__45839));
    LocalMux I__8633 (
            .O(N__45972),
            .I(N__45832));
    LocalMux I__8632 (
            .O(N__45963),
            .I(N__45832));
    Span4Mux_v I__8631 (
            .O(N__45960),
            .I(N__45832));
    LocalMux I__8630 (
            .O(N__45949),
            .I(N__45827));
    Span4Mux_v I__8629 (
            .O(N__45946),
            .I(N__45827));
    InMux I__8628 (
            .O(N__45945),
            .I(N__45824));
    Span4Mux_v I__8627 (
            .O(N__45940),
            .I(N__45821));
    LocalMux I__8626 (
            .O(N__45937),
            .I(N__45818));
    InMux I__8625 (
            .O(N__45936),
            .I(N__45815));
    LocalMux I__8624 (
            .O(N__45933),
            .I(N__45812));
    Span4Mux_v I__8623 (
            .O(N__45930),
            .I(N__45809));
    LocalMux I__8622 (
            .O(N__45927),
            .I(N__45796));
    LocalMux I__8621 (
            .O(N__45922),
            .I(N__45796));
    LocalMux I__8620 (
            .O(N__45919),
            .I(N__45796));
    LocalMux I__8619 (
            .O(N__45914),
            .I(N__45796));
    LocalMux I__8618 (
            .O(N__45907),
            .I(N__45796));
    Span4Mux_v I__8617 (
            .O(N__45902),
            .I(N__45796));
    LocalMux I__8616 (
            .O(N__45897),
            .I(N__45791));
    Span4Mux_v I__8615 (
            .O(N__45890),
            .I(N__45791));
    InMux I__8614 (
            .O(N__45889),
            .I(N__45788));
    InMux I__8613 (
            .O(N__45886),
            .I(N__45785));
    InMux I__8612 (
            .O(N__45883),
            .I(N__45782));
    InMux I__8611 (
            .O(N__45882),
            .I(N__45775));
    InMux I__8610 (
            .O(N__45881),
            .I(N__45775));
    InMux I__8609 (
            .O(N__45880),
            .I(N__45775));
    InMux I__8608 (
            .O(N__45879),
            .I(N__45766));
    InMux I__8607 (
            .O(N__45878),
            .I(N__45766));
    InMux I__8606 (
            .O(N__45877),
            .I(N__45766));
    InMux I__8605 (
            .O(N__45876),
            .I(N__45766));
    InMux I__8604 (
            .O(N__45875),
            .I(N__45755));
    InMux I__8603 (
            .O(N__45874),
            .I(N__45755));
    InMux I__8602 (
            .O(N__45873),
            .I(N__45755));
    InMux I__8601 (
            .O(N__45872),
            .I(N__45755));
    InMux I__8600 (
            .O(N__45871),
            .I(N__45755));
    LocalMux I__8599 (
            .O(N__45864),
            .I(N__45752));
    LocalMux I__8598 (
            .O(N__45859),
            .I(N__45741));
    LocalMux I__8597 (
            .O(N__45852),
            .I(N__45741));
    LocalMux I__8596 (
            .O(N__45839),
            .I(N__45741));
    Span4Mux_h I__8595 (
            .O(N__45832),
            .I(N__45741));
    Span4Mux_h I__8594 (
            .O(N__45827),
            .I(N__45741));
    LocalMux I__8593 (
            .O(N__45824),
            .I(N__45734));
    Sp12to4 I__8592 (
            .O(N__45821),
            .I(N__45734));
    Span12Mux_v I__8591 (
            .O(N__45818),
            .I(N__45734));
    LocalMux I__8590 (
            .O(N__45815),
            .I(N__45723));
    Span4Mux_v I__8589 (
            .O(N__45812),
            .I(N__45723));
    Span4Mux_h I__8588 (
            .O(N__45809),
            .I(N__45723));
    Span4Mux_v I__8587 (
            .O(N__45796),
            .I(N__45723));
    Span4Mux_v I__8586 (
            .O(N__45791),
            .I(N__45723));
    LocalMux I__8585 (
            .O(N__45788),
            .I(N__45718));
    LocalMux I__8584 (
            .O(N__45785),
            .I(N__45718));
    LocalMux I__8583 (
            .O(N__45782),
            .I(n13058));
    LocalMux I__8582 (
            .O(N__45775),
            .I(n13058));
    LocalMux I__8581 (
            .O(N__45766),
            .I(n13058));
    LocalMux I__8580 (
            .O(N__45755),
            .I(n13058));
    Odrv12 I__8579 (
            .O(N__45752),
            .I(n13058));
    Odrv4 I__8578 (
            .O(N__45741),
            .I(n13058));
    Odrv12 I__8577 (
            .O(N__45734),
            .I(n13058));
    Odrv4 I__8576 (
            .O(N__45723),
            .I(n13058));
    Odrv4 I__8575 (
            .O(N__45718),
            .I(n13058));
    InMux I__8574 (
            .O(N__45699),
            .I(N__45696));
    LocalMux I__8573 (
            .O(N__45696),
            .I(N__45693));
    Span4Mux_v I__8572 (
            .O(N__45693),
            .I(N__45689));
    CascadeMux I__8571 (
            .O(N__45692),
            .I(N__45686));
    Span4Mux_h I__8570 (
            .O(N__45689),
            .I(N__45683));
    InMux I__8569 (
            .O(N__45686),
            .I(N__45680));
    Span4Mux_v I__8568 (
            .O(N__45683),
            .I(N__45677));
    LocalMux I__8567 (
            .O(N__45680),
            .I(data_out_frame_8_6));
    Odrv4 I__8566 (
            .O(N__45677),
            .I(data_out_frame_8_6));
    CascadeMux I__8565 (
            .O(N__45672),
            .I(N__45669));
    InMux I__8564 (
            .O(N__45669),
            .I(N__45666));
    LocalMux I__8563 (
            .O(N__45666),
            .I(N__45663));
    Span4Mux_h I__8562 (
            .O(N__45663),
            .I(N__45660));
    Span4Mux_v I__8561 (
            .O(N__45660),
            .I(N__45657));
    Span4Mux_h I__8560 (
            .O(N__45657),
            .I(N__45652));
    CascadeMux I__8559 (
            .O(N__45656),
            .I(N__45649));
    InMux I__8558 (
            .O(N__45655),
            .I(N__45645));
    Span4Mux_v I__8557 (
            .O(N__45652),
            .I(N__45642));
    InMux I__8556 (
            .O(N__45649),
            .I(N__45639));
    InMux I__8555 (
            .O(N__45648),
            .I(N__45636));
    LocalMux I__8554 (
            .O(N__45645),
            .I(encoder0_position_21));
    Odrv4 I__8553 (
            .O(N__45642),
            .I(encoder0_position_21));
    LocalMux I__8552 (
            .O(N__45639),
            .I(encoder0_position_21));
    LocalMux I__8551 (
            .O(N__45636),
            .I(encoder0_position_21));
    InMux I__8550 (
            .O(N__45627),
            .I(N__45623));
    InMux I__8549 (
            .O(N__45626),
            .I(N__45620));
    LocalMux I__8548 (
            .O(N__45623),
            .I(\c0.n22252 ));
    LocalMux I__8547 (
            .O(N__45620),
            .I(\c0.n22252 ));
    CascadeMux I__8546 (
            .O(N__45615),
            .I(N__45609));
    CascadeMux I__8545 (
            .O(N__45614),
            .I(N__45606));
    CascadeMux I__8544 (
            .O(N__45613),
            .I(N__45603));
    InMux I__8543 (
            .O(N__45612),
            .I(N__45599));
    InMux I__8542 (
            .O(N__45609),
            .I(N__45595));
    InMux I__8541 (
            .O(N__45606),
            .I(N__45592));
    InMux I__8540 (
            .O(N__45603),
            .I(N__45588));
    InMux I__8539 (
            .O(N__45602),
            .I(N__45584));
    LocalMux I__8538 (
            .O(N__45599),
            .I(N__45581));
    InMux I__8537 (
            .O(N__45598),
            .I(N__45578));
    LocalMux I__8536 (
            .O(N__45595),
            .I(N__45573));
    LocalMux I__8535 (
            .O(N__45592),
            .I(N__45573));
    InMux I__8534 (
            .O(N__45591),
            .I(N__45570));
    LocalMux I__8533 (
            .O(N__45588),
            .I(N__45567));
    InMux I__8532 (
            .O(N__45587),
            .I(N__45564));
    LocalMux I__8531 (
            .O(N__45584),
            .I(N__45561));
    Span4Mux_v I__8530 (
            .O(N__45581),
            .I(N__45556));
    LocalMux I__8529 (
            .O(N__45578),
            .I(N__45556));
    Span4Mux_h I__8528 (
            .O(N__45573),
            .I(N__45549));
    LocalMux I__8527 (
            .O(N__45570),
            .I(N__45549));
    Span4Mux_h I__8526 (
            .O(N__45567),
            .I(N__45549));
    LocalMux I__8525 (
            .O(N__45564),
            .I(encoder0_position_27));
    Odrv12 I__8524 (
            .O(N__45561),
            .I(encoder0_position_27));
    Odrv4 I__8523 (
            .O(N__45556),
            .I(encoder0_position_27));
    Odrv4 I__8522 (
            .O(N__45549),
            .I(encoder0_position_27));
    InMux I__8521 (
            .O(N__45540),
            .I(N__45537));
    LocalMux I__8520 (
            .O(N__45537),
            .I(N__45534));
    Span4Mux_v I__8519 (
            .O(N__45534),
            .I(N__45530));
    InMux I__8518 (
            .O(N__45533),
            .I(N__45527));
    Span4Mux_h I__8517 (
            .O(N__45530),
            .I(N__45524));
    LocalMux I__8516 (
            .O(N__45527),
            .I(data_out_frame_6_3));
    Odrv4 I__8515 (
            .O(N__45524),
            .I(data_out_frame_6_3));
    InMux I__8514 (
            .O(N__45519),
            .I(N__45514));
    InMux I__8513 (
            .O(N__45518),
            .I(N__45511));
    CascadeMux I__8512 (
            .O(N__45517),
            .I(N__45508));
    LocalMux I__8511 (
            .O(N__45514),
            .I(N__45502));
    LocalMux I__8510 (
            .O(N__45511),
            .I(N__45499));
    InMux I__8509 (
            .O(N__45508),
            .I(N__45494));
    InMux I__8508 (
            .O(N__45507),
            .I(N__45494));
    InMux I__8507 (
            .O(N__45506),
            .I(N__45490));
    InMux I__8506 (
            .O(N__45505),
            .I(N__45487));
    Span4Mux_v I__8505 (
            .O(N__45502),
            .I(N__45480));
    Span4Mux_h I__8504 (
            .O(N__45499),
            .I(N__45480));
    LocalMux I__8503 (
            .O(N__45494),
            .I(N__45480));
    InMux I__8502 (
            .O(N__45493),
            .I(N__45476));
    LocalMux I__8501 (
            .O(N__45490),
            .I(N__45473));
    LocalMux I__8500 (
            .O(N__45487),
            .I(N__45470));
    Span4Mux_v I__8499 (
            .O(N__45480),
            .I(N__45467));
    InMux I__8498 (
            .O(N__45479),
            .I(N__45464));
    LocalMux I__8497 (
            .O(N__45476),
            .I(N__45461));
    Span12Mux_s7_v I__8496 (
            .O(N__45473),
            .I(N__45458));
    Span4Mux_v I__8495 (
            .O(N__45470),
            .I(N__45453));
    Span4Mux_h I__8494 (
            .O(N__45467),
            .I(N__45453));
    LocalMux I__8493 (
            .O(N__45464),
            .I(encoder1_position_3));
    Odrv4 I__8492 (
            .O(N__45461),
            .I(encoder1_position_3));
    Odrv12 I__8491 (
            .O(N__45458),
            .I(encoder1_position_3));
    Odrv4 I__8490 (
            .O(N__45453),
            .I(encoder1_position_3));
    InMux I__8489 (
            .O(N__45444),
            .I(N__45441));
    LocalMux I__8488 (
            .O(N__45441),
            .I(N__45433));
    InMux I__8487 (
            .O(N__45440),
            .I(N__45430));
    InMux I__8486 (
            .O(N__45439),
            .I(N__45425));
    InMux I__8485 (
            .O(N__45438),
            .I(N__45425));
    InMux I__8484 (
            .O(N__45437),
            .I(N__45422));
    InMux I__8483 (
            .O(N__45436),
            .I(N__45419));
    Span4Mux_v I__8482 (
            .O(N__45433),
            .I(N__45416));
    LocalMux I__8481 (
            .O(N__45430),
            .I(N__45411));
    LocalMux I__8480 (
            .O(N__45425),
            .I(N__45411));
    LocalMux I__8479 (
            .O(N__45422),
            .I(N__45408));
    LocalMux I__8478 (
            .O(N__45419),
            .I(\c0.n20455 ));
    Odrv4 I__8477 (
            .O(N__45416),
            .I(\c0.n20455 ));
    Odrv12 I__8476 (
            .O(N__45411),
            .I(\c0.n20455 ));
    Odrv4 I__8475 (
            .O(N__45408),
            .I(\c0.n20455 ));
    InMux I__8474 (
            .O(N__45399),
            .I(N__45396));
    LocalMux I__8473 (
            .O(N__45396),
            .I(N__45393));
    Span4Mux_v I__8472 (
            .O(N__45393),
            .I(N__45389));
    InMux I__8471 (
            .O(N__45392),
            .I(N__45386));
    Span4Mux_h I__8470 (
            .O(N__45389),
            .I(N__45383));
    LocalMux I__8469 (
            .O(N__45386),
            .I(N__45377));
    Span4Mux_v I__8468 (
            .O(N__45383),
            .I(N__45374));
    InMux I__8467 (
            .O(N__45382),
            .I(N__45371));
    InMux I__8466 (
            .O(N__45381),
            .I(N__45368));
    InMux I__8465 (
            .O(N__45380),
            .I(N__45365));
    Span4Mux_v I__8464 (
            .O(N__45377),
            .I(N__45362));
    Sp12to4 I__8463 (
            .O(N__45374),
            .I(N__45357));
    LocalMux I__8462 (
            .O(N__45371),
            .I(N__45357));
    LocalMux I__8461 (
            .O(N__45368),
            .I(encoder0_position_5));
    LocalMux I__8460 (
            .O(N__45365),
            .I(encoder0_position_5));
    Odrv4 I__8459 (
            .O(N__45362),
            .I(encoder0_position_5));
    Odrv12 I__8458 (
            .O(N__45357),
            .I(encoder0_position_5));
    InMux I__8457 (
            .O(N__45348),
            .I(N__45345));
    LocalMux I__8456 (
            .O(N__45345),
            .I(N__45341));
    CascadeMux I__8455 (
            .O(N__45344),
            .I(N__45337));
    Span4Mux_h I__8454 (
            .O(N__45341),
            .I(N__45333));
    InMux I__8453 (
            .O(N__45340),
            .I(N__45330));
    InMux I__8452 (
            .O(N__45337),
            .I(N__45327));
    InMux I__8451 (
            .O(N__45336),
            .I(N__45324));
    Span4Mux_v I__8450 (
            .O(N__45333),
            .I(N__45316));
    LocalMux I__8449 (
            .O(N__45330),
            .I(N__45316));
    LocalMux I__8448 (
            .O(N__45327),
            .I(N__45311));
    LocalMux I__8447 (
            .O(N__45324),
            .I(N__45311));
    CascadeMux I__8446 (
            .O(N__45323),
            .I(N__45308));
    InMux I__8445 (
            .O(N__45322),
            .I(N__45305));
    InMux I__8444 (
            .O(N__45321),
            .I(N__45302));
    Span4Mux_v I__8443 (
            .O(N__45316),
            .I(N__45297));
    Span4Mux_h I__8442 (
            .O(N__45311),
            .I(N__45297));
    InMux I__8441 (
            .O(N__45308),
            .I(N__45294));
    LocalMux I__8440 (
            .O(N__45305),
            .I(encoder0_position_20));
    LocalMux I__8439 (
            .O(N__45302),
            .I(encoder0_position_20));
    Odrv4 I__8438 (
            .O(N__45297),
            .I(encoder0_position_20));
    LocalMux I__8437 (
            .O(N__45294),
            .I(encoder0_position_20));
    CascadeMux I__8436 (
            .O(N__45285),
            .I(N__45282));
    InMux I__8435 (
            .O(N__45282),
            .I(N__45279));
    LocalMux I__8434 (
            .O(N__45279),
            .I(\c0.n22689 ));
    InMux I__8433 (
            .O(N__45276),
            .I(N__45273));
    LocalMux I__8432 (
            .O(N__45273),
            .I(N__45270));
    Odrv4 I__8431 (
            .O(N__45270),
            .I(\c0.n22641 ));
    CascadeMux I__8430 (
            .O(N__45267),
            .I(N__45264));
    InMux I__8429 (
            .O(N__45264),
            .I(N__45257));
    InMux I__8428 (
            .O(N__45263),
            .I(N__45254));
    InMux I__8427 (
            .O(N__45262),
            .I(N__45251));
    InMux I__8426 (
            .O(N__45261),
            .I(N__45248));
    InMux I__8425 (
            .O(N__45260),
            .I(N__45245));
    LocalMux I__8424 (
            .O(N__45257),
            .I(N__45242));
    LocalMux I__8423 (
            .O(N__45254),
            .I(N__45239));
    LocalMux I__8422 (
            .O(N__45251),
            .I(N__45236));
    LocalMux I__8421 (
            .O(N__45248),
            .I(N__45233));
    LocalMux I__8420 (
            .O(N__45245),
            .I(N__45230));
    Span4Mux_v I__8419 (
            .O(N__45242),
            .I(N__45219));
    Span4Mux_v I__8418 (
            .O(N__45239),
            .I(N__45219));
    Span4Mux_h I__8417 (
            .O(N__45236),
            .I(N__45219));
    Span4Mux_v I__8416 (
            .O(N__45233),
            .I(N__45219));
    Span4Mux_v I__8415 (
            .O(N__45230),
            .I(N__45216));
    InMux I__8414 (
            .O(N__45229),
            .I(N__45213));
    InMux I__8413 (
            .O(N__45228),
            .I(N__45210));
    Span4Mux_h I__8412 (
            .O(N__45219),
            .I(N__45207));
    Span4Mux_h I__8411 (
            .O(N__45216),
            .I(N__45204));
    LocalMux I__8410 (
            .O(N__45213),
            .I(N__45201));
    LocalMux I__8409 (
            .O(N__45210),
            .I(encoder0_position_4));
    Odrv4 I__8408 (
            .O(N__45207),
            .I(encoder0_position_4));
    Odrv4 I__8407 (
            .O(N__45204),
            .I(encoder0_position_4));
    Odrv4 I__8406 (
            .O(N__45201),
            .I(encoder0_position_4));
    CascadeMux I__8405 (
            .O(N__45192),
            .I(\c0.n22689_cascade_ ));
    CascadeMux I__8404 (
            .O(N__45189),
            .I(N__45186));
    InMux I__8403 (
            .O(N__45186),
            .I(N__45181));
    InMux I__8402 (
            .O(N__45185),
            .I(N__45178));
    InMux I__8401 (
            .O(N__45184),
            .I(N__45175));
    LocalMux I__8400 (
            .O(N__45181),
            .I(N__45170));
    LocalMux I__8399 (
            .O(N__45178),
            .I(N__45165));
    LocalMux I__8398 (
            .O(N__45175),
            .I(N__45165));
    InMux I__8397 (
            .O(N__45174),
            .I(N__45162));
    InMux I__8396 (
            .O(N__45173),
            .I(N__45159));
    Span4Mux_h I__8395 (
            .O(N__45170),
            .I(N__45155));
    Span4Mux_v I__8394 (
            .O(N__45165),
            .I(N__45152));
    LocalMux I__8393 (
            .O(N__45162),
            .I(N__45149));
    LocalMux I__8392 (
            .O(N__45159),
            .I(N__45146));
    InMux I__8391 (
            .O(N__45158),
            .I(N__45143));
    Span4Mux_h I__8390 (
            .O(N__45155),
            .I(N__45140));
    Span4Mux_v I__8389 (
            .O(N__45152),
            .I(N__45137));
    Span12Mux_h I__8388 (
            .O(N__45149),
            .I(N__45132));
    Span12Mux_v I__8387 (
            .O(N__45146),
            .I(N__45132));
    LocalMux I__8386 (
            .O(N__45143),
            .I(control_mode_0));
    Odrv4 I__8385 (
            .O(N__45140),
            .I(control_mode_0));
    Odrv4 I__8384 (
            .O(N__45137),
            .I(control_mode_0));
    Odrv12 I__8383 (
            .O(N__45132),
            .I(control_mode_0));
    InMux I__8382 (
            .O(N__45123),
            .I(N__45120));
    LocalMux I__8381 (
            .O(N__45120),
            .I(N__45117));
    Span4Mux_h I__8380 (
            .O(N__45117),
            .I(N__45113));
    InMux I__8379 (
            .O(N__45116),
            .I(N__45110));
    Odrv4 I__8378 (
            .O(N__45113),
            .I(\c0.n10455 ));
    LocalMux I__8377 (
            .O(N__45110),
            .I(\c0.n10455 ));
    InMux I__8376 (
            .O(N__45105),
            .I(N__45102));
    LocalMux I__8375 (
            .O(N__45102),
            .I(N__45099));
    Span4Mux_h I__8374 (
            .O(N__45099),
            .I(N__45095));
    InMux I__8373 (
            .O(N__45098),
            .I(N__45092));
    Odrv4 I__8372 (
            .O(N__45095),
            .I(\c0.n20312 ));
    LocalMux I__8371 (
            .O(N__45092),
            .I(\c0.n20312 ));
    CascadeMux I__8370 (
            .O(N__45087),
            .I(\c0.n20312_cascade_ ));
    InMux I__8369 (
            .O(N__45084),
            .I(N__45081));
    LocalMux I__8368 (
            .O(N__45081),
            .I(\c0.n22522 ));
    CascadeMux I__8367 (
            .O(N__45078),
            .I(\c0.n6_adj_4674_cascade_ ));
    InMux I__8366 (
            .O(N__45075),
            .I(N__45072));
    LocalMux I__8365 (
            .O(N__45072),
            .I(N__45069));
    Span4Mux_h I__8364 (
            .O(N__45069),
            .I(N__45066));
    Span4Mux_h I__8363 (
            .O(N__45066),
            .I(N__45063));
    Odrv4 I__8362 (
            .O(N__45063),
            .I(\c0.data_out_frame_29_4 ));
    CEMux I__8361 (
            .O(N__45060),
            .I(N__45056));
    CEMux I__8360 (
            .O(N__45059),
            .I(N__45051));
    LocalMux I__8359 (
            .O(N__45056),
            .I(N__45047));
    CEMux I__8358 (
            .O(N__45055),
            .I(N__45044));
    CEMux I__8357 (
            .O(N__45054),
            .I(N__45038));
    LocalMux I__8356 (
            .O(N__45051),
            .I(N__45032));
    CEMux I__8355 (
            .O(N__45050),
            .I(N__45029));
    Span4Mux_h I__8354 (
            .O(N__45047),
            .I(N__45022));
    LocalMux I__8353 (
            .O(N__45044),
            .I(N__45022));
    CEMux I__8352 (
            .O(N__45043),
            .I(N__45019));
    CEMux I__8351 (
            .O(N__45042),
            .I(N__45016));
    CEMux I__8350 (
            .O(N__45041),
            .I(N__45013));
    LocalMux I__8349 (
            .O(N__45038),
            .I(N__45010));
    CEMux I__8348 (
            .O(N__45037),
            .I(N__45007));
    CEMux I__8347 (
            .O(N__45036),
            .I(N__45004));
    CEMux I__8346 (
            .O(N__45035),
            .I(N__45001));
    Span4Mux_v I__8345 (
            .O(N__45032),
            .I(N__44996));
    LocalMux I__8344 (
            .O(N__45029),
            .I(N__44996));
    SRMux I__8343 (
            .O(N__45028),
            .I(N__44992));
    SRMux I__8342 (
            .O(N__45027),
            .I(N__44989));
    Span4Mux_h I__8341 (
            .O(N__45022),
            .I(N__44986));
    LocalMux I__8340 (
            .O(N__45019),
            .I(N__44983));
    LocalMux I__8339 (
            .O(N__45016),
            .I(N__44980));
    LocalMux I__8338 (
            .O(N__45013),
            .I(N__44975));
    Span4Mux_h I__8337 (
            .O(N__45010),
            .I(N__44975));
    LocalMux I__8336 (
            .O(N__45007),
            .I(N__44972));
    LocalMux I__8335 (
            .O(N__45004),
            .I(N__44967));
    LocalMux I__8334 (
            .O(N__45001),
            .I(N__44967));
    Span4Mux_h I__8333 (
            .O(N__44996),
            .I(N__44964));
    SRMux I__8332 (
            .O(N__44995),
            .I(N__44961));
    LocalMux I__8331 (
            .O(N__44992),
            .I(N__44956));
    LocalMux I__8330 (
            .O(N__44989),
            .I(N__44956));
    Span4Mux_v I__8329 (
            .O(N__44986),
            .I(N__44953));
    Span4Mux_v I__8328 (
            .O(N__44983),
            .I(N__44948));
    Span4Mux_v I__8327 (
            .O(N__44980),
            .I(N__44948));
    Span4Mux_v I__8326 (
            .O(N__44975),
            .I(N__44945));
    Span4Mux_h I__8325 (
            .O(N__44972),
            .I(N__44938));
    Span4Mux_h I__8324 (
            .O(N__44967),
            .I(N__44938));
    Span4Mux_h I__8323 (
            .O(N__44964),
            .I(N__44938));
    LocalMux I__8322 (
            .O(N__44961),
            .I(N__44931));
    Span4Mux_v I__8321 (
            .O(N__44956),
            .I(N__44931));
    Span4Mux_h I__8320 (
            .O(N__44953),
            .I(N__44931));
    Span4Mux_v I__8319 (
            .O(N__44948),
            .I(N__44926));
    Span4Mux_v I__8318 (
            .O(N__44945),
            .I(N__44926));
    Sp12to4 I__8317 (
            .O(N__44938),
            .I(N__44923));
    Span4Mux_v I__8316 (
            .O(N__44931),
            .I(N__44920));
    Span4Mux_h I__8315 (
            .O(N__44926),
            .I(N__44917));
    Odrv12 I__8314 (
            .O(N__44923),
            .I(\c0.n8162 ));
    Odrv4 I__8313 (
            .O(N__44920),
            .I(\c0.n8162 ));
    Odrv4 I__8312 (
            .O(N__44917),
            .I(\c0.n8162 ));
    InMux I__8311 (
            .O(N__44910),
            .I(N__44907));
    LocalMux I__8310 (
            .O(N__44907),
            .I(N__44904));
    Odrv4 I__8309 (
            .O(N__44904),
            .I(\c0.n22580 ));
    InMux I__8308 (
            .O(N__44901),
            .I(N__44896));
    InMux I__8307 (
            .O(N__44900),
            .I(N__44891));
    InMux I__8306 (
            .O(N__44899),
            .I(N__44891));
    LocalMux I__8305 (
            .O(N__44896),
            .I(N__44888));
    LocalMux I__8304 (
            .O(N__44891),
            .I(N__44883));
    Span4Mux_h I__8303 (
            .O(N__44888),
            .I(N__44883));
    Odrv4 I__8302 (
            .O(N__44883),
            .I(\c0.n10477 ));
    InMux I__8301 (
            .O(N__44880),
            .I(N__44877));
    LocalMux I__8300 (
            .O(N__44877),
            .I(N__44874));
    Odrv4 I__8299 (
            .O(N__44874),
            .I(n2339));
    CascadeMux I__8298 (
            .O(N__44871),
            .I(N__44868));
    InMux I__8297 (
            .O(N__44868),
            .I(N__44865));
    LocalMux I__8296 (
            .O(N__44865),
            .I(N__44858));
    InMux I__8295 (
            .O(N__44864),
            .I(N__44855));
    CascadeMux I__8294 (
            .O(N__44863),
            .I(N__44852));
    InMux I__8293 (
            .O(N__44862),
            .I(N__44847));
    InMux I__8292 (
            .O(N__44861),
            .I(N__44847));
    Span4Mux_h I__8291 (
            .O(N__44858),
            .I(N__44841));
    LocalMux I__8290 (
            .O(N__44855),
            .I(N__44841));
    InMux I__8289 (
            .O(N__44852),
            .I(N__44838));
    LocalMux I__8288 (
            .O(N__44847),
            .I(N__44835));
    CascadeMux I__8287 (
            .O(N__44846),
            .I(N__44832));
    Span4Mux_v I__8286 (
            .O(N__44841),
            .I(N__44827));
    LocalMux I__8285 (
            .O(N__44838),
            .I(N__44822));
    Span4Mux_v I__8284 (
            .O(N__44835),
            .I(N__44822));
    InMux I__8283 (
            .O(N__44832),
            .I(N__44815));
    InMux I__8282 (
            .O(N__44831),
            .I(N__44815));
    InMux I__8281 (
            .O(N__44830),
            .I(N__44815));
    Odrv4 I__8280 (
            .O(N__44827),
            .I(encoder0_position_18));
    Odrv4 I__8279 (
            .O(N__44822),
            .I(encoder0_position_18));
    LocalMux I__8278 (
            .O(N__44815),
            .I(encoder0_position_18));
    InMux I__8277 (
            .O(N__44808),
            .I(N__44805));
    LocalMux I__8276 (
            .O(N__44805),
            .I(\c0.n22583 ));
    CascadeMux I__8275 (
            .O(N__44802),
            .I(N__44799));
    InMux I__8274 (
            .O(N__44799),
            .I(N__44793));
    InMux I__8273 (
            .O(N__44798),
            .I(N__44793));
    LocalMux I__8272 (
            .O(N__44793),
            .I(N__44790));
    Sp12to4 I__8271 (
            .O(N__44790),
            .I(N__44787));
    Span12Mux_s9_v I__8270 (
            .O(N__44787),
            .I(N__44784));
    Odrv12 I__8269 (
            .O(N__44784),
            .I(\c0.n22149 ));
    CascadeMux I__8268 (
            .O(N__44781),
            .I(N__44778));
    InMux I__8267 (
            .O(N__44778),
            .I(N__44775));
    LocalMux I__8266 (
            .O(N__44775),
            .I(N__44770));
    InMux I__8265 (
            .O(N__44774),
            .I(N__44766));
    InMux I__8264 (
            .O(N__44773),
            .I(N__44763));
    Span4Mux_v I__8263 (
            .O(N__44770),
            .I(N__44759));
    InMux I__8262 (
            .O(N__44769),
            .I(N__44756));
    LocalMux I__8261 (
            .O(N__44766),
            .I(N__44750));
    LocalMux I__8260 (
            .O(N__44763),
            .I(N__44750));
    CascadeMux I__8259 (
            .O(N__44762),
            .I(N__44747));
    Span4Mux_v I__8258 (
            .O(N__44759),
            .I(N__44744));
    LocalMux I__8257 (
            .O(N__44756),
            .I(N__44741));
    InMux I__8256 (
            .O(N__44755),
            .I(N__44738));
    Span4Mux_v I__8255 (
            .O(N__44750),
            .I(N__44735));
    InMux I__8254 (
            .O(N__44747),
            .I(N__44732));
    Span4Mux_h I__8253 (
            .O(N__44744),
            .I(N__44727));
    Span4Mux_v I__8252 (
            .O(N__44741),
            .I(N__44727));
    LocalMux I__8251 (
            .O(N__44738),
            .I(encoder0_position_3));
    Odrv4 I__8250 (
            .O(N__44735),
            .I(encoder0_position_3));
    LocalMux I__8249 (
            .O(N__44732),
            .I(encoder0_position_3));
    Odrv4 I__8248 (
            .O(N__44727),
            .I(encoder0_position_3));
    CascadeMux I__8247 (
            .O(N__44718),
            .I(\c0.n22583_cascade_ ));
    CascadeMux I__8246 (
            .O(N__44715),
            .I(N__44712));
    InMux I__8245 (
            .O(N__44712),
            .I(N__44709));
    LocalMux I__8244 (
            .O(N__44709),
            .I(N__44704));
    InMux I__8243 (
            .O(N__44708),
            .I(N__44700));
    InMux I__8242 (
            .O(N__44707),
            .I(N__44696));
    Span4Mux_v I__8241 (
            .O(N__44704),
            .I(N__44693));
    InMux I__8240 (
            .O(N__44703),
            .I(N__44690));
    LocalMux I__8239 (
            .O(N__44700),
            .I(N__44687));
    InMux I__8238 (
            .O(N__44699),
            .I(N__44680));
    LocalMux I__8237 (
            .O(N__44696),
            .I(N__44677));
    Span4Mux_v I__8236 (
            .O(N__44693),
            .I(N__44674));
    LocalMux I__8235 (
            .O(N__44690),
            .I(N__44671));
    Span4Mux_v I__8234 (
            .O(N__44687),
            .I(N__44668));
    InMux I__8233 (
            .O(N__44686),
            .I(N__44665));
    InMux I__8232 (
            .O(N__44685),
            .I(N__44660));
    InMux I__8231 (
            .O(N__44684),
            .I(N__44660));
    InMux I__8230 (
            .O(N__44683),
            .I(N__44657));
    LocalMux I__8229 (
            .O(N__44680),
            .I(N__44652));
    Span4Mux_h I__8228 (
            .O(N__44677),
            .I(N__44652));
    Span4Mux_h I__8227 (
            .O(N__44674),
            .I(N__44645));
    Span4Mux_v I__8226 (
            .O(N__44671),
            .I(N__44645));
    Span4Mux_v I__8225 (
            .O(N__44668),
            .I(N__44645));
    LocalMux I__8224 (
            .O(N__44665),
            .I(N__44642));
    LocalMux I__8223 (
            .O(N__44660),
            .I(encoder0_position_31));
    LocalMux I__8222 (
            .O(N__44657),
            .I(encoder0_position_31));
    Odrv4 I__8221 (
            .O(N__44652),
            .I(encoder0_position_31));
    Odrv4 I__8220 (
            .O(N__44645),
            .I(encoder0_position_31));
    Odrv4 I__8219 (
            .O(N__44642),
            .I(encoder0_position_31));
    CascadeMux I__8218 (
            .O(N__44631),
            .I(N__44628));
    InMux I__8217 (
            .O(N__44628),
            .I(N__44623));
    InMux I__8216 (
            .O(N__44627),
            .I(N__44618));
    InMux I__8215 (
            .O(N__44626),
            .I(N__44618));
    LocalMux I__8214 (
            .O(N__44623),
            .I(N__44613));
    LocalMux I__8213 (
            .O(N__44618),
            .I(N__44613));
    Span4Mux_h I__8212 (
            .O(N__44613),
            .I(N__44610));
    Odrv4 I__8211 (
            .O(N__44610),
            .I(\c0.n13872 ));
    CascadeMux I__8210 (
            .O(N__44607),
            .I(N__44604));
    InMux I__8209 (
            .O(N__44604),
            .I(N__44601));
    LocalMux I__8208 (
            .O(N__44601),
            .I(N__44598));
    Span4Mux_v I__8207 (
            .O(N__44598),
            .I(N__44595));
    Span4Mux_v I__8206 (
            .O(N__44595),
            .I(N__44592));
    Odrv4 I__8205 (
            .O(N__44592),
            .I(n2337));
    InMux I__8204 (
            .O(N__44589),
            .I(N__44585));
    InMux I__8203 (
            .O(N__44588),
            .I(N__44582));
    LocalMux I__8202 (
            .O(N__44585),
            .I(N__44577));
    LocalMux I__8201 (
            .O(N__44582),
            .I(N__44577));
    Span4Mux_v I__8200 (
            .O(N__44577),
            .I(N__44574));
    Span4Mux_v I__8199 (
            .O(N__44574),
            .I(N__44571));
    Span4Mux_v I__8198 (
            .O(N__44571),
            .I(N__44568));
    Odrv4 I__8197 (
            .O(N__44568),
            .I(n17571));
    InMux I__8196 (
            .O(N__44565),
            .I(N__44562));
    LocalMux I__8195 (
            .O(N__44562),
            .I(N__44559));
    Span4Mux_h I__8194 (
            .O(N__44559),
            .I(N__44554));
    InMux I__8193 (
            .O(N__44558),
            .I(N__44549));
    InMux I__8192 (
            .O(N__44557),
            .I(N__44549));
    Sp12to4 I__8191 (
            .O(N__44554),
            .I(N__44545));
    LocalMux I__8190 (
            .O(N__44549),
            .I(N__44542));
    InMux I__8189 (
            .O(N__44548),
            .I(N__44539));
    Span12Mux_v I__8188 (
            .O(N__44545),
            .I(N__44536));
    Span4Mux_h I__8187 (
            .O(N__44542),
            .I(N__44533));
    LocalMux I__8186 (
            .O(N__44539),
            .I(data_in_1_6));
    Odrv12 I__8185 (
            .O(N__44536),
            .I(data_in_1_6));
    Odrv4 I__8184 (
            .O(N__44533),
            .I(data_in_1_6));
    InMux I__8183 (
            .O(N__44526),
            .I(N__44522));
    InMux I__8182 (
            .O(N__44525),
            .I(N__44519));
    LocalMux I__8181 (
            .O(N__44522),
            .I(N__44514));
    LocalMux I__8180 (
            .O(N__44519),
            .I(N__44514));
    Span4Mux_v I__8179 (
            .O(N__44514),
            .I(N__44510));
    InMux I__8178 (
            .O(N__44513),
            .I(N__44507));
    Span4Mux_v I__8177 (
            .O(N__44510),
            .I(N__44504));
    LocalMux I__8176 (
            .O(N__44507),
            .I(data_in_0_6));
    Odrv4 I__8175 (
            .O(N__44504),
            .I(data_in_0_6));
    InMux I__8174 (
            .O(N__44499),
            .I(N__44496));
    LocalMux I__8173 (
            .O(N__44496),
            .I(N__44493));
    Span4Mux_v I__8172 (
            .O(N__44493),
            .I(N__44489));
    CascadeMux I__8171 (
            .O(N__44492),
            .I(N__44486));
    Span4Mux_h I__8170 (
            .O(N__44489),
            .I(N__44482));
    InMux I__8169 (
            .O(N__44486),
            .I(N__44479));
    CascadeMux I__8168 (
            .O(N__44485),
            .I(N__44476));
    Sp12to4 I__8167 (
            .O(N__44482),
            .I(N__44473));
    LocalMux I__8166 (
            .O(N__44479),
            .I(N__44470));
    InMux I__8165 (
            .O(N__44476),
            .I(N__44467));
    Span12Mux_h I__8164 (
            .O(N__44473),
            .I(N__44459));
    Sp12to4 I__8163 (
            .O(N__44470),
            .I(N__44459));
    LocalMux I__8162 (
            .O(N__44467),
            .I(N__44459));
    InMux I__8161 (
            .O(N__44466),
            .I(N__44456));
    Span12Mux_v I__8160 (
            .O(N__44459),
            .I(N__44453));
    LocalMux I__8159 (
            .O(N__44456),
            .I(data_in_3_6));
    Odrv12 I__8158 (
            .O(N__44453),
            .I(data_in_3_6));
    CascadeMux I__8157 (
            .O(N__44448),
            .I(N__44445));
    InMux I__8156 (
            .O(N__44445),
            .I(N__44442));
    LocalMux I__8155 (
            .O(N__44442),
            .I(\c0.n20_adj_4726 ));
    InMux I__8154 (
            .O(N__44439),
            .I(N__44436));
    LocalMux I__8153 (
            .O(N__44436),
            .I(\c0.n27_adj_4735 ));
    InMux I__8152 (
            .O(N__44433),
            .I(N__44429));
    CascadeMux I__8151 (
            .O(N__44432),
            .I(N__44426));
    LocalMux I__8150 (
            .O(N__44429),
            .I(N__44423));
    InMux I__8149 (
            .O(N__44426),
            .I(N__44420));
    Span4Mux_v I__8148 (
            .O(N__44423),
            .I(N__44417));
    LocalMux I__8147 (
            .O(N__44420),
            .I(N__44414));
    Odrv4 I__8146 (
            .O(N__44417),
            .I(\c0.data_out_frame_29__7__N_735 ));
    Odrv12 I__8145 (
            .O(N__44414),
            .I(\c0.data_out_frame_29__7__N_735 ));
    InMux I__8144 (
            .O(N__44409),
            .I(N__44406));
    LocalMux I__8143 (
            .O(N__44406),
            .I(N__44402));
    InMux I__8142 (
            .O(N__44405),
            .I(N__44399));
    Span4Mux_h I__8141 (
            .O(N__44402),
            .I(N__44396));
    LocalMux I__8140 (
            .O(N__44399),
            .I(N__44393));
    Span4Mux_v I__8139 (
            .O(N__44396),
            .I(N__44390));
    Span4Mux_v I__8138 (
            .O(N__44393),
            .I(N__44387));
    Odrv4 I__8137 (
            .O(N__44390),
            .I(\c0.n13665 ));
    Odrv4 I__8136 (
            .O(N__44387),
            .I(\c0.n13665 ));
    InMux I__8135 (
            .O(N__44382),
            .I(N__44379));
    LocalMux I__8134 (
            .O(N__44379),
            .I(N__44376));
    Span4Mux_h I__8133 (
            .O(N__44376),
            .I(N__44373));
    Odrv4 I__8132 (
            .O(N__44373),
            .I(\c0.n22754 ));
    InMux I__8131 (
            .O(N__44370),
            .I(N__44367));
    LocalMux I__8130 (
            .O(N__44367),
            .I(N__44364));
    Span4Mux_h I__8129 (
            .O(N__44364),
            .I(N__44360));
    InMux I__8128 (
            .O(N__44363),
            .I(N__44357));
    Odrv4 I__8127 (
            .O(N__44360),
            .I(\c0.n13558 ));
    LocalMux I__8126 (
            .O(N__44357),
            .I(\c0.n13558 ));
    CascadeMux I__8125 (
            .O(N__44352),
            .I(\c0.n22754_cascade_ ));
    InMux I__8124 (
            .O(N__44349),
            .I(N__44346));
    LocalMux I__8123 (
            .O(N__44346),
            .I(N__44342));
    InMux I__8122 (
            .O(N__44345),
            .I(N__44339));
    Span4Mux_v I__8121 (
            .O(N__44342),
            .I(N__44336));
    LocalMux I__8120 (
            .O(N__44339),
            .I(\c0.n22243 ));
    Odrv4 I__8119 (
            .O(N__44336),
            .I(\c0.n22243 ));
    CascadeMux I__8118 (
            .O(N__44331),
            .I(N__44328));
    InMux I__8117 (
            .O(N__44328),
            .I(N__44322));
    InMux I__8116 (
            .O(N__44327),
            .I(N__44315));
    InMux I__8115 (
            .O(N__44326),
            .I(N__44315));
    InMux I__8114 (
            .O(N__44325),
            .I(N__44315));
    LocalMux I__8113 (
            .O(N__44322),
            .I(N__44311));
    LocalMux I__8112 (
            .O(N__44315),
            .I(N__44308));
    InMux I__8111 (
            .O(N__44314),
            .I(N__44305));
    Span4Mux_h I__8110 (
            .O(N__44311),
            .I(N__44302));
    Span4Mux_v I__8109 (
            .O(N__44308),
            .I(N__44299));
    LocalMux I__8108 (
            .O(N__44305),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv4 I__8107 (
            .O(N__44302),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv4 I__8106 (
            .O(N__44299),
            .I(\c0.FRAME_MATCHER_state_20 ));
    SRMux I__8105 (
            .O(N__44292),
            .I(N__44289));
    LocalMux I__8104 (
            .O(N__44289),
            .I(N__44286));
    Span4Mux_h I__8103 (
            .O(N__44286),
            .I(N__44283));
    Span4Mux_v I__8102 (
            .O(N__44283),
            .I(N__44280));
    Odrv4 I__8101 (
            .O(N__44280),
            .I(\c0.n8_adj_4553 ));
    InMux I__8100 (
            .O(N__44277),
            .I(N__44273));
    InMux I__8099 (
            .O(N__44276),
            .I(N__44270));
    LocalMux I__8098 (
            .O(N__44273),
            .I(N__44266));
    LocalMux I__8097 (
            .O(N__44270),
            .I(N__44263));
    InMux I__8096 (
            .O(N__44269),
            .I(N__44259));
    Span4Mux_h I__8095 (
            .O(N__44266),
            .I(N__44256));
    Span4Mux_v I__8094 (
            .O(N__44263),
            .I(N__44253));
    InMux I__8093 (
            .O(N__44262),
            .I(N__44250));
    LocalMux I__8092 (
            .O(N__44259),
            .I(N__44247));
    Odrv4 I__8091 (
            .O(N__44256),
            .I(\c0.n4_adj_4212 ));
    Odrv4 I__8090 (
            .O(N__44253),
            .I(\c0.n4_adj_4212 ));
    LocalMux I__8089 (
            .O(N__44250),
            .I(\c0.n4_adj_4212 ));
    Odrv12 I__8088 (
            .O(N__44247),
            .I(\c0.n4_adj_4212 ));
    CascadeMux I__8087 (
            .O(N__44238),
            .I(\c0.n22098_cascade_ ));
    InMux I__8086 (
            .O(N__44235),
            .I(N__44232));
    LocalMux I__8085 (
            .O(N__44232),
            .I(\c0.n4_adj_4306 ));
    CascadeMux I__8084 (
            .O(N__44229),
            .I(\c0.n63_adj_4305_cascade_ ));
    CascadeMux I__8083 (
            .O(N__44226),
            .I(N__44222));
    InMux I__8082 (
            .O(N__44225),
            .I(N__44214));
    InMux I__8081 (
            .O(N__44222),
            .I(N__44205));
    InMux I__8080 (
            .O(N__44221),
            .I(N__44205));
    InMux I__8079 (
            .O(N__44220),
            .I(N__44205));
    InMux I__8078 (
            .O(N__44219),
            .I(N__44205));
    CascadeMux I__8077 (
            .O(N__44218),
            .I(N__44202));
    CascadeMux I__8076 (
            .O(N__44217),
            .I(N__44198));
    LocalMux I__8075 (
            .O(N__44214),
            .I(N__44191));
    LocalMux I__8074 (
            .O(N__44205),
            .I(N__44188));
    InMux I__8073 (
            .O(N__44202),
            .I(N__44179));
    InMux I__8072 (
            .O(N__44201),
            .I(N__44179));
    InMux I__8071 (
            .O(N__44198),
            .I(N__44179));
    InMux I__8070 (
            .O(N__44197),
            .I(N__44179));
    InMux I__8069 (
            .O(N__44196),
            .I(N__44176));
    InMux I__8068 (
            .O(N__44195),
            .I(N__44173));
    InMux I__8067 (
            .O(N__44194),
            .I(N__44170));
    Span4Mux_v I__8066 (
            .O(N__44191),
            .I(N__44159));
    Span4Mux_h I__8065 (
            .O(N__44188),
            .I(N__44159));
    LocalMux I__8064 (
            .O(N__44179),
            .I(N__44159));
    LocalMux I__8063 (
            .O(N__44176),
            .I(N__44159));
    LocalMux I__8062 (
            .O(N__44173),
            .I(N__44159));
    LocalMux I__8061 (
            .O(N__44170),
            .I(N__44155));
    Span4Mux_h I__8060 (
            .O(N__44159),
            .I(N__44152));
    InMux I__8059 (
            .O(N__44158),
            .I(N__44149));
    Odrv4 I__8058 (
            .O(N__44155),
            .I(\c0.n13001 ));
    Odrv4 I__8057 (
            .O(N__44152),
            .I(\c0.n13001 ));
    LocalMux I__8056 (
            .O(N__44149),
            .I(\c0.n13001 ));
    CascadeMux I__8055 (
            .O(N__44142),
            .I(N__44138));
    InMux I__8054 (
            .O(N__44141),
            .I(N__44135));
    InMux I__8053 (
            .O(N__44138),
            .I(N__44132));
    LocalMux I__8052 (
            .O(N__44135),
            .I(N__44128));
    LocalMux I__8051 (
            .O(N__44132),
            .I(N__44125));
    InMux I__8050 (
            .O(N__44131),
            .I(N__44122));
    Span4Mux_h I__8049 (
            .O(N__44128),
            .I(N__44119));
    Span4Mux_h I__8048 (
            .O(N__44125),
            .I(N__44116));
    LocalMux I__8047 (
            .O(N__44122),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__8046 (
            .O(N__44119),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__8045 (
            .O(N__44116),
            .I(\c0.FRAME_MATCHER_state_0 ));
    InMux I__8044 (
            .O(N__44109),
            .I(N__44105));
    InMux I__8043 (
            .O(N__44108),
            .I(N__44100));
    LocalMux I__8042 (
            .O(N__44105),
            .I(N__44097));
    InMux I__8041 (
            .O(N__44104),
            .I(N__44094));
    InMux I__8040 (
            .O(N__44103),
            .I(N__44091));
    LocalMux I__8039 (
            .O(N__44100),
            .I(N__44088));
    Span4Mux_v I__8038 (
            .O(N__44097),
            .I(N__44079));
    LocalMux I__8037 (
            .O(N__44094),
            .I(N__44079));
    LocalMux I__8036 (
            .O(N__44091),
            .I(N__44079));
    Span4Mux_h I__8035 (
            .O(N__44088),
            .I(N__44076));
    InMux I__8034 (
            .O(N__44087),
            .I(N__44073));
    InMux I__8033 (
            .O(N__44086),
            .I(N__44070));
    Span4Mux_h I__8032 (
            .O(N__44079),
            .I(N__44067));
    Odrv4 I__8031 (
            .O(N__44076),
            .I(\c0.n9248 ));
    LocalMux I__8030 (
            .O(N__44073),
            .I(\c0.n9248 ));
    LocalMux I__8029 (
            .O(N__44070),
            .I(\c0.n9248 ));
    Odrv4 I__8028 (
            .O(N__44067),
            .I(\c0.n9248 ));
    InMux I__8027 (
            .O(N__44058),
            .I(N__44053));
    InMux I__8026 (
            .O(N__44057),
            .I(N__44050));
    InMux I__8025 (
            .O(N__44056),
            .I(N__44047));
    LocalMux I__8024 (
            .O(N__44053),
            .I(N__44040));
    LocalMux I__8023 (
            .O(N__44050),
            .I(N__44040));
    LocalMux I__8022 (
            .O(N__44047),
            .I(N__44037));
    InMux I__8021 (
            .O(N__44046),
            .I(N__44034));
    InMux I__8020 (
            .O(N__44045),
            .I(N__44031));
    Span4Mux_h I__8019 (
            .O(N__44040),
            .I(N__44028));
    Span4Mux_h I__8018 (
            .O(N__44037),
            .I(N__44025));
    LocalMux I__8017 (
            .O(N__44034),
            .I(N__44022));
    LocalMux I__8016 (
            .O(N__44031),
            .I(\c0.n13055 ));
    Odrv4 I__8015 (
            .O(N__44028),
            .I(\c0.n13055 ));
    Odrv4 I__8014 (
            .O(N__44025),
            .I(\c0.n13055 ));
    Odrv4 I__8013 (
            .O(N__44022),
            .I(\c0.n13055 ));
    InMux I__8012 (
            .O(N__44013),
            .I(N__44008));
    CascadeMux I__8011 (
            .O(N__44012),
            .I(N__44005));
    CascadeMux I__8010 (
            .O(N__44011),
            .I(N__43999));
    LocalMux I__8009 (
            .O(N__44008),
            .I(N__43994));
    InMux I__8008 (
            .O(N__44005),
            .I(N__43991));
    InMux I__8007 (
            .O(N__44004),
            .I(N__43986));
    InMux I__8006 (
            .O(N__44003),
            .I(N__43986));
    InMux I__8005 (
            .O(N__44002),
            .I(N__43983));
    InMux I__8004 (
            .O(N__43999),
            .I(N__43980));
    InMux I__8003 (
            .O(N__43998),
            .I(N__43977));
    CascadeMux I__8002 (
            .O(N__43997),
            .I(N__43974));
    Span4Mux_v I__8001 (
            .O(N__43994),
            .I(N__43969));
    LocalMux I__8000 (
            .O(N__43991),
            .I(N__43969));
    LocalMux I__7999 (
            .O(N__43986),
            .I(N__43964));
    LocalMux I__7998 (
            .O(N__43983),
            .I(N__43959));
    LocalMux I__7997 (
            .O(N__43980),
            .I(N__43959));
    LocalMux I__7996 (
            .O(N__43977),
            .I(N__43956));
    InMux I__7995 (
            .O(N__43974),
            .I(N__43953));
    Span4Mux_h I__7994 (
            .O(N__43969),
            .I(N__43950));
    InMux I__7993 (
            .O(N__43968),
            .I(N__43947));
    InMux I__7992 (
            .O(N__43967),
            .I(N__43944));
    Span4Mux_v I__7991 (
            .O(N__43964),
            .I(N__43939));
    Span4Mux_v I__7990 (
            .O(N__43959),
            .I(N__43939));
    Odrv4 I__7989 (
            .O(N__43956),
            .I(\c0.data_out_frame_29_7_N_1482_0 ));
    LocalMux I__7988 (
            .O(N__43953),
            .I(\c0.data_out_frame_29_7_N_1482_0 ));
    Odrv4 I__7987 (
            .O(N__43950),
            .I(\c0.data_out_frame_29_7_N_1482_0 ));
    LocalMux I__7986 (
            .O(N__43947),
            .I(\c0.data_out_frame_29_7_N_1482_0 ));
    LocalMux I__7985 (
            .O(N__43944),
            .I(\c0.data_out_frame_29_7_N_1482_0 ));
    Odrv4 I__7984 (
            .O(N__43939),
            .I(\c0.data_out_frame_29_7_N_1482_0 ));
    InMux I__7983 (
            .O(N__43926),
            .I(N__43918));
    InMux I__7982 (
            .O(N__43925),
            .I(N__43918));
    InMux I__7981 (
            .O(N__43924),
            .I(N__43915));
    InMux I__7980 (
            .O(N__43923),
            .I(N__43912));
    LocalMux I__7979 (
            .O(N__43918),
            .I(N__43908));
    LocalMux I__7978 (
            .O(N__43915),
            .I(N__43905));
    LocalMux I__7977 (
            .O(N__43912),
            .I(N__43902));
    InMux I__7976 (
            .O(N__43911),
            .I(N__43896));
    Span4Mux_h I__7975 (
            .O(N__43908),
            .I(N__43891));
    Span4Mux_v I__7974 (
            .O(N__43905),
            .I(N__43891));
    Span4Mux_h I__7973 (
            .O(N__43902),
            .I(N__43888));
    InMux I__7972 (
            .O(N__43901),
            .I(N__43885));
    InMux I__7971 (
            .O(N__43900),
            .I(N__43880));
    InMux I__7970 (
            .O(N__43899),
            .I(N__43880));
    LocalMux I__7969 (
            .O(N__43896),
            .I(data_out_frame_29_7_N_2878_2));
    Odrv4 I__7968 (
            .O(N__43891),
            .I(data_out_frame_29_7_N_2878_2));
    Odrv4 I__7967 (
            .O(N__43888),
            .I(data_out_frame_29_7_N_2878_2));
    LocalMux I__7966 (
            .O(N__43885),
            .I(data_out_frame_29_7_N_2878_2));
    LocalMux I__7965 (
            .O(N__43880),
            .I(data_out_frame_29_7_N_2878_2));
    InMux I__7964 (
            .O(N__43869),
            .I(N__43866));
    LocalMux I__7963 (
            .O(N__43866),
            .I(N__43862));
    InMux I__7962 (
            .O(N__43865),
            .I(N__43859));
    Span4Mux_h I__7961 (
            .O(N__43862),
            .I(N__43856));
    LocalMux I__7960 (
            .O(N__43859),
            .I(N__43853));
    Span4Mux_h I__7959 (
            .O(N__43856),
            .I(N__43850));
    Span4Mux_v I__7958 (
            .O(N__43853),
            .I(N__43847));
    Odrv4 I__7957 (
            .O(N__43850),
            .I(\c0.n9_adj_4549 ));
    Odrv4 I__7956 (
            .O(N__43847),
            .I(\c0.n9_adj_4549 ));
    CascadeMux I__7955 (
            .O(N__43842),
            .I(N__43839));
    InMux I__7954 (
            .O(N__43839),
            .I(N__43831));
    CascadeMux I__7953 (
            .O(N__43838),
            .I(N__43826));
    InMux I__7952 (
            .O(N__43837),
            .I(N__43821));
    InMux I__7951 (
            .O(N__43836),
            .I(N__43817));
    CascadeMux I__7950 (
            .O(N__43835),
            .I(N__43813));
    CascadeMux I__7949 (
            .O(N__43834),
            .I(N__43810));
    LocalMux I__7948 (
            .O(N__43831),
            .I(N__43806));
    InMux I__7947 (
            .O(N__43830),
            .I(N__43803));
    InMux I__7946 (
            .O(N__43829),
            .I(N__43800));
    InMux I__7945 (
            .O(N__43826),
            .I(N__43797));
    InMux I__7944 (
            .O(N__43825),
            .I(N__43793));
    InMux I__7943 (
            .O(N__43824),
            .I(N__43790));
    LocalMux I__7942 (
            .O(N__43821),
            .I(N__43787));
    InMux I__7941 (
            .O(N__43820),
            .I(N__43784));
    LocalMux I__7940 (
            .O(N__43817),
            .I(N__43781));
    InMux I__7939 (
            .O(N__43816),
            .I(N__43778));
    InMux I__7938 (
            .O(N__43813),
            .I(N__43773));
    InMux I__7937 (
            .O(N__43810),
            .I(N__43773));
    InMux I__7936 (
            .O(N__43809),
            .I(N__43770));
    Span4Mux_v I__7935 (
            .O(N__43806),
            .I(N__43765));
    LocalMux I__7934 (
            .O(N__43803),
            .I(N__43765));
    LocalMux I__7933 (
            .O(N__43800),
            .I(N__43760));
    LocalMux I__7932 (
            .O(N__43797),
            .I(N__43760));
    InMux I__7931 (
            .O(N__43796),
            .I(N__43757));
    LocalMux I__7930 (
            .O(N__43793),
            .I(N__43754));
    LocalMux I__7929 (
            .O(N__43790),
            .I(N__43737));
    Span4Mux_h I__7928 (
            .O(N__43787),
            .I(N__43737));
    LocalMux I__7927 (
            .O(N__43784),
            .I(N__43737));
    Span4Mux_v I__7926 (
            .O(N__43781),
            .I(N__43737));
    LocalMux I__7925 (
            .O(N__43778),
            .I(N__43737));
    LocalMux I__7924 (
            .O(N__43773),
            .I(N__43737));
    LocalMux I__7923 (
            .O(N__43770),
            .I(N__43737));
    Span4Mux_h I__7922 (
            .O(N__43765),
            .I(N__43734));
    Span4Mux_h I__7921 (
            .O(N__43760),
            .I(N__43727));
    LocalMux I__7920 (
            .O(N__43757),
            .I(N__43727));
    Span4Mux_v I__7919 (
            .O(N__43754),
            .I(N__43727));
    InMux I__7918 (
            .O(N__43753),
            .I(N__43722));
    InMux I__7917 (
            .O(N__43752),
            .I(N__43722));
    Span4Mux_v I__7916 (
            .O(N__43737),
            .I(N__43719));
    Odrv4 I__7915 (
            .O(N__43734),
            .I(n63));
    Odrv4 I__7914 (
            .O(N__43727),
            .I(n63));
    LocalMux I__7913 (
            .O(N__43722),
            .I(n63));
    Odrv4 I__7912 (
            .O(N__43719),
            .I(n63));
    InMux I__7911 (
            .O(N__43710),
            .I(N__43705));
    InMux I__7910 (
            .O(N__43709),
            .I(N__43702));
    CascadeMux I__7909 (
            .O(N__43708),
            .I(N__43699));
    LocalMux I__7908 (
            .O(N__43705),
            .I(N__43693));
    LocalMux I__7907 (
            .O(N__43702),
            .I(N__43693));
    InMux I__7906 (
            .O(N__43699),
            .I(N__43690));
    InMux I__7905 (
            .O(N__43698),
            .I(N__43687));
    Span4Mux_v I__7904 (
            .O(N__43693),
            .I(N__43682));
    LocalMux I__7903 (
            .O(N__43690),
            .I(N__43682));
    LocalMux I__7902 (
            .O(N__43687),
            .I(N__43679));
    Span4Mux_h I__7901 (
            .O(N__43682),
            .I(N__43676));
    Odrv4 I__7900 (
            .O(N__43679),
            .I(\c0.n3844 ));
    Odrv4 I__7899 (
            .O(N__43676),
            .I(\c0.n3844 ));
    InMux I__7898 (
            .O(N__43671),
            .I(N__43668));
    LocalMux I__7897 (
            .O(N__43668),
            .I(N__43664));
    InMux I__7896 (
            .O(N__43667),
            .I(N__43661));
    Span4Mux_v I__7895 (
            .O(N__43664),
            .I(N__43656));
    LocalMux I__7894 (
            .O(N__43661),
            .I(N__43656));
    Span4Mux_h I__7893 (
            .O(N__43656),
            .I(N__43651));
    InMux I__7892 (
            .O(N__43655),
            .I(N__43648));
    InMux I__7891 (
            .O(N__43654),
            .I(N__43645));
    Odrv4 I__7890 (
            .O(N__43651),
            .I(\c0.n58_adj_4706 ));
    LocalMux I__7889 (
            .O(N__43648),
            .I(\c0.n58_adj_4706 ));
    LocalMux I__7888 (
            .O(N__43645),
            .I(\c0.n58_adj_4706 ));
    CascadeMux I__7887 (
            .O(N__43638),
            .I(\c0.n24591_cascade_ ));
    InMux I__7886 (
            .O(N__43635),
            .I(N__43632));
    LocalMux I__7885 (
            .O(N__43632),
            .I(N__43629));
    Span4Mux_h I__7884 (
            .O(N__43629),
            .I(N__43626));
    Odrv4 I__7883 (
            .O(N__43626),
            .I(\c0.n6_adj_4728 ));
    InMux I__7882 (
            .O(N__43623),
            .I(N__43620));
    LocalMux I__7881 (
            .O(N__43620),
            .I(N__43617));
    Span12Mux_v I__7880 (
            .O(N__43617),
            .I(N__43614));
    Odrv12 I__7879 (
            .O(N__43614),
            .I(\c0.FRAME_MATCHER_state_2 ));
    InMux I__7878 (
            .O(N__43611),
            .I(N__43606));
    InMux I__7877 (
            .O(N__43610),
            .I(N__43599));
    InMux I__7876 (
            .O(N__43609),
            .I(N__43599));
    LocalMux I__7875 (
            .O(N__43606),
            .I(N__43595));
    InMux I__7874 (
            .O(N__43605),
            .I(N__43592));
    InMux I__7873 (
            .O(N__43604),
            .I(N__43589));
    LocalMux I__7872 (
            .O(N__43599),
            .I(N__43586));
    InMux I__7871 (
            .O(N__43598),
            .I(N__43583));
    Span4Mux_h I__7870 (
            .O(N__43595),
            .I(N__43580));
    LocalMux I__7869 (
            .O(N__43592),
            .I(N__43575));
    LocalMux I__7868 (
            .O(N__43589),
            .I(N__43575));
    Span4Mux_h I__7867 (
            .O(N__43586),
            .I(N__43572));
    LocalMux I__7866 (
            .O(N__43583),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__7865 (
            .O(N__43580),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__7864 (
            .O(N__43575),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__7863 (
            .O(N__43572),
            .I(\c0.FRAME_MATCHER_state_15 ));
    SRMux I__7862 (
            .O(N__43563),
            .I(N__43560));
    LocalMux I__7861 (
            .O(N__43560),
            .I(N__43557));
    Span12Mux_s9_v I__7860 (
            .O(N__43557),
            .I(N__43554));
    Odrv12 I__7859 (
            .O(N__43554),
            .I(\c0.n21659 ));
    InMux I__7858 (
            .O(N__43551),
            .I(N__43548));
    LocalMux I__7857 (
            .O(N__43548),
            .I(\c0.n4_adj_4721 ));
    CascadeMux I__7856 (
            .O(N__43545),
            .I(N__43542));
    InMux I__7855 (
            .O(N__43542),
            .I(N__43539));
    LocalMux I__7854 (
            .O(N__43539),
            .I(N__43536));
    Odrv12 I__7853 (
            .O(N__43536),
            .I(\c0.n937 ));
    InMux I__7852 (
            .O(N__43533),
            .I(N__43527));
    InMux I__7851 (
            .O(N__43532),
            .I(N__43523));
    InMux I__7850 (
            .O(N__43531),
            .I(N__43520));
    InMux I__7849 (
            .O(N__43530),
            .I(N__43517));
    LocalMux I__7848 (
            .O(N__43527),
            .I(N__43510));
    InMux I__7847 (
            .O(N__43526),
            .I(N__43507));
    LocalMux I__7846 (
            .O(N__43523),
            .I(N__43500));
    LocalMux I__7845 (
            .O(N__43520),
            .I(N__43500));
    LocalMux I__7844 (
            .O(N__43517),
            .I(N__43500));
    InMux I__7843 (
            .O(N__43516),
            .I(N__43497));
    InMux I__7842 (
            .O(N__43515),
            .I(N__43494));
    InMux I__7841 (
            .O(N__43514),
            .I(N__43488));
    InMux I__7840 (
            .O(N__43513),
            .I(N__43485));
    Span4Mux_v I__7839 (
            .O(N__43510),
            .I(N__43478));
    LocalMux I__7838 (
            .O(N__43507),
            .I(N__43478));
    Span4Mux_v I__7837 (
            .O(N__43500),
            .I(N__43478));
    LocalMux I__7836 (
            .O(N__43497),
            .I(N__43473));
    LocalMux I__7835 (
            .O(N__43494),
            .I(N__43473));
    InMux I__7834 (
            .O(N__43493),
            .I(N__43468));
    InMux I__7833 (
            .O(N__43492),
            .I(N__43468));
    InMux I__7832 (
            .O(N__43491),
            .I(N__43465));
    LocalMux I__7831 (
            .O(N__43488),
            .I(\c0.data_out_frame_29_7_N_1482_1 ));
    LocalMux I__7830 (
            .O(N__43485),
            .I(\c0.data_out_frame_29_7_N_1482_1 ));
    Odrv4 I__7829 (
            .O(N__43478),
            .I(\c0.data_out_frame_29_7_N_1482_1 ));
    Odrv4 I__7828 (
            .O(N__43473),
            .I(\c0.data_out_frame_29_7_N_1482_1 ));
    LocalMux I__7827 (
            .O(N__43468),
            .I(\c0.data_out_frame_29_7_N_1482_1 ));
    LocalMux I__7826 (
            .O(N__43465),
            .I(\c0.data_out_frame_29_7_N_1482_1 ));
    CascadeMux I__7825 (
            .O(N__43452),
            .I(N__43449));
    InMux I__7824 (
            .O(N__43449),
            .I(N__43446));
    LocalMux I__7823 (
            .O(N__43446),
            .I(N__43442));
    InMux I__7822 (
            .O(N__43445),
            .I(N__43439));
    Span4Mux_h I__7821 (
            .O(N__43442),
            .I(N__43436));
    LocalMux I__7820 (
            .O(N__43439),
            .I(\c0.FRAME_MATCHER_state_1 ));
    Odrv4 I__7819 (
            .O(N__43436),
            .I(\c0.FRAME_MATCHER_state_1 ));
    CascadeMux I__7818 (
            .O(N__43431),
            .I(N__43428));
    InMux I__7817 (
            .O(N__43428),
            .I(N__43425));
    LocalMux I__7816 (
            .O(N__43425),
            .I(N__43422));
    Span4Mux_h I__7815 (
            .O(N__43422),
            .I(N__43419));
    Odrv4 I__7814 (
            .O(N__43419),
            .I(\c0.n74_adj_4525 ));
    InMux I__7813 (
            .O(N__43416),
            .I(N__43412));
    InMux I__7812 (
            .O(N__43415),
            .I(N__43409));
    LocalMux I__7811 (
            .O(N__43412),
            .I(N__43403));
    LocalMux I__7810 (
            .O(N__43409),
            .I(N__43403));
    InMux I__7809 (
            .O(N__43408),
            .I(N__43400));
    Span4Mux_h I__7808 (
            .O(N__43403),
            .I(N__43397));
    LocalMux I__7807 (
            .O(N__43400),
            .I(N__43390));
    Span4Mux_v I__7806 (
            .O(N__43397),
            .I(N__43390));
    InMux I__7805 (
            .O(N__43396),
            .I(N__43387));
    InMux I__7804 (
            .O(N__43395),
            .I(N__43384));
    Span4Mux_v I__7803 (
            .O(N__43390),
            .I(N__43381));
    LocalMux I__7802 (
            .O(N__43387),
            .I(N__43378));
    LocalMux I__7801 (
            .O(N__43384),
            .I(control_mode_6));
    Odrv4 I__7800 (
            .O(N__43381),
            .I(control_mode_6));
    Odrv4 I__7799 (
            .O(N__43378),
            .I(control_mode_6));
    InMux I__7798 (
            .O(N__43371),
            .I(N__43368));
    LocalMux I__7797 (
            .O(N__43368),
            .I(N__43364));
    InMux I__7796 (
            .O(N__43367),
            .I(N__43360));
    Span4Mux_v I__7795 (
            .O(N__43364),
            .I(N__43357));
    InMux I__7794 (
            .O(N__43363),
            .I(N__43354));
    LocalMux I__7793 (
            .O(N__43360),
            .I(data_in_1_1));
    Odrv4 I__7792 (
            .O(N__43357),
            .I(data_in_1_1));
    LocalMux I__7791 (
            .O(N__43354),
            .I(data_in_1_1));
    InMux I__7790 (
            .O(N__43347),
            .I(N__43342));
    InMux I__7789 (
            .O(N__43346),
            .I(N__43339));
    InMux I__7788 (
            .O(N__43345),
            .I(N__43336));
    LocalMux I__7787 (
            .O(N__43342),
            .I(data_in_0_1));
    LocalMux I__7786 (
            .O(N__43339),
            .I(data_in_0_1));
    LocalMux I__7785 (
            .O(N__43336),
            .I(data_in_0_1));
    InMux I__7784 (
            .O(N__43329),
            .I(N__43325));
    CascadeMux I__7783 (
            .O(N__43328),
            .I(N__43322));
    LocalMux I__7782 (
            .O(N__43325),
            .I(N__43319));
    InMux I__7781 (
            .O(N__43322),
            .I(N__43314));
    Span4Mux_h I__7780 (
            .O(N__43319),
            .I(N__43311));
    InMux I__7779 (
            .O(N__43318),
            .I(N__43308));
    InMux I__7778 (
            .O(N__43317),
            .I(N__43305));
    LocalMux I__7777 (
            .O(N__43314),
            .I(data_in_3_2));
    Odrv4 I__7776 (
            .O(N__43311),
            .I(data_in_3_2));
    LocalMux I__7775 (
            .O(N__43308),
            .I(data_in_3_2));
    LocalMux I__7774 (
            .O(N__43305),
            .I(data_in_3_2));
    CascadeMux I__7773 (
            .O(N__43296),
            .I(N__43293));
    InMux I__7772 (
            .O(N__43293),
            .I(N__43289));
    InMux I__7771 (
            .O(N__43292),
            .I(N__43286));
    LocalMux I__7770 (
            .O(N__43289),
            .I(N__43282));
    LocalMux I__7769 (
            .O(N__43286),
            .I(N__43279));
    InMux I__7768 (
            .O(N__43285),
            .I(N__43276));
    Span4Mux_v I__7767 (
            .O(N__43282),
            .I(N__43271));
    Span4Mux_v I__7766 (
            .O(N__43279),
            .I(N__43268));
    LocalMux I__7765 (
            .O(N__43276),
            .I(N__43265));
    InMux I__7764 (
            .O(N__43275),
            .I(N__43262));
    InMux I__7763 (
            .O(N__43274),
            .I(N__43259));
    Span4Mux_v I__7762 (
            .O(N__43271),
            .I(N__43256));
    Span4Mux_h I__7761 (
            .O(N__43268),
            .I(N__43253));
    Span12Mux_h I__7760 (
            .O(N__43265),
            .I(N__43248));
    LocalMux I__7759 (
            .O(N__43262),
            .I(N__43248));
    LocalMux I__7758 (
            .O(N__43259),
            .I(control_mode_4));
    Odrv4 I__7757 (
            .O(N__43256),
            .I(control_mode_4));
    Odrv4 I__7756 (
            .O(N__43253),
            .I(control_mode_4));
    Odrv12 I__7755 (
            .O(N__43248),
            .I(control_mode_4));
    InMux I__7754 (
            .O(N__43239),
            .I(N__43235));
    InMux I__7753 (
            .O(N__43238),
            .I(N__43224));
    LocalMux I__7752 (
            .O(N__43235),
            .I(N__43213));
    InMux I__7751 (
            .O(N__43234),
            .I(N__43210));
    InMux I__7750 (
            .O(N__43233),
            .I(N__43207));
    InMux I__7749 (
            .O(N__43232),
            .I(N__43193));
    InMux I__7748 (
            .O(N__43231),
            .I(N__43193));
    InMux I__7747 (
            .O(N__43230),
            .I(N__43193));
    InMux I__7746 (
            .O(N__43229),
            .I(N__43193));
    InMux I__7745 (
            .O(N__43228),
            .I(N__43193));
    InMux I__7744 (
            .O(N__43227),
            .I(N__43193));
    LocalMux I__7743 (
            .O(N__43224),
            .I(N__43190));
    InMux I__7742 (
            .O(N__43223),
            .I(N__43187));
    InMux I__7741 (
            .O(N__43222),
            .I(N__43183));
    InMux I__7740 (
            .O(N__43221),
            .I(N__43172));
    InMux I__7739 (
            .O(N__43220),
            .I(N__43168));
    InMux I__7738 (
            .O(N__43219),
            .I(N__43165));
    InMux I__7737 (
            .O(N__43218),
            .I(N__43161));
    InMux I__7736 (
            .O(N__43217),
            .I(N__43157));
    InMux I__7735 (
            .O(N__43216),
            .I(N__43154));
    Span4Mux_v I__7734 (
            .O(N__43213),
            .I(N__43149));
    LocalMux I__7733 (
            .O(N__43210),
            .I(N__43149));
    LocalMux I__7732 (
            .O(N__43207),
            .I(N__43146));
    InMux I__7731 (
            .O(N__43206),
            .I(N__43143));
    LocalMux I__7730 (
            .O(N__43193),
            .I(N__43138));
    Span4Mux_v I__7729 (
            .O(N__43190),
            .I(N__43138));
    LocalMux I__7728 (
            .O(N__43187),
            .I(N__43135));
    InMux I__7727 (
            .O(N__43186),
            .I(N__43132));
    LocalMux I__7726 (
            .O(N__43183),
            .I(N__43129));
    InMux I__7725 (
            .O(N__43182),
            .I(N__43126));
    InMux I__7724 (
            .O(N__43181),
            .I(N__43122));
    InMux I__7723 (
            .O(N__43180),
            .I(N__43119));
    InMux I__7722 (
            .O(N__43179),
            .I(N__43114));
    InMux I__7721 (
            .O(N__43178),
            .I(N__43114));
    InMux I__7720 (
            .O(N__43177),
            .I(N__43109));
    InMux I__7719 (
            .O(N__43176),
            .I(N__43109));
    InMux I__7718 (
            .O(N__43175),
            .I(N__43106));
    LocalMux I__7717 (
            .O(N__43172),
            .I(N__43103));
    InMux I__7716 (
            .O(N__43171),
            .I(N__43100));
    LocalMux I__7715 (
            .O(N__43168),
            .I(N__43097));
    LocalMux I__7714 (
            .O(N__43165),
            .I(N__43094));
    InMux I__7713 (
            .O(N__43164),
            .I(N__43091));
    LocalMux I__7712 (
            .O(N__43161),
            .I(N__43088));
    InMux I__7711 (
            .O(N__43160),
            .I(N__43081));
    LocalMux I__7710 (
            .O(N__43157),
            .I(N__43068));
    LocalMux I__7709 (
            .O(N__43154),
            .I(N__43068));
    Span4Mux_h I__7708 (
            .O(N__43149),
            .I(N__43068));
    Span4Mux_v I__7707 (
            .O(N__43146),
            .I(N__43068));
    LocalMux I__7706 (
            .O(N__43143),
            .I(N__43068));
    Span4Mux_v I__7705 (
            .O(N__43138),
            .I(N__43068));
    Span4Mux_v I__7704 (
            .O(N__43135),
            .I(N__43063));
    LocalMux I__7703 (
            .O(N__43132),
            .I(N__43063));
    Span4Mux_v I__7702 (
            .O(N__43129),
            .I(N__43055));
    LocalMux I__7701 (
            .O(N__43126),
            .I(N__43055));
    InMux I__7700 (
            .O(N__43125),
            .I(N__43050));
    LocalMux I__7699 (
            .O(N__43122),
            .I(N__43047));
    LocalMux I__7698 (
            .O(N__43119),
            .I(N__43044));
    LocalMux I__7697 (
            .O(N__43114),
            .I(N__43035));
    LocalMux I__7696 (
            .O(N__43109),
            .I(N__43035));
    LocalMux I__7695 (
            .O(N__43106),
            .I(N__43035));
    Span4Mux_h I__7694 (
            .O(N__43103),
            .I(N__43035));
    LocalMux I__7693 (
            .O(N__43100),
            .I(N__43029));
    Span4Mux_h I__7692 (
            .O(N__43097),
            .I(N__43024));
    Span4Mux_h I__7691 (
            .O(N__43094),
            .I(N__43024));
    LocalMux I__7690 (
            .O(N__43091),
            .I(N__43021));
    Span4Mux_v I__7689 (
            .O(N__43088),
            .I(N__43018));
    InMux I__7688 (
            .O(N__43087),
            .I(N__43009));
    InMux I__7687 (
            .O(N__43086),
            .I(N__43009));
    InMux I__7686 (
            .O(N__43085),
            .I(N__43009));
    InMux I__7685 (
            .O(N__43084),
            .I(N__43009));
    LocalMux I__7684 (
            .O(N__43081),
            .I(N__43006));
    Span4Mux_v I__7683 (
            .O(N__43068),
            .I(N__43001));
    Span4Mux_v I__7682 (
            .O(N__43063),
            .I(N__43001));
    InMux I__7681 (
            .O(N__43062),
            .I(N__42998));
    InMux I__7680 (
            .O(N__43061),
            .I(N__42993));
    InMux I__7679 (
            .O(N__43060),
            .I(N__42993));
    Sp12to4 I__7678 (
            .O(N__43055),
            .I(N__42990));
    InMux I__7677 (
            .O(N__43054),
            .I(N__42987));
    InMux I__7676 (
            .O(N__43053),
            .I(N__42984));
    LocalMux I__7675 (
            .O(N__43050),
            .I(N__42979));
    Span4Mux_h I__7674 (
            .O(N__43047),
            .I(N__42979));
    Span4Mux_h I__7673 (
            .O(N__43044),
            .I(N__42974));
    Span4Mux_h I__7672 (
            .O(N__43035),
            .I(N__42974));
    InMux I__7671 (
            .O(N__43034),
            .I(N__42967));
    InMux I__7670 (
            .O(N__43033),
            .I(N__42967));
    InMux I__7669 (
            .O(N__43032),
            .I(N__42967));
    Span4Mux_h I__7668 (
            .O(N__43029),
            .I(N__42960));
    Span4Mux_v I__7667 (
            .O(N__43024),
            .I(N__42960));
    Span4Mux_h I__7666 (
            .O(N__43021),
            .I(N__42960));
    Span4Mux_v I__7665 (
            .O(N__43018),
            .I(N__42953));
    LocalMux I__7664 (
            .O(N__43009),
            .I(N__42953));
    Span4Mux_v I__7663 (
            .O(N__43006),
            .I(N__42953));
    Sp12to4 I__7662 (
            .O(N__43001),
            .I(N__42948));
    LocalMux I__7661 (
            .O(N__42998),
            .I(N__42948));
    LocalMux I__7660 (
            .O(N__42993),
            .I(N__42943));
    Span12Mux_h I__7659 (
            .O(N__42990),
            .I(N__42943));
    LocalMux I__7658 (
            .O(N__42987),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__7657 (
            .O(N__42984),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7656 (
            .O(N__42979),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7655 (
            .O(N__42974),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__7654 (
            .O(N__42967),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7653 (
            .O(N__42960),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7652 (
            .O(N__42953),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__7651 (
            .O(N__42948),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__7650 (
            .O(N__42943),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__7649 (
            .O(N__42924),
            .I(N__42920));
    InMux I__7648 (
            .O(N__42923),
            .I(N__42917));
    LocalMux I__7647 (
            .O(N__42920),
            .I(N__42914));
    LocalMux I__7646 (
            .O(N__42917),
            .I(data_out_frame_9_4));
    Odrv12 I__7645 (
            .O(N__42914),
            .I(data_out_frame_9_4));
    InMux I__7644 (
            .O(N__42909),
            .I(N__42906));
    LocalMux I__7643 (
            .O(N__42906),
            .I(N__42902));
    InMux I__7642 (
            .O(N__42905),
            .I(N__42899));
    Span4Mux_v I__7641 (
            .O(N__42902),
            .I(N__42896));
    LocalMux I__7640 (
            .O(N__42899),
            .I(data_out_frame_8_4));
    Odrv4 I__7639 (
            .O(N__42896),
            .I(data_out_frame_8_4));
    InMux I__7638 (
            .O(N__42891),
            .I(N__42888));
    LocalMux I__7637 (
            .O(N__42888),
            .I(N__42885));
    Odrv4 I__7636 (
            .O(N__42885),
            .I(\c0.n24782 ));
    CascadeMux I__7635 (
            .O(N__42882),
            .I(N__42878));
    CascadeMux I__7634 (
            .O(N__42881),
            .I(N__42875));
    InMux I__7633 (
            .O(N__42878),
            .I(N__42872));
    InMux I__7632 (
            .O(N__42875),
            .I(N__42869));
    LocalMux I__7631 (
            .O(N__42872),
            .I(N__42866));
    LocalMux I__7630 (
            .O(N__42869),
            .I(N__42863));
    Span4Mux_v I__7629 (
            .O(N__42866),
            .I(N__42860));
    Span4Mux_v I__7628 (
            .O(N__42863),
            .I(N__42857));
    Span4Mux_h I__7627 (
            .O(N__42860),
            .I(N__42852));
    Span4Mux_v I__7626 (
            .O(N__42857),
            .I(N__42849));
    InMux I__7625 (
            .O(N__42856),
            .I(N__42846));
    InMux I__7624 (
            .O(N__42855),
            .I(N__42842));
    Sp12to4 I__7623 (
            .O(N__42852),
            .I(N__42839));
    Span4Mux_h I__7622 (
            .O(N__42849),
            .I(N__42834));
    LocalMux I__7621 (
            .O(N__42846),
            .I(N__42834));
    InMux I__7620 (
            .O(N__42845),
            .I(N__42831));
    LocalMux I__7619 (
            .O(N__42842),
            .I(encoder0_position_8));
    Odrv12 I__7618 (
            .O(N__42839),
            .I(encoder0_position_8));
    Odrv4 I__7617 (
            .O(N__42834),
            .I(encoder0_position_8));
    LocalMux I__7616 (
            .O(N__42831),
            .I(encoder0_position_8));
    InMux I__7615 (
            .O(N__42822),
            .I(N__42819));
    LocalMux I__7614 (
            .O(N__42819),
            .I(N__42815));
    InMux I__7613 (
            .O(N__42818),
            .I(N__42812));
    Span4Mux_h I__7612 (
            .O(N__42815),
            .I(N__42809));
    LocalMux I__7611 (
            .O(N__42812),
            .I(N__42806));
    Span4Mux_v I__7610 (
            .O(N__42809),
            .I(N__42803));
    Span4Mux_h I__7609 (
            .O(N__42806),
            .I(N__42800));
    Span4Mux_v I__7608 (
            .O(N__42803),
            .I(N__42797));
    Span4Mux_v I__7607 (
            .O(N__42800),
            .I(N__42794));
    Odrv4 I__7606 (
            .O(N__42797),
            .I(\c0.n22423 ));
    Odrv4 I__7605 (
            .O(N__42794),
            .I(\c0.n22423 ));
    CascadeMux I__7604 (
            .O(N__42789),
            .I(N__42784));
    CascadeMux I__7603 (
            .O(N__42788),
            .I(N__42781));
    InMux I__7602 (
            .O(N__42787),
            .I(N__42778));
    InMux I__7601 (
            .O(N__42784),
            .I(N__42775));
    InMux I__7600 (
            .O(N__42781),
            .I(N__42772));
    LocalMux I__7599 (
            .O(N__42778),
            .I(N__42767));
    LocalMux I__7598 (
            .O(N__42775),
            .I(N__42764));
    LocalMux I__7597 (
            .O(N__42772),
            .I(N__42761));
    InMux I__7596 (
            .O(N__42771),
            .I(N__42758));
    InMux I__7595 (
            .O(N__42770),
            .I(N__42755));
    Span4Mux_v I__7594 (
            .O(N__42767),
            .I(N__42752));
    Span4Mux_v I__7593 (
            .O(N__42764),
            .I(N__42749));
    Span4Mux_h I__7592 (
            .O(N__42761),
            .I(N__42746));
    LocalMux I__7591 (
            .O(N__42758),
            .I(N__42743));
    LocalMux I__7590 (
            .O(N__42755),
            .I(N__42738));
    Span4Mux_v I__7589 (
            .O(N__42752),
            .I(N__42738));
    Span4Mux_v I__7588 (
            .O(N__42749),
            .I(N__42733));
    Span4Mux_h I__7587 (
            .O(N__42746),
            .I(N__42733));
    Odrv4 I__7586 (
            .O(N__42743),
            .I(encoder0_position_6));
    Odrv4 I__7585 (
            .O(N__42738),
            .I(encoder0_position_6));
    Odrv4 I__7584 (
            .O(N__42733),
            .I(encoder0_position_6));
    InMux I__7583 (
            .O(N__42726),
            .I(N__42723));
    LocalMux I__7582 (
            .O(N__42723),
            .I(\c0.n6_adj_4293 ));
    CascadeMux I__7581 (
            .O(N__42720),
            .I(N__42717));
    InMux I__7580 (
            .O(N__42717),
            .I(N__42713));
    CascadeMux I__7579 (
            .O(N__42716),
            .I(N__42710));
    LocalMux I__7578 (
            .O(N__42713),
            .I(N__42707));
    InMux I__7577 (
            .O(N__42710),
            .I(N__42704));
    Span4Mux_h I__7576 (
            .O(N__42707),
            .I(N__42698));
    LocalMux I__7575 (
            .O(N__42704),
            .I(N__42695));
    InMux I__7574 (
            .O(N__42703),
            .I(N__42692));
    InMux I__7573 (
            .O(N__42702),
            .I(N__42689));
    InMux I__7572 (
            .O(N__42701),
            .I(N__42685));
    Span4Mux_h I__7571 (
            .O(N__42698),
            .I(N__42680));
    Span4Mux_v I__7570 (
            .O(N__42695),
            .I(N__42680));
    LocalMux I__7569 (
            .O(N__42692),
            .I(N__42675));
    LocalMux I__7568 (
            .O(N__42689),
            .I(N__42675));
    InMux I__7567 (
            .O(N__42688),
            .I(N__42672));
    LocalMux I__7566 (
            .O(N__42685),
            .I(encoder0_position_23));
    Odrv4 I__7565 (
            .O(N__42680),
            .I(encoder0_position_23));
    Odrv4 I__7564 (
            .O(N__42675),
            .I(encoder0_position_23));
    LocalMux I__7563 (
            .O(N__42672),
            .I(encoder0_position_23));
    InMux I__7562 (
            .O(N__42663),
            .I(N__42660));
    LocalMux I__7561 (
            .O(N__42660),
            .I(N__42652));
    InMux I__7560 (
            .O(N__42659),
            .I(N__42649));
    InMux I__7559 (
            .O(N__42658),
            .I(N__42646));
    InMux I__7558 (
            .O(N__42657),
            .I(N__42643));
    InMux I__7557 (
            .O(N__42656),
            .I(N__42640));
    InMux I__7556 (
            .O(N__42655),
            .I(N__42637));
    Sp12to4 I__7555 (
            .O(N__42652),
            .I(N__42632));
    LocalMux I__7554 (
            .O(N__42649),
            .I(N__42632));
    LocalMux I__7553 (
            .O(N__42646),
            .I(N__42629));
    LocalMux I__7552 (
            .O(N__42643),
            .I(encoder0_position_9));
    LocalMux I__7551 (
            .O(N__42640),
            .I(encoder0_position_9));
    LocalMux I__7550 (
            .O(N__42637),
            .I(encoder0_position_9));
    Odrv12 I__7549 (
            .O(N__42632),
            .I(encoder0_position_9));
    Odrv12 I__7548 (
            .O(N__42629),
            .I(encoder0_position_9));
    CascadeMux I__7547 (
            .O(N__42618),
            .I(N__42615));
    InMux I__7546 (
            .O(N__42615),
            .I(N__42612));
    LocalMux I__7545 (
            .O(N__42612),
            .I(N__42608));
    CascadeMux I__7544 (
            .O(N__42611),
            .I(N__42605));
    Span4Mux_v I__7543 (
            .O(N__42608),
            .I(N__42602));
    InMux I__7542 (
            .O(N__42605),
            .I(N__42598));
    Span4Mux_h I__7541 (
            .O(N__42602),
            .I(N__42594));
    InMux I__7540 (
            .O(N__42601),
            .I(N__42591));
    LocalMux I__7539 (
            .O(N__42598),
            .I(N__42588));
    InMux I__7538 (
            .O(N__42597),
            .I(N__42585));
    Span4Mux_h I__7537 (
            .O(N__42594),
            .I(N__42580));
    LocalMux I__7536 (
            .O(N__42591),
            .I(N__42580));
    Span12Mux_v I__7535 (
            .O(N__42588),
            .I(N__42577));
    LocalMux I__7534 (
            .O(N__42585),
            .I(control_mode_7));
    Odrv4 I__7533 (
            .O(N__42580),
            .I(control_mode_7));
    Odrv12 I__7532 (
            .O(N__42577),
            .I(control_mode_7));
    CascadeMux I__7531 (
            .O(N__42570),
            .I(\c0.n22385_cascade_ ));
    CascadeMux I__7530 (
            .O(N__42567),
            .I(N__42564));
    InMux I__7529 (
            .O(N__42564),
            .I(N__42561));
    LocalMux I__7528 (
            .O(N__42561),
            .I(N__42556));
    InMux I__7527 (
            .O(N__42560),
            .I(N__42553));
    InMux I__7526 (
            .O(N__42559),
            .I(N__42549));
    Span4Mux_h I__7525 (
            .O(N__42556),
            .I(N__42544));
    LocalMux I__7524 (
            .O(N__42553),
            .I(N__42544));
    InMux I__7523 (
            .O(N__42552),
            .I(N__42541));
    LocalMux I__7522 (
            .O(N__42549),
            .I(N__42538));
    Span4Mux_v I__7521 (
            .O(N__42544),
            .I(N__42532));
    LocalMux I__7520 (
            .O(N__42541),
            .I(N__42529));
    Span4Mux_h I__7519 (
            .O(N__42538),
            .I(N__42526));
    InMux I__7518 (
            .O(N__42537),
            .I(N__42523));
    InMux I__7517 (
            .O(N__42536),
            .I(N__42520));
    InMux I__7516 (
            .O(N__42535),
            .I(N__42517));
    Span4Mux_v I__7515 (
            .O(N__42532),
            .I(N__42514));
    Span4Mux_h I__7514 (
            .O(N__42529),
            .I(N__42509));
    Span4Mux_v I__7513 (
            .O(N__42526),
            .I(N__42509));
    LocalMux I__7512 (
            .O(N__42523),
            .I(encoder0_position_24));
    LocalMux I__7511 (
            .O(N__42520),
            .I(encoder0_position_24));
    LocalMux I__7510 (
            .O(N__42517),
            .I(encoder0_position_24));
    Odrv4 I__7509 (
            .O(N__42514),
            .I(encoder0_position_24));
    Odrv4 I__7508 (
            .O(N__42509),
            .I(encoder0_position_24));
    InMux I__7507 (
            .O(N__42498),
            .I(N__42494));
    InMux I__7506 (
            .O(N__42497),
            .I(N__42491));
    LocalMux I__7505 (
            .O(N__42494),
            .I(N__42488));
    LocalMux I__7504 (
            .O(N__42491),
            .I(N__42485));
    Span4Mux_h I__7503 (
            .O(N__42488),
            .I(N__42482));
    Span4Mux_v I__7502 (
            .O(N__42485),
            .I(N__42479));
    Span4Mux_v I__7501 (
            .O(N__42482),
            .I(N__42474));
    Span4Mux_h I__7500 (
            .O(N__42479),
            .I(N__42474));
    Odrv4 I__7499 (
            .O(N__42474),
            .I(\c0.n20325 ));
    InMux I__7498 (
            .O(N__42471),
            .I(N__42467));
    CascadeMux I__7497 (
            .O(N__42470),
            .I(N__42463));
    LocalMux I__7496 (
            .O(N__42467),
            .I(N__42459));
    InMux I__7495 (
            .O(N__42466),
            .I(N__42454));
    InMux I__7494 (
            .O(N__42463),
            .I(N__42454));
    InMux I__7493 (
            .O(N__42462),
            .I(N__42451));
    Span4Mux_v I__7492 (
            .O(N__42459),
            .I(N__42448));
    LocalMux I__7491 (
            .O(N__42454),
            .I(N__42445));
    LocalMux I__7490 (
            .O(N__42451),
            .I(data_in_2_5));
    Odrv4 I__7489 (
            .O(N__42448),
            .I(data_in_2_5));
    Odrv4 I__7488 (
            .O(N__42445),
            .I(data_in_2_5));
    InMux I__7487 (
            .O(N__42438),
            .I(N__42431));
    InMux I__7486 (
            .O(N__42437),
            .I(N__42431));
    InMux I__7485 (
            .O(N__42436),
            .I(N__42428));
    LocalMux I__7484 (
            .O(N__42431),
            .I(N__42424));
    LocalMux I__7483 (
            .O(N__42428),
            .I(N__42421));
    InMux I__7482 (
            .O(N__42427),
            .I(N__42418));
    Span4Mux_h I__7481 (
            .O(N__42424),
            .I(N__42415));
    Odrv4 I__7480 (
            .O(N__42421),
            .I(data_in_1_5));
    LocalMux I__7479 (
            .O(N__42418),
            .I(data_in_1_5));
    Odrv4 I__7478 (
            .O(N__42415),
            .I(data_in_1_5));
    CascadeMux I__7477 (
            .O(N__42408),
            .I(N__42405));
    InMux I__7476 (
            .O(N__42405),
            .I(N__42402));
    LocalMux I__7475 (
            .O(N__42402),
            .I(N__42397));
    InMux I__7474 (
            .O(N__42401),
            .I(N__42394));
    InMux I__7473 (
            .O(N__42400),
            .I(N__42391));
    Span4Mux_v I__7472 (
            .O(N__42397),
            .I(N__42382));
    LocalMux I__7471 (
            .O(N__42394),
            .I(N__42382));
    LocalMux I__7470 (
            .O(N__42391),
            .I(N__42382));
    InMux I__7469 (
            .O(N__42390),
            .I(N__42377));
    InMux I__7468 (
            .O(N__42389),
            .I(N__42374));
    Span4Mux_h I__7467 (
            .O(N__42382),
            .I(N__42371));
    InMux I__7466 (
            .O(N__42381),
            .I(N__42366));
    InMux I__7465 (
            .O(N__42380),
            .I(N__42366));
    LocalMux I__7464 (
            .O(N__42377),
            .I(N__42363));
    LocalMux I__7463 (
            .O(N__42374),
            .I(encoder0_position_19));
    Odrv4 I__7462 (
            .O(N__42371),
            .I(encoder0_position_19));
    LocalMux I__7461 (
            .O(N__42366),
            .I(encoder0_position_19));
    Odrv12 I__7460 (
            .O(N__42363),
            .I(encoder0_position_19));
    CascadeMux I__7459 (
            .O(N__42354),
            .I(\c0.n22199_cascade_ ));
    InMux I__7458 (
            .O(N__42351),
            .I(N__42348));
    LocalMux I__7457 (
            .O(N__42348),
            .I(N__42345));
    Span4Mux_h I__7456 (
            .O(N__42345),
            .I(N__42342));
    Span4Mux_v I__7455 (
            .O(N__42342),
            .I(N__42338));
    InMux I__7454 (
            .O(N__42341),
            .I(N__42335));
    Odrv4 I__7453 (
            .O(N__42338),
            .I(\c0.n22834 ));
    LocalMux I__7452 (
            .O(N__42335),
            .I(\c0.n22834 ));
    InMux I__7451 (
            .O(N__42330),
            .I(N__42325));
    CascadeMux I__7450 (
            .O(N__42329),
            .I(N__42322));
    InMux I__7449 (
            .O(N__42328),
            .I(N__42319));
    LocalMux I__7448 (
            .O(N__42325),
            .I(N__42316));
    InMux I__7447 (
            .O(N__42322),
            .I(N__42313));
    LocalMux I__7446 (
            .O(N__42319),
            .I(N__42308));
    Span4Mux_h I__7445 (
            .O(N__42316),
            .I(N__42308));
    LocalMux I__7444 (
            .O(N__42313),
            .I(N__42304));
    Span4Mux_v I__7443 (
            .O(N__42308),
            .I(N__42301));
    InMux I__7442 (
            .O(N__42307),
            .I(N__42298));
    Span4Mux_v I__7441 (
            .O(N__42304),
            .I(N__42292));
    Span4Mux_v I__7440 (
            .O(N__42301),
            .I(N__42292));
    LocalMux I__7439 (
            .O(N__42298),
            .I(N__42289));
    InMux I__7438 (
            .O(N__42297),
            .I(N__42285));
    Span4Mux_h I__7437 (
            .O(N__42292),
            .I(N__42282));
    Sp12to4 I__7436 (
            .O(N__42289),
            .I(N__42279));
    InMux I__7435 (
            .O(N__42288),
            .I(N__42276));
    LocalMux I__7434 (
            .O(N__42285),
            .I(encoder0_position_13));
    Odrv4 I__7433 (
            .O(N__42282),
            .I(encoder0_position_13));
    Odrv12 I__7432 (
            .O(N__42279),
            .I(encoder0_position_13));
    LocalMux I__7431 (
            .O(N__42276),
            .I(encoder0_position_13));
    InMux I__7430 (
            .O(N__42267),
            .I(N__42264));
    LocalMux I__7429 (
            .O(N__42264),
            .I(N__42258));
    InMux I__7428 (
            .O(N__42263),
            .I(N__42254));
    InMux I__7427 (
            .O(N__42262),
            .I(N__42251));
    InMux I__7426 (
            .O(N__42261),
            .I(N__42248));
    Span4Mux_h I__7425 (
            .O(N__42258),
            .I(N__42244));
    InMux I__7424 (
            .O(N__42257),
            .I(N__42241));
    LocalMux I__7423 (
            .O(N__42254),
            .I(N__42238));
    LocalMux I__7422 (
            .O(N__42251),
            .I(N__42235));
    LocalMux I__7421 (
            .O(N__42248),
            .I(N__42232));
    InMux I__7420 (
            .O(N__42247),
            .I(N__42229));
    Span4Mux_v I__7419 (
            .O(N__42244),
            .I(N__42226));
    LocalMux I__7418 (
            .O(N__42241),
            .I(N__42223));
    Span4Mux_v I__7417 (
            .O(N__42238),
            .I(N__42216));
    Span4Mux_v I__7416 (
            .O(N__42235),
            .I(N__42216));
    Span4Mux_v I__7415 (
            .O(N__42232),
            .I(N__42216));
    LocalMux I__7414 (
            .O(N__42229),
            .I(encoder0_position_22));
    Odrv4 I__7413 (
            .O(N__42226),
            .I(encoder0_position_22));
    Odrv4 I__7412 (
            .O(N__42223),
            .I(encoder0_position_22));
    Odrv4 I__7411 (
            .O(N__42216),
            .I(encoder0_position_22));
    InMux I__7410 (
            .O(N__42207),
            .I(N__42204));
    LocalMux I__7409 (
            .O(N__42204),
            .I(\c0.n6_adj_4366 ));
    InMux I__7408 (
            .O(N__42201),
            .I(N__42195));
    InMux I__7407 (
            .O(N__42200),
            .I(N__42195));
    LocalMux I__7406 (
            .O(N__42195),
            .I(N__42190));
    InMux I__7405 (
            .O(N__42194),
            .I(N__42187));
    InMux I__7404 (
            .O(N__42193),
            .I(N__42184));
    Sp12to4 I__7403 (
            .O(N__42190),
            .I(N__42181));
    LocalMux I__7402 (
            .O(N__42187),
            .I(data_in_2_0));
    LocalMux I__7401 (
            .O(N__42184),
            .I(data_in_2_0));
    Odrv12 I__7400 (
            .O(N__42181),
            .I(data_in_2_0));
    CascadeMux I__7399 (
            .O(N__42174),
            .I(N__42171));
    InMux I__7398 (
            .O(N__42171),
            .I(N__42167));
    InMux I__7397 (
            .O(N__42170),
            .I(N__42164));
    LocalMux I__7396 (
            .O(N__42167),
            .I(N__42161));
    LocalMux I__7395 (
            .O(N__42164),
            .I(N__42158));
    Span4Mux_h I__7394 (
            .O(N__42161),
            .I(N__42155));
    Odrv12 I__7393 (
            .O(N__42158),
            .I(\c0.n22635 ));
    Odrv4 I__7392 (
            .O(N__42155),
            .I(\c0.n22635 ));
    CascadeMux I__7391 (
            .O(N__42150),
            .I(\c0.n22256_cascade_ ));
    InMux I__7390 (
            .O(N__42147),
            .I(N__42144));
    LocalMux I__7389 (
            .O(N__42144),
            .I(N__42140));
    InMux I__7388 (
            .O(N__42143),
            .I(N__42137));
    Span4Mux_v I__7387 (
            .O(N__42140),
            .I(N__42134));
    LocalMux I__7386 (
            .O(N__42137),
            .I(N__42131));
    Span4Mux_h I__7385 (
            .O(N__42134),
            .I(N__42128));
    Odrv12 I__7384 (
            .O(N__42131),
            .I(\c0.n22772 ));
    Odrv4 I__7383 (
            .O(N__42128),
            .I(\c0.n22772 ));
    InMux I__7382 (
            .O(N__42123),
            .I(N__42118));
    CascadeMux I__7381 (
            .O(N__42122),
            .I(N__42115));
    InMux I__7380 (
            .O(N__42121),
            .I(N__42111));
    LocalMux I__7379 (
            .O(N__42118),
            .I(N__42108));
    InMux I__7378 (
            .O(N__42115),
            .I(N__42105));
    InMux I__7377 (
            .O(N__42114),
            .I(N__42102));
    LocalMux I__7376 (
            .O(N__42111),
            .I(data_in_1_3));
    Odrv4 I__7375 (
            .O(N__42108),
            .I(data_in_1_3));
    LocalMux I__7374 (
            .O(N__42105),
            .I(data_in_1_3));
    LocalMux I__7373 (
            .O(N__42102),
            .I(data_in_1_3));
    InMux I__7372 (
            .O(N__42093),
            .I(N__42088));
    InMux I__7371 (
            .O(N__42092),
            .I(N__42083));
    InMux I__7370 (
            .O(N__42091),
            .I(N__42083));
    LocalMux I__7369 (
            .O(N__42088),
            .I(data_in_3_4));
    LocalMux I__7368 (
            .O(N__42083),
            .I(data_in_3_4));
    InMux I__7367 (
            .O(N__42078),
            .I(N__42075));
    LocalMux I__7366 (
            .O(N__42075),
            .I(N__42072));
    Span4Mux_v I__7365 (
            .O(N__42072),
            .I(N__42069));
    Odrv4 I__7364 (
            .O(N__42069),
            .I(n2334));
    CascadeMux I__7363 (
            .O(N__42066),
            .I(N__42060));
    InMux I__7362 (
            .O(N__42065),
            .I(N__42057));
    InMux I__7361 (
            .O(N__42064),
            .I(N__42054));
    InMux I__7360 (
            .O(N__42063),
            .I(N__42049));
    InMux I__7359 (
            .O(N__42060),
            .I(N__42049));
    LocalMux I__7358 (
            .O(N__42057),
            .I(data_in_1_0));
    LocalMux I__7357 (
            .O(N__42054),
            .I(data_in_1_0));
    LocalMux I__7356 (
            .O(N__42049),
            .I(data_in_1_0));
    InMux I__7355 (
            .O(N__42042),
            .I(N__42039));
    LocalMux I__7354 (
            .O(N__42039),
            .I(N__42036));
    Span4Mux_v I__7353 (
            .O(N__42036),
            .I(N__42033));
    Span4Mux_v I__7352 (
            .O(N__42033),
            .I(N__42030));
    Odrv4 I__7351 (
            .O(N__42030),
            .I(n2349));
    InMux I__7350 (
            .O(N__42027),
            .I(N__42023));
    InMux I__7349 (
            .O(N__42026),
            .I(N__42019));
    LocalMux I__7348 (
            .O(N__42023),
            .I(N__42014));
    InMux I__7347 (
            .O(N__42022),
            .I(N__42011));
    LocalMux I__7346 (
            .O(N__42019),
            .I(N__42008));
    InMux I__7345 (
            .O(N__42018),
            .I(N__42004));
    InMux I__7344 (
            .O(N__42017),
            .I(N__42001));
    Span4Mux_v I__7343 (
            .O(N__42014),
            .I(N__41996));
    LocalMux I__7342 (
            .O(N__42011),
            .I(N__41996));
    Span4Mux_v I__7341 (
            .O(N__42008),
            .I(N__41993));
    InMux I__7340 (
            .O(N__42007),
            .I(N__41990));
    LocalMux I__7339 (
            .O(N__42004),
            .I(N__41987));
    LocalMux I__7338 (
            .O(N__42001),
            .I(N__41984));
    Span4Mux_v I__7337 (
            .O(N__41996),
            .I(N__41981));
    Sp12to4 I__7336 (
            .O(N__41993),
            .I(N__41978));
    LocalMux I__7335 (
            .O(N__41990),
            .I(N__41975));
    Span4Mux_h I__7334 (
            .O(N__41987),
            .I(N__41972));
    Span4Mux_v I__7333 (
            .O(N__41984),
            .I(N__41967));
    Span4Mux_v I__7332 (
            .O(N__41981),
            .I(N__41967));
    Span12Mux_h I__7331 (
            .O(N__41978),
            .I(N__41964));
    Span4Mux_h I__7330 (
            .O(N__41975),
            .I(N__41959));
    Span4Mux_v I__7329 (
            .O(N__41972),
            .I(N__41959));
    Odrv4 I__7328 (
            .O(N__41967),
            .I(\c0.rx.r_SM_Main_2_N_3680_2 ));
    Odrv12 I__7327 (
            .O(N__41964),
            .I(\c0.rx.r_SM_Main_2_N_3680_2 ));
    Odrv4 I__7326 (
            .O(N__41959),
            .I(\c0.rx.r_SM_Main_2_N_3680_2 ));
    CascadeMux I__7325 (
            .O(N__41952),
            .I(N__41949));
    InMux I__7324 (
            .O(N__41949),
            .I(N__41946));
    LocalMux I__7323 (
            .O(N__41946),
            .I(N__41940));
    InMux I__7322 (
            .O(N__41945),
            .I(N__41935));
    InMux I__7321 (
            .O(N__41944),
            .I(N__41935));
    InMux I__7320 (
            .O(N__41943),
            .I(N__41932));
    Odrv4 I__7319 (
            .O(N__41940),
            .I(\c0.n24028 ));
    LocalMux I__7318 (
            .O(N__41935),
            .I(\c0.n24028 ));
    LocalMux I__7317 (
            .O(N__41932),
            .I(\c0.n24028 ));
    CascadeMux I__7316 (
            .O(N__41925),
            .I(\c0.n14_adj_4478_cascade_ ));
    InMux I__7315 (
            .O(N__41922),
            .I(N__41916));
    InMux I__7314 (
            .O(N__41921),
            .I(N__41916));
    LocalMux I__7313 (
            .O(N__41916),
            .I(\c0.n22193 ));
    InMux I__7312 (
            .O(N__41913),
            .I(N__41908));
    InMux I__7311 (
            .O(N__41912),
            .I(N__41904));
    InMux I__7310 (
            .O(N__41911),
            .I(N__41901));
    LocalMux I__7309 (
            .O(N__41908),
            .I(N__41898));
    InMux I__7308 (
            .O(N__41907),
            .I(N__41895));
    LocalMux I__7307 (
            .O(N__41904),
            .I(N__41890));
    LocalMux I__7306 (
            .O(N__41901),
            .I(N__41890));
    Span12Mux_v I__7305 (
            .O(N__41898),
            .I(N__41885));
    LocalMux I__7304 (
            .O(N__41895),
            .I(N__41885));
    Span4Mux_v I__7303 (
            .O(N__41890),
            .I(N__41882));
    Odrv12 I__7302 (
            .O(N__41885),
            .I(\c0.n13422 ));
    Odrv4 I__7301 (
            .O(N__41882),
            .I(\c0.n13422 ));
    CascadeMux I__7300 (
            .O(N__41877),
            .I(N__41874));
    InMux I__7299 (
            .O(N__41874),
            .I(N__41871));
    LocalMux I__7298 (
            .O(N__41871),
            .I(N__41868));
    Odrv4 I__7297 (
            .O(N__41868),
            .I(\c0.n22722 ));
    InMux I__7296 (
            .O(N__41865),
            .I(N__41862));
    LocalMux I__7295 (
            .O(N__41862),
            .I(N__41858));
    InMux I__7294 (
            .O(N__41861),
            .I(N__41855));
    Odrv4 I__7293 (
            .O(N__41858),
            .I(data_out_frame_29__2__N_1748));
    LocalMux I__7292 (
            .O(N__41855),
            .I(data_out_frame_29__2__N_1748));
    InMux I__7291 (
            .O(N__41850),
            .I(N__41847));
    LocalMux I__7290 (
            .O(N__41847),
            .I(N__41844));
    Span12Mux_v I__7289 (
            .O(N__41844),
            .I(N__41841));
    Odrv12 I__7288 (
            .O(N__41841),
            .I(\c0.n19_adj_4720 ));
    CascadeMux I__7287 (
            .O(N__41838),
            .I(N__41834));
    InMux I__7286 (
            .O(N__41837),
            .I(N__41831));
    InMux I__7285 (
            .O(N__41834),
            .I(N__41828));
    LocalMux I__7284 (
            .O(N__41831),
            .I(N__41825));
    LocalMux I__7283 (
            .O(N__41828),
            .I(N__41822));
    Span4Mux_h I__7282 (
            .O(N__41825),
            .I(N__41815));
    Span4Mux_v I__7281 (
            .O(N__41822),
            .I(N__41815));
    InMux I__7280 (
            .O(N__41821),
            .I(N__41810));
    InMux I__7279 (
            .O(N__41820),
            .I(N__41810));
    Odrv4 I__7278 (
            .O(N__41815),
            .I(data_in_2_1));
    LocalMux I__7277 (
            .O(N__41810),
            .I(data_in_2_1));
    InMux I__7276 (
            .O(N__41805),
            .I(N__41802));
    LocalMux I__7275 (
            .O(N__41802),
            .I(N__41798));
    CascadeMux I__7274 (
            .O(N__41801),
            .I(N__41795));
    Span4Mux_h I__7273 (
            .O(N__41798),
            .I(N__41792));
    InMux I__7272 (
            .O(N__41795),
            .I(N__41789));
    Span4Mux_v I__7271 (
            .O(N__41792),
            .I(N__41786));
    LocalMux I__7270 (
            .O(N__41789),
            .I(data_out_frame_29_3));
    Odrv4 I__7269 (
            .O(N__41786),
            .I(data_out_frame_29_3));
    CascadeMux I__7268 (
            .O(N__41781),
            .I(N__41776));
    CascadeMux I__7267 (
            .O(N__41780),
            .I(N__41773));
    CascadeMux I__7266 (
            .O(N__41779),
            .I(N__41770));
    InMux I__7265 (
            .O(N__41776),
            .I(N__41767));
    InMux I__7264 (
            .O(N__41773),
            .I(N__41764));
    InMux I__7263 (
            .O(N__41770),
            .I(N__41761));
    LocalMux I__7262 (
            .O(N__41767),
            .I(N__41757));
    LocalMux I__7261 (
            .O(N__41764),
            .I(N__41754));
    LocalMux I__7260 (
            .O(N__41761),
            .I(N__41749));
    InMux I__7259 (
            .O(N__41760),
            .I(N__41746));
    Span12Mux_v I__7258 (
            .O(N__41757),
            .I(N__41743));
    Span12Mux_h I__7257 (
            .O(N__41754),
            .I(N__41740));
    InMux I__7256 (
            .O(N__41753),
            .I(N__41737));
    InMux I__7255 (
            .O(N__41752),
            .I(N__41734));
    Span4Mux_v I__7254 (
            .O(N__41749),
            .I(N__41731));
    LocalMux I__7253 (
            .O(N__41746),
            .I(encoder1_position_12));
    Odrv12 I__7252 (
            .O(N__41743),
            .I(encoder1_position_12));
    Odrv12 I__7251 (
            .O(N__41740),
            .I(encoder1_position_12));
    LocalMux I__7250 (
            .O(N__41737),
            .I(encoder1_position_12));
    LocalMux I__7249 (
            .O(N__41734),
            .I(encoder1_position_12));
    Odrv4 I__7248 (
            .O(N__41731),
            .I(encoder1_position_12));
    InMux I__7247 (
            .O(N__41718),
            .I(N__41715));
    LocalMux I__7246 (
            .O(N__41715),
            .I(N__41711));
    InMux I__7245 (
            .O(N__41714),
            .I(N__41708));
    Span4Mux_v I__7244 (
            .O(N__41711),
            .I(N__41705));
    LocalMux I__7243 (
            .O(N__41708),
            .I(data_out_frame_12_4));
    Odrv4 I__7242 (
            .O(N__41705),
            .I(data_out_frame_12_4));
    InMux I__7241 (
            .O(N__41700),
            .I(N__41695));
    InMux I__7240 (
            .O(N__41699),
            .I(N__41692));
    InMux I__7239 (
            .O(N__41698),
            .I(N__41689));
    LocalMux I__7238 (
            .O(N__41695),
            .I(data_in_0_3));
    LocalMux I__7237 (
            .O(N__41692),
            .I(data_in_0_3));
    LocalMux I__7236 (
            .O(N__41689),
            .I(data_in_0_3));
    InMux I__7235 (
            .O(N__41682),
            .I(N__41679));
    LocalMux I__7234 (
            .O(N__41679),
            .I(N__41676));
    Span4Mux_h I__7233 (
            .O(N__41676),
            .I(N__41673));
    Odrv4 I__7232 (
            .O(N__41673),
            .I(\c0.n15 ));
    CascadeMux I__7231 (
            .O(N__41670),
            .I(\c0.n21311_cascade_ ));
    InMux I__7230 (
            .O(N__41667),
            .I(N__41664));
    LocalMux I__7229 (
            .O(N__41664),
            .I(N__41661));
    Span4Mux_v I__7228 (
            .O(N__41661),
            .I(N__41658));
    Span4Mux_h I__7227 (
            .O(N__41658),
            .I(N__41654));
    InMux I__7226 (
            .O(N__41657),
            .I(N__41651));
    Odrv4 I__7225 (
            .O(N__41654),
            .I(\c0.n21244 ));
    LocalMux I__7224 (
            .O(N__41651),
            .I(\c0.n21244 ));
    InMux I__7223 (
            .O(N__41646),
            .I(N__41643));
    LocalMux I__7222 (
            .O(N__41643),
            .I(N__41640));
    Span4Mux_h I__7221 (
            .O(N__41640),
            .I(N__41636));
    InMux I__7220 (
            .O(N__41639),
            .I(N__41633));
    Span4Mux_h I__7219 (
            .O(N__41636),
            .I(N__41630));
    LocalMux I__7218 (
            .O(N__41633),
            .I(\c0.n21496 ));
    Odrv4 I__7217 (
            .O(N__41630),
            .I(\c0.n21496 ));
    CascadeMux I__7216 (
            .O(N__41625),
            .I(\c0.n21273_cascade_ ));
    InMux I__7215 (
            .O(N__41622),
            .I(N__41619));
    LocalMux I__7214 (
            .O(N__41619),
            .I(N__41616));
    Span4Mux_h I__7213 (
            .O(N__41616),
            .I(N__41613));
    Odrv4 I__7212 (
            .O(N__41613),
            .I(\c0.data_out_frame_29_6 ));
    InMux I__7211 (
            .O(N__41610),
            .I(N__41607));
    LocalMux I__7210 (
            .O(N__41607),
            .I(N__41604));
    Odrv4 I__7209 (
            .O(N__41604),
            .I(\c0.data_out_frame_28_6 ));
    InMux I__7208 (
            .O(N__41601),
            .I(N__41598));
    LocalMux I__7207 (
            .O(N__41598),
            .I(N__41595));
    Span12Mux_h I__7206 (
            .O(N__41595),
            .I(N__41592));
    Odrv12 I__7205 (
            .O(N__41592),
            .I(\c0.n26_adj_4702 ));
    InMux I__7204 (
            .O(N__41589),
            .I(N__41585));
    InMux I__7203 (
            .O(N__41588),
            .I(N__41582));
    LocalMux I__7202 (
            .O(N__41585),
            .I(N__41577));
    LocalMux I__7201 (
            .O(N__41582),
            .I(N__41577));
    Span4Mux_h I__7200 (
            .O(N__41577),
            .I(N__41574));
    Odrv4 I__7199 (
            .O(N__41574),
            .I(\c0.n22617 ));
    InMux I__7198 (
            .O(N__41571),
            .I(N__41568));
    LocalMux I__7197 (
            .O(N__41568),
            .I(N__41565));
    Span4Mux_v I__7196 (
            .O(N__41565),
            .I(N__41559));
    InMux I__7195 (
            .O(N__41564),
            .I(N__41556));
    InMux I__7194 (
            .O(N__41563),
            .I(N__41551));
    InMux I__7193 (
            .O(N__41562),
            .I(N__41551));
    Span4Mux_h I__7192 (
            .O(N__41559),
            .I(N__41546));
    LocalMux I__7191 (
            .O(N__41556),
            .I(N__41546));
    LocalMux I__7190 (
            .O(N__41551),
            .I(\c0.n20341 ));
    Odrv4 I__7189 (
            .O(N__41546),
            .I(\c0.n20341 ));
    CascadeMux I__7188 (
            .O(N__41541),
            .I(\c0.n18_adj_4684_cascade_ ));
    InMux I__7187 (
            .O(N__41538),
            .I(N__41532));
    InMux I__7186 (
            .O(N__41537),
            .I(N__41529));
    InMux I__7185 (
            .O(N__41536),
            .I(N__41524));
    InMux I__7184 (
            .O(N__41535),
            .I(N__41524));
    LocalMux I__7183 (
            .O(N__41532),
            .I(\c0.n13268 ));
    LocalMux I__7182 (
            .O(N__41529),
            .I(\c0.n13268 ));
    LocalMux I__7181 (
            .O(N__41524),
            .I(\c0.n13268 ));
    InMux I__7180 (
            .O(N__41517),
            .I(N__41514));
    LocalMux I__7179 (
            .O(N__41514),
            .I(N__41511));
    Span4Mux_v I__7178 (
            .O(N__41511),
            .I(N__41508));
    Odrv4 I__7177 (
            .O(N__41508),
            .I(\c0.n15_adj_4686 ));
    CascadeMux I__7176 (
            .O(N__41505),
            .I(\c0.n20_adj_4685_cascade_ ));
    InMux I__7175 (
            .O(N__41502),
            .I(N__41499));
    LocalMux I__7174 (
            .O(N__41499),
            .I(N__41496));
    Span4Mux_h I__7173 (
            .O(N__41496),
            .I(N__41492));
    InMux I__7172 (
            .O(N__41495),
            .I(N__41488));
    Span4Mux_h I__7171 (
            .O(N__41492),
            .I(N__41485));
    InMux I__7170 (
            .O(N__41491),
            .I(N__41482));
    LocalMux I__7169 (
            .O(N__41488),
            .I(N__41479));
    Odrv4 I__7168 (
            .O(N__41485),
            .I(\c0.n21475 ));
    LocalMux I__7167 (
            .O(N__41482),
            .I(\c0.n21475 ));
    Odrv4 I__7166 (
            .O(N__41479),
            .I(\c0.n21475 ));
    InMux I__7165 (
            .O(N__41472),
            .I(N__41469));
    LocalMux I__7164 (
            .O(N__41469),
            .I(N__41466));
    Span4Mux_v I__7163 (
            .O(N__41466),
            .I(N__41463));
    Span4Mux_h I__7162 (
            .O(N__41463),
            .I(N__41460));
    Sp12to4 I__7161 (
            .O(N__41460),
            .I(N__41457));
    Odrv12 I__7160 (
            .O(N__41457),
            .I(\c0.data_out_frame_28_7 ));
    InMux I__7159 (
            .O(N__41454),
            .I(N__41451));
    LocalMux I__7158 (
            .O(N__41451),
            .I(\c0.n22461 ));
    InMux I__7157 (
            .O(N__41448),
            .I(N__41444));
    InMux I__7156 (
            .O(N__41447),
            .I(N__41441));
    LocalMux I__7155 (
            .O(N__41444),
            .I(\c0.n21358 ));
    LocalMux I__7154 (
            .O(N__41441),
            .I(\c0.n21358 ));
    CascadeMux I__7153 (
            .O(N__41436),
            .I(\c0.n22461_cascade_ ));
    InMux I__7152 (
            .O(N__41433),
            .I(N__41426));
    InMux I__7151 (
            .O(N__41432),
            .I(N__41423));
    InMux I__7150 (
            .O(N__41431),
            .I(N__41420));
    InMux I__7149 (
            .O(N__41430),
            .I(N__41417));
    InMux I__7148 (
            .O(N__41429),
            .I(N__41414));
    LocalMux I__7147 (
            .O(N__41426),
            .I(N__41409));
    LocalMux I__7146 (
            .O(N__41423),
            .I(N__41400));
    LocalMux I__7145 (
            .O(N__41420),
            .I(N__41400));
    LocalMux I__7144 (
            .O(N__41417),
            .I(N__41400));
    LocalMux I__7143 (
            .O(N__41414),
            .I(N__41400));
    InMux I__7142 (
            .O(N__41413),
            .I(N__41397));
    InMux I__7141 (
            .O(N__41412),
            .I(N__41394));
    Span4Mux_v I__7140 (
            .O(N__41409),
            .I(N__41391));
    Span4Mux_v I__7139 (
            .O(N__41400),
            .I(N__41386));
    LocalMux I__7138 (
            .O(N__41397),
            .I(N__41386));
    LocalMux I__7137 (
            .O(N__41394),
            .I(N__41383));
    Span4Mux_v I__7136 (
            .O(N__41391),
            .I(N__41378));
    Span4Mux_v I__7135 (
            .O(N__41386),
            .I(N__41378));
    Span4Mux_h I__7134 (
            .O(N__41383),
            .I(N__41375));
    Odrv4 I__7133 (
            .O(N__41378),
            .I(\c0.n21406 ));
    Odrv4 I__7132 (
            .O(N__41375),
            .I(\c0.n21406 ));
    InMux I__7131 (
            .O(N__41370),
            .I(N__41367));
    LocalMux I__7130 (
            .O(N__41367),
            .I(N__41361));
    InMux I__7129 (
            .O(N__41366),
            .I(N__41358));
    InMux I__7128 (
            .O(N__41365),
            .I(N__41355));
    InMux I__7127 (
            .O(N__41364),
            .I(N__41352));
    Span4Mux_v I__7126 (
            .O(N__41361),
            .I(N__41347));
    LocalMux I__7125 (
            .O(N__41358),
            .I(N__41347));
    LocalMux I__7124 (
            .O(N__41355),
            .I(N__41342));
    LocalMux I__7123 (
            .O(N__41352),
            .I(N__41342));
    Span4Mux_h I__7122 (
            .O(N__41347),
            .I(N__41339));
    Odrv12 I__7121 (
            .O(N__41342),
            .I(\c0.n21441 ));
    Odrv4 I__7120 (
            .O(N__41339),
            .I(\c0.n21441 ));
    CascadeMux I__7119 (
            .O(N__41334),
            .I(N__41331));
    InMux I__7118 (
            .O(N__41331),
            .I(N__41328));
    LocalMux I__7117 (
            .O(N__41328),
            .I(N__41322));
    CascadeMux I__7116 (
            .O(N__41327),
            .I(N__41319));
    InMux I__7115 (
            .O(N__41326),
            .I(N__41314));
    InMux I__7114 (
            .O(N__41325),
            .I(N__41311));
    Span4Mux_h I__7113 (
            .O(N__41322),
            .I(N__41308));
    InMux I__7112 (
            .O(N__41319),
            .I(N__41305));
    InMux I__7111 (
            .O(N__41318),
            .I(N__41302));
    InMux I__7110 (
            .O(N__41317),
            .I(N__41299));
    LocalMux I__7109 (
            .O(N__41314),
            .I(N__41296));
    LocalMux I__7108 (
            .O(N__41311),
            .I(encoder0_position_25));
    Odrv4 I__7107 (
            .O(N__41308),
            .I(encoder0_position_25));
    LocalMux I__7106 (
            .O(N__41305),
            .I(encoder0_position_25));
    LocalMux I__7105 (
            .O(N__41302),
            .I(encoder0_position_25));
    LocalMux I__7104 (
            .O(N__41299),
            .I(encoder0_position_25));
    Odrv4 I__7103 (
            .O(N__41296),
            .I(encoder0_position_25));
    InMux I__7102 (
            .O(N__41283),
            .I(N__41280));
    LocalMux I__7101 (
            .O(N__41280),
            .I(N__41277));
    Span4Mux_v I__7100 (
            .O(N__41277),
            .I(N__41273));
    InMux I__7099 (
            .O(N__41276),
            .I(N__41270));
    Span4Mux_h I__7098 (
            .O(N__41273),
            .I(N__41267));
    LocalMux I__7097 (
            .O(N__41270),
            .I(data_out_frame_6_1));
    Odrv4 I__7096 (
            .O(N__41267),
            .I(data_out_frame_6_1));
    InMux I__7095 (
            .O(N__41262),
            .I(N__41258));
    CascadeMux I__7094 (
            .O(N__41261),
            .I(N__41255));
    LocalMux I__7093 (
            .O(N__41258),
            .I(N__41252));
    InMux I__7092 (
            .O(N__41255),
            .I(N__41249));
    Span4Mux_h I__7091 (
            .O(N__41252),
            .I(N__41246));
    LocalMux I__7090 (
            .O(N__41249),
            .I(data_out_frame_29_2));
    Odrv4 I__7089 (
            .O(N__41246),
            .I(data_out_frame_29_2));
    InMux I__7088 (
            .O(N__41241),
            .I(N__41238));
    LocalMux I__7087 (
            .O(N__41238),
            .I(\c0.n12_adj_4312 ));
    CascadeMux I__7086 (
            .O(N__41235),
            .I(\c0.n24113_cascade_ ));
    InMux I__7085 (
            .O(N__41232),
            .I(N__41226));
    InMux I__7084 (
            .O(N__41231),
            .I(N__41223));
    InMux I__7083 (
            .O(N__41230),
            .I(N__41220));
    InMux I__7082 (
            .O(N__41229),
            .I(N__41217));
    LocalMux I__7081 (
            .O(N__41226),
            .I(N__41214));
    LocalMux I__7080 (
            .O(N__41223),
            .I(N__41211));
    LocalMux I__7079 (
            .O(N__41220),
            .I(N__41208));
    LocalMux I__7078 (
            .O(N__41217),
            .I(N__41205));
    Span4Mux_h I__7077 (
            .O(N__41214),
            .I(N__41202));
    Span4Mux_v I__7076 (
            .O(N__41211),
            .I(N__41197));
    Span4Mux_v I__7075 (
            .O(N__41208),
            .I(N__41197));
    Odrv4 I__7074 (
            .O(N__41205),
            .I(\c0.n10529 ));
    Odrv4 I__7073 (
            .O(N__41202),
            .I(\c0.n10529 ));
    Odrv4 I__7072 (
            .O(N__41197),
            .I(\c0.n10529 ));
    InMux I__7071 (
            .O(N__41190),
            .I(N__41186));
    CascadeMux I__7070 (
            .O(N__41189),
            .I(N__41182));
    LocalMux I__7069 (
            .O(N__41186),
            .I(N__41176));
    InMux I__7068 (
            .O(N__41185),
            .I(N__41173));
    InMux I__7067 (
            .O(N__41182),
            .I(N__41169));
    InMux I__7066 (
            .O(N__41181),
            .I(N__41164));
    InMux I__7065 (
            .O(N__41180),
            .I(N__41164));
    InMux I__7064 (
            .O(N__41179),
            .I(N__41161));
    Span4Mux_v I__7063 (
            .O(N__41176),
            .I(N__41156));
    LocalMux I__7062 (
            .O(N__41173),
            .I(N__41156));
    CascadeMux I__7061 (
            .O(N__41172),
            .I(N__41153));
    LocalMux I__7060 (
            .O(N__41169),
            .I(N__41148));
    LocalMux I__7059 (
            .O(N__41164),
            .I(N__41148));
    LocalMux I__7058 (
            .O(N__41161),
            .I(N__41143));
    Span4Mux_v I__7057 (
            .O(N__41156),
            .I(N__41143));
    InMux I__7056 (
            .O(N__41153),
            .I(N__41140));
    Span4Mux_v I__7055 (
            .O(N__41148),
            .I(N__41136));
    Span4Mux_h I__7054 (
            .O(N__41143),
            .I(N__41131));
    LocalMux I__7053 (
            .O(N__41140),
            .I(N__41131));
    InMux I__7052 (
            .O(N__41139),
            .I(N__41128));
    Span4Mux_h I__7051 (
            .O(N__41136),
            .I(N__41125));
    Span4Mux_h I__7050 (
            .O(N__41131),
            .I(N__41122));
    LocalMux I__7049 (
            .O(N__41128),
            .I(encoder1_position_5));
    Odrv4 I__7048 (
            .O(N__41125),
            .I(encoder1_position_5));
    Odrv4 I__7047 (
            .O(N__41122),
            .I(encoder1_position_5));
    CascadeMux I__7046 (
            .O(N__41115),
            .I(N__41112));
    InMux I__7045 (
            .O(N__41112),
            .I(N__41109));
    LocalMux I__7044 (
            .O(N__41109),
            .I(N__41099));
    InMux I__7043 (
            .O(N__41108),
            .I(N__41094));
    InMux I__7042 (
            .O(N__41107),
            .I(N__41094));
    InMux I__7041 (
            .O(N__41106),
            .I(N__41089));
    InMux I__7040 (
            .O(N__41105),
            .I(N__41089));
    InMux I__7039 (
            .O(N__41104),
            .I(N__41086));
    InMux I__7038 (
            .O(N__41103),
            .I(N__41081));
    InMux I__7037 (
            .O(N__41102),
            .I(N__41081));
    Span4Mux_h I__7036 (
            .O(N__41099),
            .I(N__41074));
    LocalMux I__7035 (
            .O(N__41094),
            .I(N__41074));
    LocalMux I__7034 (
            .O(N__41089),
            .I(N__41074));
    LocalMux I__7033 (
            .O(N__41086),
            .I(\c0.n21364 ));
    LocalMux I__7032 (
            .O(N__41081),
            .I(\c0.n21364 ));
    Odrv4 I__7031 (
            .O(N__41074),
            .I(\c0.n21364 ));
    InMux I__7030 (
            .O(N__41067),
            .I(N__41063));
    InMux I__7029 (
            .O(N__41066),
            .I(N__41060));
    LocalMux I__7028 (
            .O(N__41063),
            .I(\c0.n24113 ));
    LocalMux I__7027 (
            .O(N__41060),
            .I(\c0.n24113 ));
    InMux I__7026 (
            .O(N__41055),
            .I(N__41050));
    InMux I__7025 (
            .O(N__41054),
            .I(N__41047));
    InMux I__7024 (
            .O(N__41053),
            .I(N__41042));
    LocalMux I__7023 (
            .O(N__41050),
            .I(N__41039));
    LocalMux I__7022 (
            .O(N__41047),
            .I(N__41035));
    InMux I__7021 (
            .O(N__41046),
            .I(N__41030));
    InMux I__7020 (
            .O(N__41045),
            .I(N__41027));
    LocalMux I__7019 (
            .O(N__41042),
            .I(N__41014));
    Span4Mux_v I__7018 (
            .O(N__41039),
            .I(N__41011));
    InMux I__7017 (
            .O(N__41038),
            .I(N__41005));
    Span4Mux_v I__7016 (
            .O(N__41035),
            .I(N__41002));
    InMux I__7015 (
            .O(N__41034),
            .I(N__40997));
    CascadeMux I__7014 (
            .O(N__41033),
            .I(N__40991));
    LocalMux I__7013 (
            .O(N__41030),
            .I(N__40986));
    LocalMux I__7012 (
            .O(N__41027),
            .I(N__40986));
    InMux I__7011 (
            .O(N__41026),
            .I(N__40983));
    InMux I__7010 (
            .O(N__41025),
            .I(N__40980));
    InMux I__7009 (
            .O(N__41024),
            .I(N__40973));
    InMux I__7008 (
            .O(N__41023),
            .I(N__40973));
    InMux I__7007 (
            .O(N__41022),
            .I(N__40973));
    InMux I__7006 (
            .O(N__41021),
            .I(N__40966));
    InMux I__7005 (
            .O(N__41020),
            .I(N__40966));
    InMux I__7004 (
            .O(N__41019),
            .I(N__40966));
    InMux I__7003 (
            .O(N__41018),
            .I(N__40961));
    InMux I__7002 (
            .O(N__41017),
            .I(N__40961));
    Span4Mux_v I__7001 (
            .O(N__41014),
            .I(N__40958));
    Span4Mux_v I__7000 (
            .O(N__41011),
            .I(N__40955));
    InMux I__6999 (
            .O(N__41010),
            .I(N__40950));
    InMux I__6998 (
            .O(N__41009),
            .I(N__40950));
    InMux I__6997 (
            .O(N__41008),
            .I(N__40946));
    LocalMux I__6996 (
            .O(N__41005),
            .I(N__40941));
    Span4Mux_v I__6995 (
            .O(N__41002),
            .I(N__40941));
    InMux I__6994 (
            .O(N__41001),
            .I(N__40936));
    InMux I__6993 (
            .O(N__41000),
            .I(N__40936));
    LocalMux I__6992 (
            .O(N__40997),
            .I(N__40933));
    InMux I__6991 (
            .O(N__40996),
            .I(N__40930));
    InMux I__6990 (
            .O(N__40995),
            .I(N__40926));
    InMux I__6989 (
            .O(N__40994),
            .I(N__40923));
    InMux I__6988 (
            .O(N__40991),
            .I(N__40920));
    Span4Mux_v I__6987 (
            .O(N__40986),
            .I(N__40913));
    LocalMux I__6986 (
            .O(N__40983),
            .I(N__40913));
    LocalMux I__6985 (
            .O(N__40980),
            .I(N__40913));
    LocalMux I__6984 (
            .O(N__40973),
            .I(N__40904));
    LocalMux I__6983 (
            .O(N__40966),
            .I(N__40904));
    LocalMux I__6982 (
            .O(N__40961),
            .I(N__40904));
    Span4Mux_v I__6981 (
            .O(N__40958),
            .I(N__40904));
    Span4Mux_v I__6980 (
            .O(N__40955),
            .I(N__40901));
    LocalMux I__6979 (
            .O(N__40950),
            .I(N__40898));
    InMux I__6978 (
            .O(N__40949),
            .I(N__40895));
    LocalMux I__6977 (
            .O(N__40946),
            .I(N__40890));
    Span4Mux_h I__6976 (
            .O(N__40941),
            .I(N__40890));
    LocalMux I__6975 (
            .O(N__40936),
            .I(N__40883));
    Span4Mux_h I__6974 (
            .O(N__40933),
            .I(N__40883));
    LocalMux I__6973 (
            .O(N__40930),
            .I(N__40883));
    InMux I__6972 (
            .O(N__40929),
            .I(N__40880));
    LocalMux I__6971 (
            .O(N__40926),
            .I(N__40867));
    LocalMux I__6970 (
            .O(N__40923),
            .I(N__40867));
    LocalMux I__6969 (
            .O(N__40920),
            .I(N__40867));
    Span4Mux_v I__6968 (
            .O(N__40913),
            .I(N__40867));
    Span4Mux_v I__6967 (
            .O(N__40904),
            .I(N__40867));
    Span4Mux_h I__6966 (
            .O(N__40901),
            .I(N__40867));
    Odrv12 I__6965 (
            .O(N__40898),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__6964 (
            .O(N__40895),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__6963 (
            .O(N__40890),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__6962 (
            .O(N__40883),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__6961 (
            .O(N__40880),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__6960 (
            .O(N__40867),
            .I(\c0.byte_transmit_counter_2 ));
    InMux I__6959 (
            .O(N__40854),
            .I(N__40851));
    LocalMux I__6958 (
            .O(N__40851),
            .I(N__40848));
    Span4Mux_h I__6957 (
            .O(N__40848),
            .I(N__40845));
    Span4Mux_v I__6956 (
            .O(N__40845),
            .I(N__40842));
    Span4Mux_v I__6955 (
            .O(N__40842),
            .I(N__40839));
    Odrv4 I__6954 (
            .O(N__40839),
            .I(\c0.n5_adj_4217 ));
    CascadeMux I__6953 (
            .O(N__40836),
            .I(N__40832));
    InMux I__6952 (
            .O(N__40835),
            .I(N__40829));
    InMux I__6951 (
            .O(N__40832),
            .I(N__40826));
    LocalMux I__6950 (
            .O(N__40829),
            .I(N__40823));
    LocalMux I__6949 (
            .O(N__40826),
            .I(N__40812));
    Span4Mux_v I__6948 (
            .O(N__40823),
            .I(N__40801));
    InMux I__6947 (
            .O(N__40822),
            .I(N__40796));
    InMux I__6946 (
            .O(N__40821),
            .I(N__40796));
    InMux I__6945 (
            .O(N__40820),
            .I(N__40793));
    InMux I__6944 (
            .O(N__40819),
            .I(N__40790));
    InMux I__6943 (
            .O(N__40818),
            .I(N__40787));
    InMux I__6942 (
            .O(N__40817),
            .I(N__40782));
    InMux I__6941 (
            .O(N__40816),
            .I(N__40782));
    CascadeMux I__6940 (
            .O(N__40815),
            .I(N__40764));
    Span4Mux_v I__6939 (
            .O(N__40812),
            .I(N__40761));
    InMux I__6938 (
            .O(N__40811),
            .I(N__40758));
    InMux I__6937 (
            .O(N__40810),
            .I(N__40755));
    InMux I__6936 (
            .O(N__40809),
            .I(N__40746));
    InMux I__6935 (
            .O(N__40808),
            .I(N__40746));
    InMux I__6934 (
            .O(N__40807),
            .I(N__40746));
    InMux I__6933 (
            .O(N__40806),
            .I(N__40746));
    InMux I__6932 (
            .O(N__40805),
            .I(N__40741));
    InMux I__6931 (
            .O(N__40804),
            .I(N__40741));
    Span4Mux_v I__6930 (
            .O(N__40801),
            .I(N__40736));
    LocalMux I__6929 (
            .O(N__40796),
            .I(N__40736));
    LocalMux I__6928 (
            .O(N__40793),
            .I(N__40727));
    LocalMux I__6927 (
            .O(N__40790),
            .I(N__40727));
    LocalMux I__6926 (
            .O(N__40787),
            .I(N__40727));
    LocalMux I__6925 (
            .O(N__40782),
            .I(N__40727));
    InMux I__6924 (
            .O(N__40781),
            .I(N__40720));
    InMux I__6923 (
            .O(N__40780),
            .I(N__40720));
    InMux I__6922 (
            .O(N__40779),
            .I(N__40720));
    InMux I__6921 (
            .O(N__40778),
            .I(N__40715));
    InMux I__6920 (
            .O(N__40777),
            .I(N__40715));
    InMux I__6919 (
            .O(N__40776),
            .I(N__40706));
    InMux I__6918 (
            .O(N__40775),
            .I(N__40706));
    InMux I__6917 (
            .O(N__40774),
            .I(N__40706));
    InMux I__6916 (
            .O(N__40773),
            .I(N__40706));
    InMux I__6915 (
            .O(N__40772),
            .I(N__40703));
    InMux I__6914 (
            .O(N__40771),
            .I(N__40694));
    InMux I__6913 (
            .O(N__40770),
            .I(N__40694));
    InMux I__6912 (
            .O(N__40769),
            .I(N__40694));
    InMux I__6911 (
            .O(N__40768),
            .I(N__40694));
    InMux I__6910 (
            .O(N__40767),
            .I(N__40689));
    InMux I__6909 (
            .O(N__40764),
            .I(N__40689));
    Span4Mux_h I__6908 (
            .O(N__40761),
            .I(N__40686));
    LocalMux I__6907 (
            .O(N__40758),
            .I(N__40681));
    LocalMux I__6906 (
            .O(N__40755),
            .I(N__40672));
    LocalMux I__6905 (
            .O(N__40746),
            .I(N__40672));
    LocalMux I__6904 (
            .O(N__40741),
            .I(N__40672));
    Span4Mux_h I__6903 (
            .O(N__40736),
            .I(N__40672));
    Span4Mux_v I__6902 (
            .O(N__40727),
            .I(N__40667));
    LocalMux I__6901 (
            .O(N__40720),
            .I(N__40667));
    LocalMux I__6900 (
            .O(N__40715),
            .I(N__40654));
    LocalMux I__6899 (
            .O(N__40706),
            .I(N__40654));
    LocalMux I__6898 (
            .O(N__40703),
            .I(N__40654));
    LocalMux I__6897 (
            .O(N__40694),
            .I(N__40654));
    LocalMux I__6896 (
            .O(N__40689),
            .I(N__40654));
    Span4Mux_v I__6895 (
            .O(N__40686),
            .I(N__40654));
    CascadeMux I__6894 (
            .O(N__40685),
            .I(N__40651));
    InMux I__6893 (
            .O(N__40684),
            .I(N__40645));
    Span4Mux_v I__6892 (
            .O(N__40681),
            .I(N__40642));
    Span4Mux_h I__6891 (
            .O(N__40672),
            .I(N__40639));
    Span4Mux_v I__6890 (
            .O(N__40667),
            .I(N__40634));
    Span4Mux_v I__6889 (
            .O(N__40654),
            .I(N__40634));
    InMux I__6888 (
            .O(N__40651),
            .I(N__40627));
    InMux I__6887 (
            .O(N__40650),
            .I(N__40627));
    InMux I__6886 (
            .O(N__40649),
            .I(N__40627));
    InMux I__6885 (
            .O(N__40648),
            .I(N__40624));
    LocalMux I__6884 (
            .O(N__40645),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6883 (
            .O(N__40642),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6882 (
            .O(N__40639),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6881 (
            .O(N__40634),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__6880 (
            .O(N__40627),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__6879 (
            .O(N__40624),
            .I(\c0.byte_transmit_counter_1 ));
    InMux I__6878 (
            .O(N__40611),
            .I(N__40608));
    LocalMux I__6877 (
            .O(N__40608),
            .I(N__40605));
    Span4Mux_h I__6876 (
            .O(N__40605),
            .I(N__40602));
    Odrv4 I__6875 (
            .O(N__40602),
            .I(\c0.n24901 ));
    InMux I__6874 (
            .O(N__40599),
            .I(N__40596));
    LocalMux I__6873 (
            .O(N__40596),
            .I(N__40593));
    Odrv12 I__6872 (
            .O(N__40593),
            .I(\c0.n25062 ));
    InMux I__6871 (
            .O(N__40590),
            .I(N__40587));
    LocalMux I__6870 (
            .O(N__40587),
            .I(N__40584));
    Span4Mux_h I__6869 (
            .O(N__40584),
            .I(N__40581));
    Span4Mux_v I__6868 (
            .O(N__40581),
            .I(N__40578));
    Odrv4 I__6867 (
            .O(N__40578),
            .I(n2260));
    CascadeMux I__6866 (
            .O(N__40575),
            .I(N__40570));
    InMux I__6865 (
            .O(N__40574),
            .I(N__40559));
    InMux I__6864 (
            .O(N__40573),
            .I(N__40555));
    InMux I__6863 (
            .O(N__40570),
            .I(N__40552));
    InMux I__6862 (
            .O(N__40569),
            .I(N__40549));
    InMux I__6861 (
            .O(N__40568),
            .I(N__40546));
    InMux I__6860 (
            .O(N__40567),
            .I(N__40537));
    CascadeMux I__6859 (
            .O(N__40566),
            .I(N__40532));
    InMux I__6858 (
            .O(N__40565),
            .I(N__40529));
    InMux I__6857 (
            .O(N__40564),
            .I(N__40519));
    InMux I__6856 (
            .O(N__40563),
            .I(N__40519));
    InMux I__6855 (
            .O(N__40562),
            .I(N__40519));
    LocalMux I__6854 (
            .O(N__40559),
            .I(N__40516));
    InMux I__6853 (
            .O(N__40558),
            .I(N__40513));
    LocalMux I__6852 (
            .O(N__40555),
            .I(N__40504));
    LocalMux I__6851 (
            .O(N__40552),
            .I(N__40504));
    LocalMux I__6850 (
            .O(N__40549),
            .I(N__40504));
    LocalMux I__6849 (
            .O(N__40546),
            .I(N__40504));
    InMux I__6848 (
            .O(N__40545),
            .I(N__40499));
    InMux I__6847 (
            .O(N__40544),
            .I(N__40499));
    InMux I__6846 (
            .O(N__40543),
            .I(N__40494));
    InMux I__6845 (
            .O(N__40542),
            .I(N__40494));
    InMux I__6844 (
            .O(N__40541),
            .I(N__40489));
    InMux I__6843 (
            .O(N__40540),
            .I(N__40489));
    LocalMux I__6842 (
            .O(N__40537),
            .I(N__40486));
    InMux I__6841 (
            .O(N__40536),
            .I(N__40480));
    InMux I__6840 (
            .O(N__40535),
            .I(N__40480));
    InMux I__6839 (
            .O(N__40532),
            .I(N__40476));
    LocalMux I__6838 (
            .O(N__40529),
            .I(N__40473));
    InMux I__6837 (
            .O(N__40528),
            .I(N__40468));
    InMux I__6836 (
            .O(N__40527),
            .I(N__40468));
    InMux I__6835 (
            .O(N__40526),
            .I(N__40464));
    LocalMux I__6834 (
            .O(N__40519),
            .I(N__40457));
    Span4Mux_v I__6833 (
            .O(N__40516),
            .I(N__40457));
    LocalMux I__6832 (
            .O(N__40513),
            .I(N__40457));
    Span4Mux_v I__6831 (
            .O(N__40504),
            .I(N__40452));
    LocalMux I__6830 (
            .O(N__40499),
            .I(N__40452));
    LocalMux I__6829 (
            .O(N__40494),
            .I(N__40447));
    LocalMux I__6828 (
            .O(N__40489),
            .I(N__40447));
    Span4Mux_h I__6827 (
            .O(N__40486),
            .I(N__40444));
    InMux I__6826 (
            .O(N__40485),
            .I(N__40441));
    LocalMux I__6825 (
            .O(N__40480),
            .I(N__40437));
    InMux I__6824 (
            .O(N__40479),
            .I(N__40434));
    LocalMux I__6823 (
            .O(N__40476),
            .I(N__40431));
    Span4Mux_v I__6822 (
            .O(N__40473),
            .I(N__40426));
    LocalMux I__6821 (
            .O(N__40468),
            .I(N__40426));
    InMux I__6820 (
            .O(N__40467),
            .I(N__40423));
    LocalMux I__6819 (
            .O(N__40464),
            .I(N__40420));
    Span4Mux_v I__6818 (
            .O(N__40457),
            .I(N__40417));
    Span4Mux_h I__6817 (
            .O(N__40452),
            .I(N__40414));
    Span4Mux_h I__6816 (
            .O(N__40447),
            .I(N__40402));
    Span4Mux_h I__6815 (
            .O(N__40444),
            .I(N__40402));
    LocalMux I__6814 (
            .O(N__40441),
            .I(N__40402));
    InMux I__6813 (
            .O(N__40440),
            .I(N__40399));
    Span4Mux_v I__6812 (
            .O(N__40437),
            .I(N__40396));
    LocalMux I__6811 (
            .O(N__40434),
            .I(N__40391));
    Span4Mux_v I__6810 (
            .O(N__40431),
            .I(N__40391));
    Span4Mux_h I__6809 (
            .O(N__40426),
            .I(N__40380));
    LocalMux I__6808 (
            .O(N__40423),
            .I(N__40380));
    Span4Mux_h I__6807 (
            .O(N__40420),
            .I(N__40380));
    Span4Mux_h I__6806 (
            .O(N__40417),
            .I(N__40380));
    Span4Mux_v I__6805 (
            .O(N__40414),
            .I(N__40380));
    InMux I__6804 (
            .O(N__40413),
            .I(N__40377));
    InMux I__6803 (
            .O(N__40412),
            .I(N__40374));
    InMux I__6802 (
            .O(N__40411),
            .I(N__40371));
    InMux I__6801 (
            .O(N__40410),
            .I(N__40368));
    InMux I__6800 (
            .O(N__40409),
            .I(N__40365));
    Span4Mux_v I__6799 (
            .O(N__40402),
            .I(N__40362));
    LocalMux I__6798 (
            .O(N__40399),
            .I(N__40355));
    Span4Mux_v I__6797 (
            .O(N__40396),
            .I(N__40355));
    Span4Mux_h I__6796 (
            .O(N__40391),
            .I(N__40355));
    Span4Mux_v I__6795 (
            .O(N__40380),
            .I(N__40352));
    LocalMux I__6794 (
            .O(N__40377),
            .I(count_enable_adj_4769));
    LocalMux I__6793 (
            .O(N__40374),
            .I(count_enable_adj_4769));
    LocalMux I__6792 (
            .O(N__40371),
            .I(count_enable_adj_4769));
    LocalMux I__6791 (
            .O(N__40368),
            .I(count_enable_adj_4769));
    LocalMux I__6790 (
            .O(N__40365),
            .I(count_enable_adj_4769));
    Odrv4 I__6789 (
            .O(N__40362),
            .I(count_enable_adj_4769));
    Odrv4 I__6788 (
            .O(N__40355),
            .I(count_enable_adj_4769));
    Odrv4 I__6787 (
            .O(N__40352),
            .I(count_enable_adj_4769));
    CascadeMux I__6786 (
            .O(N__40335),
            .I(N__40332));
    InMux I__6785 (
            .O(N__40332),
            .I(N__40328));
    InMux I__6784 (
            .O(N__40331),
            .I(N__40325));
    LocalMux I__6783 (
            .O(N__40328),
            .I(N__40321));
    LocalMux I__6782 (
            .O(N__40325),
            .I(N__40318));
    InMux I__6781 (
            .O(N__40324),
            .I(N__40315));
    Sp12to4 I__6780 (
            .O(N__40321),
            .I(N__40311));
    Span4Mux_v I__6779 (
            .O(N__40318),
            .I(N__40308));
    LocalMux I__6778 (
            .O(N__40315),
            .I(N__40305));
    InMux I__6777 (
            .O(N__40314),
            .I(N__40302));
    Span12Mux_h I__6776 (
            .O(N__40311),
            .I(N__40299));
    Span4Mux_h I__6775 (
            .O(N__40308),
            .I(N__40296));
    Span4Mux_v I__6774 (
            .O(N__40305),
            .I(N__40293));
    LocalMux I__6773 (
            .O(N__40302),
            .I(encoder1_position_31));
    Odrv12 I__6772 (
            .O(N__40299),
            .I(encoder1_position_31));
    Odrv4 I__6771 (
            .O(N__40296),
            .I(encoder1_position_31));
    Odrv4 I__6770 (
            .O(N__40293),
            .I(encoder1_position_31));
    InMux I__6769 (
            .O(N__40284),
            .I(N__40281));
    LocalMux I__6768 (
            .O(N__40281),
            .I(n2338));
    CascadeMux I__6767 (
            .O(N__40278),
            .I(N__40275));
    InMux I__6766 (
            .O(N__40275),
            .I(N__40271));
    InMux I__6765 (
            .O(N__40274),
            .I(N__40268));
    LocalMux I__6764 (
            .O(N__40271),
            .I(N__40261));
    LocalMux I__6763 (
            .O(N__40268),
            .I(N__40258));
    InMux I__6762 (
            .O(N__40267),
            .I(N__40255));
    InMux I__6761 (
            .O(N__40266),
            .I(N__40252));
    InMux I__6760 (
            .O(N__40265),
            .I(N__40249));
    InMux I__6759 (
            .O(N__40264),
            .I(N__40246));
    Span4Mux_h I__6758 (
            .O(N__40261),
            .I(N__40241));
    Span4Mux_h I__6757 (
            .O(N__40258),
            .I(N__40241));
    LocalMux I__6756 (
            .O(N__40255),
            .I(N__40236));
    LocalMux I__6755 (
            .O(N__40252),
            .I(N__40236));
    LocalMux I__6754 (
            .O(N__40249),
            .I(encoder1_position_21));
    LocalMux I__6753 (
            .O(N__40246),
            .I(encoder1_position_21));
    Odrv4 I__6752 (
            .O(N__40241),
            .I(encoder1_position_21));
    Odrv12 I__6751 (
            .O(N__40236),
            .I(encoder1_position_21));
    CascadeMux I__6750 (
            .O(N__40227),
            .I(N__40224));
    InMux I__6749 (
            .O(N__40224),
            .I(N__40221));
    LocalMux I__6748 (
            .O(N__40221),
            .I(N__40218));
    Span4Mux_v I__6747 (
            .O(N__40218),
            .I(N__40215));
    Sp12to4 I__6746 (
            .O(N__40215),
            .I(N__40210));
    InMux I__6745 (
            .O(N__40214),
            .I(N__40207));
    InMux I__6744 (
            .O(N__40213),
            .I(N__40201));
    Span12Mux_h I__6743 (
            .O(N__40210),
            .I(N__40196));
    LocalMux I__6742 (
            .O(N__40207),
            .I(N__40196));
    InMux I__6741 (
            .O(N__40206),
            .I(N__40193));
    InMux I__6740 (
            .O(N__40205),
            .I(N__40188));
    InMux I__6739 (
            .O(N__40204),
            .I(N__40188));
    LocalMux I__6738 (
            .O(N__40201),
            .I(encoder0_position_17));
    Odrv12 I__6737 (
            .O(N__40196),
            .I(encoder0_position_17));
    LocalMux I__6736 (
            .O(N__40193),
            .I(encoder0_position_17));
    LocalMux I__6735 (
            .O(N__40188),
            .I(encoder0_position_17));
    CascadeMux I__6734 (
            .O(N__40179),
            .I(N__40175));
    InMux I__6733 (
            .O(N__40178),
            .I(N__40171));
    InMux I__6732 (
            .O(N__40175),
            .I(N__40168));
    CascadeMux I__6731 (
            .O(N__40174),
            .I(N__40165));
    LocalMux I__6730 (
            .O(N__40171),
            .I(N__40162));
    LocalMux I__6729 (
            .O(N__40168),
            .I(N__40159));
    InMux I__6728 (
            .O(N__40165),
            .I(N__40156));
    Span4Mux_h I__6727 (
            .O(N__40162),
            .I(N__40153));
    Span4Mux_v I__6726 (
            .O(N__40159),
            .I(N__40148));
    LocalMux I__6725 (
            .O(N__40156),
            .I(N__40148));
    Span4Mux_h I__6724 (
            .O(N__40153),
            .I(N__40145));
    Span4Mux_v I__6723 (
            .O(N__40148),
            .I(N__40138));
    Span4Mux_h I__6722 (
            .O(N__40145),
            .I(N__40138));
    InMux I__6721 (
            .O(N__40144),
            .I(N__40133));
    InMux I__6720 (
            .O(N__40143),
            .I(N__40133));
    Odrv4 I__6719 (
            .O(N__40138),
            .I(encoder1_position_8));
    LocalMux I__6718 (
            .O(N__40133),
            .I(encoder1_position_8));
    InMux I__6717 (
            .O(N__40128),
            .I(N__40124));
    InMux I__6716 (
            .O(N__40127),
            .I(N__40121));
    LocalMux I__6715 (
            .O(N__40124),
            .I(N__40118));
    LocalMux I__6714 (
            .O(N__40121),
            .I(N__40115));
    Span4Mux_h I__6713 (
            .O(N__40118),
            .I(N__40112));
    Span4Mux_h I__6712 (
            .O(N__40115),
            .I(N__40109));
    Span4Mux_h I__6711 (
            .O(N__40112),
            .I(N__40106));
    Span4Mux_v I__6710 (
            .O(N__40109),
            .I(N__40103));
    Odrv4 I__6709 (
            .O(N__40106),
            .I(\c0.n22593 ));
    Odrv4 I__6708 (
            .O(N__40103),
            .I(\c0.n22593 ));
    CascadeMux I__6707 (
            .O(N__40098),
            .I(N__40095));
    InMux I__6706 (
            .O(N__40095),
            .I(N__40091));
    CascadeMux I__6705 (
            .O(N__40094),
            .I(N__40088));
    LocalMux I__6704 (
            .O(N__40091),
            .I(N__40085));
    InMux I__6703 (
            .O(N__40088),
            .I(N__40081));
    Span4Mux_v I__6702 (
            .O(N__40085),
            .I(N__40076));
    InMux I__6701 (
            .O(N__40084),
            .I(N__40073));
    LocalMux I__6700 (
            .O(N__40081),
            .I(N__40070));
    InMux I__6699 (
            .O(N__40080),
            .I(N__40065));
    InMux I__6698 (
            .O(N__40079),
            .I(N__40065));
    Span4Mux_h I__6697 (
            .O(N__40076),
            .I(N__40059));
    LocalMux I__6696 (
            .O(N__40073),
            .I(N__40059));
    Span4Mux_h I__6695 (
            .O(N__40070),
            .I(N__40054));
    LocalMux I__6694 (
            .O(N__40065),
            .I(N__40054));
    InMux I__6693 (
            .O(N__40064),
            .I(N__40051));
    Span4Mux_v I__6692 (
            .O(N__40059),
            .I(N__40048));
    Span4Mux_h I__6691 (
            .O(N__40054),
            .I(N__40045));
    LocalMux I__6690 (
            .O(N__40051),
            .I(encoder1_position_9));
    Odrv4 I__6689 (
            .O(N__40048),
            .I(encoder1_position_9));
    Odrv4 I__6688 (
            .O(N__40045),
            .I(encoder1_position_9));
    InMux I__6687 (
            .O(N__40038),
            .I(N__40035));
    LocalMux I__6686 (
            .O(N__40035),
            .I(\c0.n6_adj_4276 ));
    CascadeMux I__6685 (
            .O(N__40032),
            .I(N__40029));
    InMux I__6684 (
            .O(N__40029),
            .I(N__40026));
    LocalMux I__6683 (
            .O(N__40026),
            .I(N__40023));
    Span4Mux_v I__6682 (
            .O(N__40023),
            .I(N__40018));
    CascadeMux I__6681 (
            .O(N__40022),
            .I(N__40015));
    InMux I__6680 (
            .O(N__40021),
            .I(N__40012));
    Span4Mux_h I__6679 (
            .O(N__40018),
            .I(N__40009));
    InMux I__6678 (
            .O(N__40015),
            .I(N__40006));
    LocalMux I__6677 (
            .O(N__40012),
            .I(N__40003));
    Span4Mux_h I__6676 (
            .O(N__40009),
            .I(N__40000));
    LocalMux I__6675 (
            .O(N__40006),
            .I(N__39995));
    Span4Mux_v I__6674 (
            .O(N__40003),
            .I(N__39995));
    Odrv4 I__6673 (
            .O(N__40000),
            .I(\c0.n22372 ));
    Odrv4 I__6672 (
            .O(N__39995),
            .I(\c0.n22372 ));
    CascadeMux I__6671 (
            .O(N__39990),
            .I(N__39986));
    CascadeMux I__6670 (
            .O(N__39989),
            .I(N__39983));
    InMux I__6669 (
            .O(N__39986),
            .I(N__39979));
    InMux I__6668 (
            .O(N__39983),
            .I(N__39976));
    InMux I__6667 (
            .O(N__39982),
            .I(N__39973));
    LocalMux I__6666 (
            .O(N__39979),
            .I(N__39969));
    LocalMux I__6665 (
            .O(N__39976),
            .I(N__39966));
    LocalMux I__6664 (
            .O(N__39973),
            .I(N__39963));
    CascadeMux I__6663 (
            .O(N__39972),
            .I(N__39959));
    Span4Mux_h I__6662 (
            .O(N__39969),
            .I(N__39956));
    Span4Mux_h I__6661 (
            .O(N__39966),
            .I(N__39953));
    Span4Mux_h I__6660 (
            .O(N__39963),
            .I(N__39950));
    InMux I__6659 (
            .O(N__39962),
            .I(N__39947));
    InMux I__6658 (
            .O(N__39959),
            .I(N__39944));
    Span4Mux_v I__6657 (
            .O(N__39956),
            .I(N__39939));
    Span4Mux_v I__6656 (
            .O(N__39953),
            .I(N__39939));
    Span4Mux_v I__6655 (
            .O(N__39950),
            .I(N__39936));
    LocalMux I__6654 (
            .O(N__39947),
            .I(encoder1_position_28));
    LocalMux I__6653 (
            .O(N__39944),
            .I(encoder1_position_28));
    Odrv4 I__6652 (
            .O(N__39939),
            .I(encoder1_position_28));
    Odrv4 I__6651 (
            .O(N__39936),
            .I(encoder1_position_28));
    InMux I__6650 (
            .O(N__39927),
            .I(N__39924));
    LocalMux I__6649 (
            .O(N__39924),
            .I(N__39921));
    Span4Mux_v I__6648 (
            .O(N__39921),
            .I(N__39918));
    Odrv4 I__6647 (
            .O(N__39918),
            .I(\c0.n31_adj_4325 ));
    InMux I__6646 (
            .O(N__39915),
            .I(N__39911));
    InMux I__6645 (
            .O(N__39914),
            .I(N__39908));
    LocalMux I__6644 (
            .O(N__39911),
            .I(N__39905));
    LocalMux I__6643 (
            .O(N__39908),
            .I(N__39902));
    Span4Mux_h I__6642 (
            .O(N__39905),
            .I(N__39899));
    Span4Mux_h I__6641 (
            .O(N__39902),
            .I(N__39896));
    Odrv4 I__6640 (
            .O(N__39899),
            .I(\c0.n22775 ));
    Odrv4 I__6639 (
            .O(N__39896),
            .I(\c0.n22775 ));
    InMux I__6638 (
            .O(N__39891),
            .I(N__39888));
    LocalMux I__6637 (
            .O(N__39888),
            .I(n2348));
    InMux I__6636 (
            .O(N__39885),
            .I(N__39882));
    LocalMux I__6635 (
            .O(N__39882),
            .I(n2336));
    InMux I__6634 (
            .O(N__39879),
            .I(N__39876));
    LocalMux I__6633 (
            .O(N__39876),
            .I(N__39872));
    InMux I__6632 (
            .O(N__39875),
            .I(N__39869));
    Span4Mux_h I__6631 (
            .O(N__39872),
            .I(N__39864));
    LocalMux I__6630 (
            .O(N__39869),
            .I(N__39864));
    Odrv4 I__6629 (
            .O(N__39864),
            .I(\c0.n22608 ));
    CascadeMux I__6628 (
            .O(N__39861),
            .I(N__39858));
    InMux I__6627 (
            .O(N__39858),
            .I(N__39855));
    LocalMux I__6626 (
            .O(N__39855),
            .I(N__39852));
    Span4Mux_h I__6625 (
            .O(N__39852),
            .I(N__39849));
    Span4Mux_v I__6624 (
            .O(N__39849),
            .I(N__39845));
    InMux I__6623 (
            .O(N__39848),
            .I(N__39842));
    Span4Mux_v I__6622 (
            .O(N__39845),
            .I(N__39837));
    LocalMux I__6621 (
            .O(N__39842),
            .I(N__39832));
    InMux I__6620 (
            .O(N__39841),
            .I(N__39829));
    InMux I__6619 (
            .O(N__39840),
            .I(N__39826));
    Span4Mux_v I__6618 (
            .O(N__39837),
            .I(N__39823));
    InMux I__6617 (
            .O(N__39836),
            .I(N__39820));
    InMux I__6616 (
            .O(N__39835),
            .I(N__39817));
    Span4Mux_v I__6615 (
            .O(N__39832),
            .I(N__39814));
    LocalMux I__6614 (
            .O(N__39829),
            .I(N__39811));
    LocalMux I__6613 (
            .O(N__39826),
            .I(encoder0_position_2));
    Odrv4 I__6612 (
            .O(N__39823),
            .I(encoder0_position_2));
    LocalMux I__6611 (
            .O(N__39820),
            .I(encoder0_position_2));
    LocalMux I__6610 (
            .O(N__39817),
            .I(encoder0_position_2));
    Odrv4 I__6609 (
            .O(N__39814),
            .I(encoder0_position_2));
    Odrv4 I__6608 (
            .O(N__39811),
            .I(encoder0_position_2));
    InMux I__6607 (
            .O(N__39798),
            .I(N__39794));
    InMux I__6606 (
            .O(N__39797),
            .I(N__39791));
    LocalMux I__6605 (
            .O(N__39794),
            .I(N__39788));
    LocalMux I__6604 (
            .O(N__39791),
            .I(N__39785));
    Odrv4 I__6603 (
            .O(N__39788),
            .I(\c0.n22785 ));
    Odrv12 I__6602 (
            .O(N__39785),
            .I(\c0.n22785 ));
    InMux I__6601 (
            .O(N__39780),
            .I(N__39776));
    InMux I__6600 (
            .O(N__39779),
            .I(N__39773));
    LocalMux I__6599 (
            .O(N__39776),
            .I(N__39770));
    LocalMux I__6598 (
            .O(N__39773),
            .I(N__39767));
    Odrv4 I__6597 (
            .O(N__39770),
            .I(\c0.n13630 ));
    Odrv4 I__6596 (
            .O(N__39767),
            .I(\c0.n13630 ));
    InMux I__6595 (
            .O(N__39762),
            .I(N__39759));
    LocalMux I__6594 (
            .O(N__39759),
            .I(n2340));
    InMux I__6593 (
            .O(N__39756),
            .I(N__39751));
    InMux I__6592 (
            .O(N__39755),
            .I(N__39746));
    InMux I__6591 (
            .O(N__39754),
            .I(N__39746));
    LocalMux I__6590 (
            .O(N__39751),
            .I(N__39741));
    LocalMux I__6589 (
            .O(N__39746),
            .I(N__39738));
    InMux I__6588 (
            .O(N__39745),
            .I(N__39735));
    InMux I__6587 (
            .O(N__39744),
            .I(N__39732));
    Span4Mux_h I__6586 (
            .O(N__39741),
            .I(N__39729));
    Span4Mux_h I__6585 (
            .O(N__39738),
            .I(N__39726));
    LocalMux I__6584 (
            .O(N__39735),
            .I(\c0.FRAME_MATCHER_state_18 ));
    LocalMux I__6583 (
            .O(N__39732),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__6582 (
            .O(N__39729),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__6581 (
            .O(N__39726),
            .I(\c0.FRAME_MATCHER_state_18 ));
    SRMux I__6580 (
            .O(N__39717),
            .I(N__39714));
    LocalMux I__6579 (
            .O(N__39714),
            .I(N__39711));
    Span4Mux_h I__6578 (
            .O(N__39711),
            .I(N__39708));
    Odrv4 I__6577 (
            .O(N__39708),
            .I(\c0.n21639 ));
    CascadeMux I__6576 (
            .O(N__39705),
            .I(N__39701));
    InMux I__6575 (
            .O(N__39704),
            .I(N__39698));
    InMux I__6574 (
            .O(N__39701),
            .I(N__39695));
    LocalMux I__6573 (
            .O(N__39698),
            .I(N__39691));
    LocalMux I__6572 (
            .O(N__39695),
            .I(N__39688));
    InMux I__6571 (
            .O(N__39694),
            .I(N__39685));
    Span4Mux_v I__6570 (
            .O(N__39691),
            .I(N__39682));
    Span4Mux_h I__6569 (
            .O(N__39688),
            .I(N__39679));
    LocalMux I__6568 (
            .O(N__39685),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__6567 (
            .O(N__39682),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__6566 (
            .O(N__39679),
            .I(\c0.FRAME_MATCHER_state_12 ));
    SRMux I__6565 (
            .O(N__39672),
            .I(N__39669));
    LocalMux I__6564 (
            .O(N__39669),
            .I(N__39666));
    Span4Mux_h I__6563 (
            .O(N__39666),
            .I(N__39663));
    Span4Mux_v I__6562 (
            .O(N__39663),
            .I(N__39660));
    Odrv4 I__6561 (
            .O(N__39660),
            .I(\c0.n8_adj_4555 ));
    SRMux I__6560 (
            .O(N__39657),
            .I(N__39654));
    LocalMux I__6559 (
            .O(N__39654),
            .I(N__39651));
    Span4Mux_h I__6558 (
            .O(N__39651),
            .I(N__39648));
    Odrv4 I__6557 (
            .O(N__39648),
            .I(\c0.n21641 ));
    CascadeMux I__6556 (
            .O(N__39645),
            .I(N__39642));
    InMux I__6555 (
            .O(N__39642),
            .I(N__39639));
    LocalMux I__6554 (
            .O(N__39639),
            .I(N__39636));
    Span4Mux_v I__6553 (
            .O(N__39636),
            .I(N__39633));
    Span4Mux_h I__6552 (
            .O(N__39633),
            .I(N__39630));
    Span4Mux_v I__6551 (
            .O(N__39630),
            .I(N__39627));
    Span4Mux_v I__6550 (
            .O(N__39627),
            .I(N__39620));
    InMux I__6549 (
            .O(N__39626),
            .I(N__39617));
    InMux I__6548 (
            .O(N__39625),
            .I(N__39614));
    InMux I__6547 (
            .O(N__39624),
            .I(N__39609));
    InMux I__6546 (
            .O(N__39623),
            .I(N__39606));
    Span4Mux_h I__6545 (
            .O(N__39620),
            .I(N__39599));
    LocalMux I__6544 (
            .O(N__39617),
            .I(N__39599));
    LocalMux I__6543 (
            .O(N__39614),
            .I(N__39599));
    InMux I__6542 (
            .O(N__39613),
            .I(N__39596));
    InMux I__6541 (
            .O(N__39612),
            .I(N__39592));
    LocalMux I__6540 (
            .O(N__39609),
            .I(N__39589));
    LocalMux I__6539 (
            .O(N__39606),
            .I(N__39586));
    Span4Mux_v I__6538 (
            .O(N__39599),
            .I(N__39581));
    LocalMux I__6537 (
            .O(N__39596),
            .I(N__39581));
    InMux I__6536 (
            .O(N__39595),
            .I(N__39578));
    LocalMux I__6535 (
            .O(N__39592),
            .I(encoder0_position_30));
    Odrv12 I__6534 (
            .O(N__39589),
            .I(encoder0_position_30));
    Odrv4 I__6533 (
            .O(N__39586),
            .I(encoder0_position_30));
    Odrv4 I__6532 (
            .O(N__39581),
            .I(encoder0_position_30));
    LocalMux I__6531 (
            .O(N__39578),
            .I(encoder0_position_30));
    InMux I__6530 (
            .O(N__39567),
            .I(N__39564));
    LocalMux I__6529 (
            .O(N__39564),
            .I(N__39561));
    Odrv4 I__6528 (
            .O(N__39561),
            .I(n2342));
    InMux I__6527 (
            .O(N__39558),
            .I(N__39555));
    LocalMux I__6526 (
            .O(N__39555),
            .I(N__39550));
    InMux I__6525 (
            .O(N__39554),
            .I(N__39546));
    InMux I__6524 (
            .O(N__39553),
            .I(N__39543));
    Sp12to4 I__6523 (
            .O(N__39550),
            .I(N__39539));
    InMux I__6522 (
            .O(N__39549),
            .I(N__39536));
    LocalMux I__6521 (
            .O(N__39546),
            .I(N__39533));
    LocalMux I__6520 (
            .O(N__39543),
            .I(N__39530));
    InMux I__6519 (
            .O(N__39542),
            .I(N__39526));
    Span12Mux_v I__6518 (
            .O(N__39539),
            .I(N__39521));
    LocalMux I__6517 (
            .O(N__39536),
            .I(N__39521));
    Span4Mux_v I__6516 (
            .O(N__39533),
            .I(N__39516));
    Span4Mux_h I__6515 (
            .O(N__39530),
            .I(N__39516));
    InMux I__6514 (
            .O(N__39529),
            .I(N__39513));
    LocalMux I__6513 (
            .O(N__39526),
            .I(encoder0_position_15));
    Odrv12 I__6512 (
            .O(N__39521),
            .I(encoder0_position_15));
    Odrv4 I__6511 (
            .O(N__39516),
            .I(encoder0_position_15));
    LocalMux I__6510 (
            .O(N__39513),
            .I(encoder0_position_15));
    InMux I__6509 (
            .O(N__39504),
            .I(N__39501));
    LocalMux I__6508 (
            .O(N__39501),
            .I(n2352));
    CascadeMux I__6507 (
            .O(N__39498),
            .I(\c0.n30_adj_4730_cascade_ ));
    InMux I__6506 (
            .O(N__39495),
            .I(N__39492));
    LocalMux I__6505 (
            .O(N__39492),
            .I(N__39489));
    Span4Mux_h I__6504 (
            .O(N__39489),
            .I(N__39485));
    InMux I__6503 (
            .O(N__39488),
            .I(N__39482));
    Span4Mux_v I__6502 (
            .O(N__39485),
            .I(N__39479));
    LocalMux I__6501 (
            .O(N__39482),
            .I(N__39476));
    Span4Mux_v I__6500 (
            .O(N__39479),
            .I(N__39473));
    Span12Mux_v I__6499 (
            .O(N__39476),
            .I(N__39470));
    Odrv4 I__6498 (
            .O(N__39473),
            .I(\c0.n17539 ));
    Odrv12 I__6497 (
            .O(N__39470),
            .I(\c0.n17539 ));
    InMux I__6496 (
            .O(N__39465),
            .I(N__39462));
    LocalMux I__6495 (
            .O(N__39462),
            .I(N__39459));
    Span4Mux_v I__6494 (
            .O(N__39459),
            .I(N__39455));
    CascadeMux I__6493 (
            .O(N__39458),
            .I(N__39452));
    Span4Mux_h I__6492 (
            .O(N__39455),
            .I(N__39448));
    InMux I__6491 (
            .O(N__39452),
            .I(N__39445));
    InMux I__6490 (
            .O(N__39451),
            .I(N__39442));
    Span4Mux_v I__6489 (
            .O(N__39448),
            .I(N__39434));
    LocalMux I__6488 (
            .O(N__39445),
            .I(N__39434));
    LocalMux I__6487 (
            .O(N__39442),
            .I(N__39434));
    InMux I__6486 (
            .O(N__39441),
            .I(N__39431));
    Span4Mux_v I__6485 (
            .O(N__39434),
            .I(N__39428));
    LocalMux I__6484 (
            .O(N__39431),
            .I(\c0.n17846 ));
    Odrv4 I__6483 (
            .O(N__39428),
            .I(\c0.n17846 ));
    InMux I__6482 (
            .O(N__39423),
            .I(N__39418));
    InMux I__6481 (
            .O(N__39422),
            .I(N__39413));
    InMux I__6480 (
            .O(N__39421),
            .I(N__39413));
    LocalMux I__6479 (
            .O(N__39418),
            .I(N__39407));
    LocalMux I__6478 (
            .O(N__39413),
            .I(N__39407));
    InMux I__6477 (
            .O(N__39412),
            .I(N__39404));
    Odrv4 I__6476 (
            .O(N__39407),
            .I(\c0.n4_adj_4654 ));
    LocalMux I__6475 (
            .O(N__39404),
            .I(\c0.n4_adj_4654 ));
    CascadeMux I__6474 (
            .O(N__39399),
            .I(N__39396));
    InMux I__6473 (
            .O(N__39396),
            .I(N__39393));
    LocalMux I__6472 (
            .O(N__39393),
            .I(N__39389));
    CascadeMux I__6471 (
            .O(N__39392),
            .I(N__39386));
    Span4Mux_h I__6470 (
            .O(N__39389),
            .I(N__39383));
    InMux I__6469 (
            .O(N__39386),
            .I(N__39380));
    Odrv4 I__6468 (
            .O(N__39383),
            .I(\c0.n17533 ));
    LocalMux I__6467 (
            .O(N__39380),
            .I(\c0.n17533 ));
    InMux I__6466 (
            .O(N__39375),
            .I(N__39372));
    LocalMux I__6465 (
            .O(N__39372),
            .I(N__39367));
    InMux I__6464 (
            .O(N__39371),
            .I(N__39364));
    InMux I__6463 (
            .O(N__39370),
            .I(N__39361));
    Span4Mux_h I__6462 (
            .O(N__39367),
            .I(N__39358));
    LocalMux I__6461 (
            .O(N__39364),
            .I(N__39353));
    LocalMux I__6460 (
            .O(N__39361),
            .I(N__39353));
    Odrv4 I__6459 (
            .O(N__39358),
            .I(\c0.n22907 ));
    Odrv12 I__6458 (
            .O(N__39353),
            .I(\c0.n22907 ));
    InMux I__6457 (
            .O(N__39348),
            .I(N__39345));
    LocalMux I__6456 (
            .O(N__39345),
            .I(N__39342));
    Odrv4 I__6455 (
            .O(N__39342),
            .I(\c0.n24422 ));
    CascadeMux I__6454 (
            .O(N__39339),
            .I(\c0.n24596_cascade_ ));
    InMux I__6453 (
            .O(N__39336),
            .I(N__39330));
    InMux I__6452 (
            .O(N__39335),
            .I(N__39327));
    InMux I__6451 (
            .O(N__39334),
            .I(N__39322));
    InMux I__6450 (
            .O(N__39333),
            .I(N__39322));
    LocalMux I__6449 (
            .O(N__39330),
            .I(\c0.n2004 ));
    LocalMux I__6448 (
            .O(N__39327),
            .I(\c0.n2004 ));
    LocalMux I__6447 (
            .O(N__39322),
            .I(\c0.n2004 ));
    InMux I__6446 (
            .O(N__39315),
            .I(N__39311));
    InMux I__6445 (
            .O(N__39314),
            .I(N__39308));
    LocalMux I__6444 (
            .O(N__39311),
            .I(N__39305));
    LocalMux I__6443 (
            .O(N__39308),
            .I(N__39302));
    Span12Mux_s10_h I__6442 (
            .O(N__39305),
            .I(N__39297));
    Span4Mux_h I__6441 (
            .O(N__39302),
            .I(N__39294));
    InMux I__6440 (
            .O(N__39301),
            .I(N__39289));
    InMux I__6439 (
            .O(N__39300),
            .I(N__39289));
    Odrv12 I__6438 (
            .O(N__39297),
            .I(\c0.rx.r_SM_Main_2_N_3686_0 ));
    Odrv4 I__6437 (
            .O(N__39294),
            .I(\c0.rx.r_SM_Main_2_N_3686_0 ));
    LocalMux I__6436 (
            .O(N__39289),
            .I(\c0.rx.r_SM_Main_2_N_3686_0 ));
    CascadeMux I__6435 (
            .O(N__39282),
            .I(\c0.rx.n6_cascade_ ));
    CEMux I__6434 (
            .O(N__39279),
            .I(N__39276));
    LocalMux I__6433 (
            .O(N__39276),
            .I(N__39272));
    InMux I__6432 (
            .O(N__39275),
            .I(N__39269));
    Span12Mux_h I__6431 (
            .O(N__39272),
            .I(N__39266));
    LocalMux I__6430 (
            .O(N__39269),
            .I(N__39263));
    Odrv12 I__6429 (
            .O(N__39266),
            .I(n14439));
    Odrv12 I__6428 (
            .O(N__39263),
            .I(n14439));
    InMux I__6427 (
            .O(N__39258),
            .I(N__39254));
    InMux I__6426 (
            .O(N__39257),
            .I(N__39251));
    LocalMux I__6425 (
            .O(N__39254),
            .I(N__39247));
    LocalMux I__6424 (
            .O(N__39251),
            .I(N__39244));
    InMux I__6423 (
            .O(N__39250),
            .I(N__39241));
    Span4Mux_v I__6422 (
            .O(N__39247),
            .I(N__39237));
    Span4Mux_h I__6421 (
            .O(N__39244),
            .I(N__39234));
    LocalMux I__6420 (
            .O(N__39241),
            .I(N__39231));
    InMux I__6419 (
            .O(N__39240),
            .I(N__39228));
    Odrv4 I__6418 (
            .O(N__39237),
            .I(\c0.n7570 ));
    Odrv4 I__6417 (
            .O(N__39234),
            .I(\c0.n7570 ));
    Odrv12 I__6416 (
            .O(N__39231),
            .I(\c0.n7570 ));
    LocalMux I__6415 (
            .O(N__39228),
            .I(\c0.n7570 ));
    InMux I__6414 (
            .O(N__39219),
            .I(N__39216));
    LocalMux I__6413 (
            .O(N__39216),
            .I(N__39213));
    Odrv4 I__6412 (
            .O(N__39213),
            .I(\c0.n24386 ));
    CascadeMux I__6411 (
            .O(N__39210),
            .I(\c0.n24302_cascade_ ));
    InMux I__6410 (
            .O(N__39207),
            .I(N__39203));
    InMux I__6409 (
            .O(N__39206),
            .I(N__39199));
    LocalMux I__6408 (
            .O(N__39203),
            .I(N__39196));
    InMux I__6407 (
            .O(N__39202),
            .I(N__39193));
    LocalMux I__6406 (
            .O(N__39199),
            .I(\c0.FRAME_MATCHER_state_10 ));
    Odrv4 I__6405 (
            .O(N__39196),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__6404 (
            .O(N__39193),
            .I(\c0.FRAME_MATCHER_state_10 ));
    SRMux I__6403 (
            .O(N__39186),
            .I(N__39183));
    LocalMux I__6402 (
            .O(N__39183),
            .I(N__39180));
    Span4Mux_h I__6401 (
            .O(N__39180),
            .I(N__39177));
    Span4Mux_h I__6400 (
            .O(N__39177),
            .I(N__39174));
    Odrv4 I__6399 (
            .O(N__39174),
            .I(\c0.n8_adj_4556 ));
    InMux I__6398 (
            .O(N__39171),
            .I(N__39165));
    InMux I__6397 (
            .O(N__39170),
            .I(N__39162));
    InMux I__6396 (
            .O(N__39169),
            .I(N__39157));
    InMux I__6395 (
            .O(N__39168),
            .I(N__39157));
    LocalMux I__6394 (
            .O(N__39165),
            .I(N__39154));
    LocalMux I__6393 (
            .O(N__39162),
            .I(N__39151));
    LocalMux I__6392 (
            .O(N__39157),
            .I(data_in_3_5));
    Odrv4 I__6391 (
            .O(N__39154),
            .I(data_in_3_5));
    Odrv12 I__6390 (
            .O(N__39151),
            .I(data_in_3_5));
    InMux I__6389 (
            .O(N__39144),
            .I(N__39140));
    InMux I__6388 (
            .O(N__39143),
            .I(N__39137));
    LocalMux I__6387 (
            .O(N__39140),
            .I(N__39134));
    LocalMux I__6386 (
            .O(N__39137),
            .I(N__39129));
    Span4Mux_v I__6385 (
            .O(N__39134),
            .I(N__39129));
    Span4Mux_h I__6384 (
            .O(N__39129),
            .I(N__39126));
    Odrv4 I__6383 (
            .O(N__39126),
            .I(\c0.n13063 ));
    CascadeMux I__6382 (
            .O(N__39123),
            .I(\c0.n13063_cascade_ ));
    InMux I__6381 (
            .O(N__39120),
            .I(N__39117));
    LocalMux I__6380 (
            .O(N__39117),
            .I(\c0.n6_adj_4263 ));
    InMux I__6379 (
            .O(N__39114),
            .I(N__39103));
    InMux I__6378 (
            .O(N__39113),
            .I(N__39103));
    InMux I__6377 (
            .O(N__39112),
            .I(N__39098));
    InMux I__6376 (
            .O(N__39111),
            .I(N__39098));
    InMux I__6375 (
            .O(N__39110),
            .I(N__39094));
    InMux I__6374 (
            .O(N__39109),
            .I(N__39091));
    InMux I__6373 (
            .O(N__39108),
            .I(N__39085));
    LocalMux I__6372 (
            .O(N__39103),
            .I(N__39080));
    LocalMux I__6371 (
            .O(N__39098),
            .I(N__39080));
    InMux I__6370 (
            .O(N__39097),
            .I(N__39077));
    LocalMux I__6369 (
            .O(N__39094),
            .I(N__39072));
    LocalMux I__6368 (
            .O(N__39091),
            .I(N__39072));
    InMux I__6367 (
            .O(N__39090),
            .I(N__39068));
    InMux I__6366 (
            .O(N__39089),
            .I(N__39063));
    InMux I__6365 (
            .O(N__39088),
            .I(N__39063));
    LocalMux I__6364 (
            .O(N__39085),
            .I(N__39056));
    Span4Mux_v I__6363 (
            .O(N__39080),
            .I(N__39056));
    LocalMux I__6362 (
            .O(N__39077),
            .I(N__39056));
    Span4Mux_h I__6361 (
            .O(N__39072),
            .I(N__39053));
    InMux I__6360 (
            .O(N__39071),
            .I(N__39050));
    LocalMux I__6359 (
            .O(N__39068),
            .I(\c0.n9706 ));
    LocalMux I__6358 (
            .O(N__39063),
            .I(\c0.n9706 ));
    Odrv4 I__6357 (
            .O(N__39056),
            .I(\c0.n9706 ));
    Odrv4 I__6356 (
            .O(N__39053),
            .I(\c0.n9706 ));
    LocalMux I__6355 (
            .O(N__39050),
            .I(\c0.n9706 ));
    InMux I__6354 (
            .O(N__39039),
            .I(N__39035));
    InMux I__6353 (
            .O(N__39038),
            .I(N__39032));
    LocalMux I__6352 (
            .O(N__39035),
            .I(N__39029));
    LocalMux I__6351 (
            .O(N__39032),
            .I(N__39026));
    Span4Mux_v I__6350 (
            .O(N__39029),
            .I(N__39021));
    Span4Mux_v I__6349 (
            .O(N__39026),
            .I(N__39021));
    Span4Mux_h I__6348 (
            .O(N__39021),
            .I(N__39017));
    InMux I__6347 (
            .O(N__39020),
            .I(N__39014));
    Odrv4 I__6346 (
            .O(N__39017),
            .I(\c0.n3325 ));
    LocalMux I__6345 (
            .O(N__39014),
            .I(\c0.n3325 ));
    InMux I__6344 (
            .O(N__39009),
            .I(N__39004));
    InMux I__6343 (
            .O(N__39008),
            .I(N__39001));
    InMux I__6342 (
            .O(N__39007),
            .I(N__38998));
    LocalMux I__6341 (
            .O(N__39004),
            .I(N__38995));
    LocalMux I__6340 (
            .O(N__39001),
            .I(data_in_2_7));
    LocalMux I__6339 (
            .O(N__38998),
            .I(data_in_2_7));
    Odrv12 I__6338 (
            .O(N__38995),
            .I(data_in_2_7));
    InMux I__6337 (
            .O(N__38988),
            .I(N__38982));
    InMux I__6336 (
            .O(N__38987),
            .I(N__38982));
    LocalMux I__6335 (
            .O(N__38982),
            .I(N__38978));
    InMux I__6334 (
            .O(N__38981),
            .I(N__38975));
    Sp12to4 I__6333 (
            .O(N__38978),
            .I(N__38972));
    LocalMux I__6332 (
            .O(N__38975),
            .I(data_in_1_7));
    Odrv12 I__6331 (
            .O(N__38972),
            .I(data_in_1_7));
    InMux I__6330 (
            .O(N__38967),
            .I(N__38961));
    InMux I__6329 (
            .O(N__38966),
            .I(N__38961));
    LocalMux I__6328 (
            .O(N__38961),
            .I(N__38958));
    Odrv4 I__6327 (
            .O(N__38958),
            .I(\c0.n17682 ));
    InMux I__6326 (
            .O(N__38955),
            .I(N__38948));
    InMux I__6325 (
            .O(N__38954),
            .I(N__38935));
    InMux I__6324 (
            .O(N__38953),
            .I(N__38935));
    InMux I__6323 (
            .O(N__38952),
            .I(N__38935));
    InMux I__6322 (
            .O(N__38951),
            .I(N__38935));
    LocalMux I__6321 (
            .O(N__38948),
            .I(N__38930));
    InMux I__6320 (
            .O(N__38947),
            .I(N__38921));
    InMux I__6319 (
            .O(N__38946),
            .I(N__38921));
    InMux I__6318 (
            .O(N__38945),
            .I(N__38921));
    InMux I__6317 (
            .O(N__38944),
            .I(N__38921));
    LocalMux I__6316 (
            .O(N__38935),
            .I(N__38918));
    InMux I__6315 (
            .O(N__38934),
            .I(N__38915));
    InMux I__6314 (
            .O(N__38933),
            .I(N__38910));
    Span4Mux_v I__6313 (
            .O(N__38930),
            .I(N__38905));
    LocalMux I__6312 (
            .O(N__38921),
            .I(N__38905));
    Span4Mux_h I__6311 (
            .O(N__38918),
            .I(N__38900));
    LocalMux I__6310 (
            .O(N__38915),
            .I(N__38900));
    InMux I__6309 (
            .O(N__38914),
            .I(N__38895));
    InMux I__6308 (
            .O(N__38913),
            .I(N__38895));
    LocalMux I__6307 (
            .O(N__38910),
            .I(\c0.n1 ));
    Odrv4 I__6306 (
            .O(N__38905),
            .I(\c0.n1 ));
    Odrv4 I__6305 (
            .O(N__38900),
            .I(\c0.n1 ));
    LocalMux I__6304 (
            .O(N__38895),
            .I(\c0.n1 ));
    InMux I__6303 (
            .O(N__38886),
            .I(N__38883));
    LocalMux I__6302 (
            .O(N__38883),
            .I(\c0.n24745 ));
    CascadeMux I__6301 (
            .O(N__38880),
            .I(N__38876));
    InMux I__6300 (
            .O(N__38879),
            .I(N__38872));
    InMux I__6299 (
            .O(N__38876),
            .I(N__38869));
    InMux I__6298 (
            .O(N__38875),
            .I(N__38865));
    LocalMux I__6297 (
            .O(N__38872),
            .I(N__38860));
    LocalMux I__6296 (
            .O(N__38869),
            .I(N__38860));
    InMux I__6295 (
            .O(N__38868),
            .I(N__38857));
    LocalMux I__6294 (
            .O(N__38865),
            .I(N__38852));
    Span4Mux_v I__6293 (
            .O(N__38860),
            .I(N__38852));
    LocalMux I__6292 (
            .O(N__38857),
            .I(data_in_2_6));
    Odrv4 I__6291 (
            .O(N__38852),
            .I(data_in_2_6));
    InMux I__6290 (
            .O(N__38847),
            .I(N__38842));
    InMux I__6289 (
            .O(N__38846),
            .I(N__38839));
    InMux I__6288 (
            .O(N__38845),
            .I(N__38836));
    LocalMux I__6287 (
            .O(N__38842),
            .I(data_in_0_5));
    LocalMux I__6286 (
            .O(N__38839),
            .I(data_in_0_5));
    LocalMux I__6285 (
            .O(N__38836),
            .I(data_in_0_5));
    InMux I__6284 (
            .O(N__38829),
            .I(N__38826));
    LocalMux I__6283 (
            .O(N__38826),
            .I(\c0.n17_adj_4232 ));
    InMux I__6282 (
            .O(N__38823),
            .I(N__38820));
    LocalMux I__6281 (
            .O(N__38820),
            .I(N__38817));
    Span4Mux_v I__6280 (
            .O(N__38817),
            .I(N__38814));
    Odrv4 I__6279 (
            .O(N__38814),
            .I(n2261));
    CascadeMux I__6278 (
            .O(N__38811),
            .I(N__38805));
    InMux I__6277 (
            .O(N__38810),
            .I(N__38802));
    InMux I__6276 (
            .O(N__38809),
            .I(N__38799));
    InMux I__6275 (
            .O(N__38808),
            .I(N__38796));
    InMux I__6274 (
            .O(N__38805),
            .I(N__38793));
    LocalMux I__6273 (
            .O(N__38802),
            .I(N__38788));
    LocalMux I__6272 (
            .O(N__38799),
            .I(N__38788));
    LocalMux I__6271 (
            .O(N__38796),
            .I(N__38782));
    LocalMux I__6270 (
            .O(N__38793),
            .I(N__38782));
    Span12Mux_h I__6269 (
            .O(N__38788),
            .I(N__38779));
    InMux I__6268 (
            .O(N__38787),
            .I(N__38776));
    Span4Mux_h I__6267 (
            .O(N__38782),
            .I(N__38773));
    Span12Mux_v I__6266 (
            .O(N__38779),
            .I(N__38770));
    LocalMux I__6265 (
            .O(N__38776),
            .I(encoder1_position_30));
    Odrv4 I__6264 (
            .O(N__38773),
            .I(encoder1_position_30));
    Odrv12 I__6263 (
            .O(N__38770),
            .I(encoder1_position_30));
    InMux I__6262 (
            .O(N__38763),
            .I(N__38758));
    CascadeMux I__6261 (
            .O(N__38762),
            .I(N__38755));
    InMux I__6260 (
            .O(N__38761),
            .I(N__38751));
    LocalMux I__6259 (
            .O(N__38758),
            .I(N__38748));
    InMux I__6258 (
            .O(N__38755),
            .I(N__38743));
    InMux I__6257 (
            .O(N__38754),
            .I(N__38743));
    LocalMux I__6256 (
            .O(N__38751),
            .I(data_in_3_7));
    Odrv4 I__6255 (
            .O(N__38748),
            .I(data_in_3_7));
    LocalMux I__6254 (
            .O(N__38743),
            .I(data_in_3_7));
    InMux I__6253 (
            .O(N__38736),
            .I(N__38731));
    InMux I__6252 (
            .O(N__38735),
            .I(N__38728));
    InMux I__6251 (
            .O(N__38734),
            .I(N__38725));
    LocalMux I__6250 (
            .O(N__38731),
            .I(N__38722));
    LocalMux I__6249 (
            .O(N__38728),
            .I(N__38719));
    LocalMux I__6248 (
            .O(N__38725),
            .I(N__38713));
    Span4Mux_h I__6247 (
            .O(N__38722),
            .I(N__38713));
    Span4Mux_h I__6246 (
            .O(N__38719),
            .I(N__38710));
    InMux I__6245 (
            .O(N__38718),
            .I(N__38707));
    Span4Mux_v I__6244 (
            .O(N__38713),
            .I(N__38704));
    Odrv4 I__6243 (
            .O(N__38710),
            .I(data_in_2_2));
    LocalMux I__6242 (
            .O(N__38707),
            .I(data_in_2_2));
    Odrv4 I__6241 (
            .O(N__38704),
            .I(data_in_2_2));
    CascadeMux I__6240 (
            .O(N__38697),
            .I(N__38694));
    InMux I__6239 (
            .O(N__38694),
            .I(N__38688));
    InMux I__6238 (
            .O(N__38693),
            .I(N__38688));
    LocalMux I__6237 (
            .O(N__38688),
            .I(data_out_frame_8_1));
    CascadeMux I__6236 (
            .O(N__38685),
            .I(N__38682));
    InMux I__6235 (
            .O(N__38682),
            .I(N__38679));
    LocalMux I__6234 (
            .O(N__38679),
            .I(N__38676));
    Span4Mux_h I__6233 (
            .O(N__38676),
            .I(N__38670));
    InMux I__6232 (
            .O(N__38675),
            .I(N__38667));
    InMux I__6231 (
            .O(N__38674),
            .I(N__38664));
    InMux I__6230 (
            .O(N__38673),
            .I(N__38661));
    Span4Mux_v I__6229 (
            .O(N__38670),
            .I(N__38658));
    LocalMux I__6228 (
            .O(N__38667),
            .I(encoder1_position_29));
    LocalMux I__6227 (
            .O(N__38664),
            .I(encoder1_position_29));
    LocalMux I__6226 (
            .O(N__38661),
            .I(encoder1_position_29));
    Odrv4 I__6225 (
            .O(N__38658),
            .I(encoder1_position_29));
    CascadeMux I__6224 (
            .O(N__38649),
            .I(N__38645));
    InMux I__6223 (
            .O(N__38648),
            .I(N__38642));
    InMux I__6222 (
            .O(N__38645),
            .I(N__38639));
    LocalMux I__6221 (
            .O(N__38642),
            .I(N__38636));
    LocalMux I__6220 (
            .O(N__38639),
            .I(data_out_frame_10_5));
    Odrv12 I__6219 (
            .O(N__38636),
            .I(data_out_frame_10_5));
    InMux I__6218 (
            .O(N__38631),
            .I(N__38627));
    InMux I__6217 (
            .O(N__38630),
            .I(N__38624));
    LocalMux I__6216 (
            .O(N__38627),
            .I(N__38619));
    LocalMux I__6215 (
            .O(N__38624),
            .I(N__38619));
    Odrv12 I__6214 (
            .O(N__38619),
            .I(\c0.n13046 ));
    InMux I__6213 (
            .O(N__38616),
            .I(N__38613));
    LocalMux I__6212 (
            .O(N__38613),
            .I(N__38609));
    InMux I__6211 (
            .O(N__38612),
            .I(N__38606));
    Span4Mux_v I__6210 (
            .O(N__38609),
            .I(N__38601));
    LocalMux I__6209 (
            .O(N__38606),
            .I(N__38601));
    Odrv4 I__6208 (
            .O(N__38601),
            .I(\c0.n12898 ));
    CascadeMux I__6207 (
            .O(N__38598),
            .I(\c0.n20_adj_4308_cascade_ ));
    InMux I__6206 (
            .O(N__38595),
            .I(N__38592));
    LocalMux I__6205 (
            .O(N__38592),
            .I(\c0.n19_adj_4307 ));
    CascadeMux I__6204 (
            .O(N__38589),
            .I(\c0.n16_adj_4231_cascade_ ));
    CascadeMux I__6203 (
            .O(N__38586),
            .I(N__38582));
    InMux I__6202 (
            .O(N__38585),
            .I(N__38579));
    InMux I__6201 (
            .O(N__38582),
            .I(N__38576));
    LocalMux I__6200 (
            .O(N__38579),
            .I(N__38571));
    LocalMux I__6199 (
            .O(N__38576),
            .I(N__38571));
    Odrv12 I__6198 (
            .O(N__38571),
            .I(\c0.n12986 ));
    InMux I__6197 (
            .O(N__38568),
            .I(N__38565));
    LocalMux I__6196 (
            .O(N__38565),
            .I(\c0.n17_adj_4234 ));
    InMux I__6195 (
            .O(N__38562),
            .I(N__38559));
    LocalMux I__6194 (
            .O(N__38559),
            .I(N__38556));
    Odrv4 I__6193 (
            .O(N__38556),
            .I(n2268));
    CascadeMux I__6192 (
            .O(N__38553),
            .I(N__38548));
    InMux I__6191 (
            .O(N__38552),
            .I(N__38543));
    InMux I__6190 (
            .O(N__38551),
            .I(N__38543));
    InMux I__6189 (
            .O(N__38548),
            .I(N__38539));
    LocalMux I__6188 (
            .O(N__38543),
            .I(N__38536));
    InMux I__6187 (
            .O(N__38542),
            .I(N__38532));
    LocalMux I__6186 (
            .O(N__38539),
            .I(N__38529));
    Span4Mux_h I__6185 (
            .O(N__38536),
            .I(N__38526));
    InMux I__6184 (
            .O(N__38535),
            .I(N__38523));
    LocalMux I__6183 (
            .O(N__38532),
            .I(N__38520));
    Span4Mux_v I__6182 (
            .O(N__38529),
            .I(N__38515));
    Span4Mux_v I__6181 (
            .O(N__38526),
            .I(N__38515));
    LocalMux I__6180 (
            .O(N__38523),
            .I(encoder1_position_23));
    Odrv4 I__6179 (
            .O(N__38520),
            .I(encoder1_position_23));
    Odrv4 I__6178 (
            .O(N__38515),
            .I(encoder1_position_23));
    InMux I__6177 (
            .O(N__38508),
            .I(N__38505));
    LocalMux I__6176 (
            .O(N__38505),
            .I(N__38502));
    Span4Mux_v I__6175 (
            .O(N__38502),
            .I(N__38499));
    Span4Mux_v I__6174 (
            .O(N__38499),
            .I(N__38496));
    Odrv4 I__6173 (
            .O(N__38496),
            .I(n2344));
    InMux I__6172 (
            .O(N__38493),
            .I(N__38490));
    LocalMux I__6171 (
            .O(N__38490),
            .I(N__38487));
    Odrv12 I__6170 (
            .O(N__38487),
            .I(\c0.n10_adj_4240 ));
    CEMux I__6169 (
            .O(N__38484),
            .I(N__38479));
    CEMux I__6168 (
            .O(N__38483),
            .I(N__38475));
    InMux I__6167 (
            .O(N__38482),
            .I(N__38472));
    LocalMux I__6166 (
            .O(N__38479),
            .I(N__38468));
    CascadeMux I__6165 (
            .O(N__38478),
            .I(N__38464));
    LocalMux I__6164 (
            .O(N__38475),
            .I(N__38460));
    LocalMux I__6163 (
            .O(N__38472),
            .I(N__38457));
    InMux I__6162 (
            .O(N__38471),
            .I(N__38454));
    Span4Mux_v I__6161 (
            .O(N__38468),
            .I(N__38451));
    InMux I__6160 (
            .O(N__38467),
            .I(N__38446));
    InMux I__6159 (
            .O(N__38464),
            .I(N__38446));
    InMux I__6158 (
            .O(N__38463),
            .I(N__38443));
    Span4Mux_v I__6157 (
            .O(N__38460),
            .I(N__38438));
    Span4Mux_v I__6156 (
            .O(N__38457),
            .I(N__38438));
    LocalMux I__6155 (
            .O(N__38454),
            .I(N__38435));
    Span4Mux_h I__6154 (
            .O(N__38451),
            .I(N__38430));
    LocalMux I__6153 (
            .O(N__38446),
            .I(N__38430));
    LocalMux I__6152 (
            .O(N__38443),
            .I(N__38427));
    Span4Mux_h I__6151 (
            .O(N__38438),
            .I(N__38420));
    Span4Mux_v I__6150 (
            .O(N__38435),
            .I(N__38420));
    Span4Mux_v I__6149 (
            .O(N__38430),
            .I(N__38420));
    Odrv4 I__6148 (
            .O(N__38427),
            .I(n14374));
    Odrv4 I__6147 (
            .O(N__38420),
            .I(n14374));
    InMux I__6146 (
            .O(N__38415),
            .I(N__38412));
    LocalMux I__6145 (
            .O(N__38412),
            .I(N__38409));
    Span4Mux_h I__6144 (
            .O(N__38409),
            .I(N__38406));
    Span4Mux_h I__6143 (
            .O(N__38406),
            .I(N__38403));
    Odrv4 I__6142 (
            .O(N__38403),
            .I(\c0.tx.n24889 ));
    InMux I__6141 (
            .O(N__38400),
            .I(N__38397));
    LocalMux I__6140 (
            .O(N__38397),
            .I(N__38394));
    Span4Mux_v I__6139 (
            .O(N__38394),
            .I(N__38390));
    InMux I__6138 (
            .O(N__38393),
            .I(N__38387));
    Sp12to4 I__6137 (
            .O(N__38390),
            .I(N__38384));
    LocalMux I__6136 (
            .O(N__38387),
            .I(\c0.tx.r_Clock_Count_0 ));
    Odrv12 I__6135 (
            .O(N__38384),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__6134 (
            .O(N__38379),
            .I(N__38376));
    LocalMux I__6133 (
            .O(N__38376),
            .I(N__38373));
    Span4Mux_h I__6132 (
            .O(N__38373),
            .I(N__38370));
    Odrv4 I__6131 (
            .O(N__38370),
            .I(n2265));
    CascadeMux I__6130 (
            .O(N__38367),
            .I(N__38362));
    CascadeMux I__6129 (
            .O(N__38366),
            .I(N__38359));
    CascadeMux I__6128 (
            .O(N__38365),
            .I(N__38356));
    InMux I__6127 (
            .O(N__38362),
            .I(N__38353));
    InMux I__6126 (
            .O(N__38359),
            .I(N__38350));
    InMux I__6125 (
            .O(N__38356),
            .I(N__38347));
    LocalMux I__6124 (
            .O(N__38353),
            .I(N__38344));
    LocalMux I__6123 (
            .O(N__38350),
            .I(N__38338));
    LocalMux I__6122 (
            .O(N__38347),
            .I(N__38338));
    Span4Mux_h I__6121 (
            .O(N__38344),
            .I(N__38335));
    InMux I__6120 (
            .O(N__38343),
            .I(N__38332));
    Span4Mux_v I__6119 (
            .O(N__38338),
            .I(N__38329));
    Span4Mux_v I__6118 (
            .O(N__38335),
            .I(N__38326));
    LocalMux I__6117 (
            .O(N__38332),
            .I(encoder1_position_26));
    Odrv4 I__6116 (
            .O(N__38329),
            .I(encoder1_position_26));
    Odrv4 I__6115 (
            .O(N__38326),
            .I(encoder1_position_26));
    InMux I__6114 (
            .O(N__38319),
            .I(N__38315));
    InMux I__6113 (
            .O(N__38318),
            .I(N__38312));
    LocalMux I__6112 (
            .O(N__38315),
            .I(data_out_frame_10_1));
    LocalMux I__6111 (
            .O(N__38312),
            .I(data_out_frame_10_1));
    CascadeMux I__6110 (
            .O(N__38307),
            .I(N__38303));
    InMux I__6109 (
            .O(N__38306),
            .I(N__38300));
    InMux I__6108 (
            .O(N__38303),
            .I(N__38297));
    LocalMux I__6107 (
            .O(N__38300),
            .I(data_out_frame_11_1));
    LocalMux I__6106 (
            .O(N__38297),
            .I(data_out_frame_11_1));
    CascadeMux I__6105 (
            .O(N__38292),
            .I(\c0.n25116_cascade_ ));
    InMux I__6104 (
            .O(N__38289),
            .I(N__38285));
    InMux I__6103 (
            .O(N__38288),
            .I(N__38282));
    LocalMux I__6102 (
            .O(N__38285),
            .I(N__38279));
    LocalMux I__6101 (
            .O(N__38282),
            .I(data_out_frame_9_1));
    Odrv4 I__6100 (
            .O(N__38279),
            .I(data_out_frame_9_1));
    InMux I__6099 (
            .O(N__38274),
            .I(N__38271));
    LocalMux I__6098 (
            .O(N__38271),
            .I(N__38268));
    Odrv12 I__6097 (
            .O(N__38268),
            .I(\c0.n25119 ));
    CascadeMux I__6096 (
            .O(N__38265),
            .I(N__38259));
    CascadeMux I__6095 (
            .O(N__38264),
            .I(N__38255));
    CascadeMux I__6094 (
            .O(N__38263),
            .I(N__38251));
    InMux I__6093 (
            .O(N__38262),
            .I(N__38248));
    InMux I__6092 (
            .O(N__38259),
            .I(N__38245));
    InMux I__6091 (
            .O(N__38258),
            .I(N__38242));
    InMux I__6090 (
            .O(N__38255),
            .I(N__38239));
    InMux I__6089 (
            .O(N__38254),
            .I(N__38234));
    InMux I__6088 (
            .O(N__38251),
            .I(N__38234));
    LocalMux I__6087 (
            .O(N__38248),
            .I(N__38229));
    LocalMux I__6086 (
            .O(N__38245),
            .I(N__38229));
    LocalMux I__6085 (
            .O(N__38242),
            .I(N__38223));
    LocalMux I__6084 (
            .O(N__38239),
            .I(N__38220));
    LocalMux I__6083 (
            .O(N__38234),
            .I(N__38217));
    Span4Mux_v I__6082 (
            .O(N__38229),
            .I(N__38214));
    InMux I__6081 (
            .O(N__38228),
            .I(N__38209));
    InMux I__6080 (
            .O(N__38227),
            .I(N__38209));
    InMux I__6079 (
            .O(N__38226),
            .I(N__38206));
    Span4Mux_v I__6078 (
            .O(N__38223),
            .I(N__38203));
    Odrv4 I__6077 (
            .O(N__38220),
            .I(\c0.n22291 ));
    Odrv4 I__6076 (
            .O(N__38217),
            .I(\c0.n22291 ));
    Odrv4 I__6075 (
            .O(N__38214),
            .I(\c0.n22291 ));
    LocalMux I__6074 (
            .O(N__38209),
            .I(\c0.n22291 ));
    LocalMux I__6073 (
            .O(N__38206),
            .I(\c0.n22291 ));
    Odrv4 I__6072 (
            .O(N__38203),
            .I(\c0.n22291 ));
    CascadeMux I__6071 (
            .O(N__38190),
            .I(N__38186));
    CascadeMux I__6070 (
            .O(N__38189),
            .I(N__38181));
    InMux I__6069 (
            .O(N__38186),
            .I(N__38169));
    InMux I__6068 (
            .O(N__38185),
            .I(N__38169));
    InMux I__6067 (
            .O(N__38184),
            .I(N__38166));
    InMux I__6066 (
            .O(N__38181),
            .I(N__38155));
    InMux I__6065 (
            .O(N__38180),
            .I(N__38155));
    InMux I__6064 (
            .O(N__38179),
            .I(N__38155));
    InMux I__6063 (
            .O(N__38178),
            .I(N__38155));
    InMux I__6062 (
            .O(N__38177),
            .I(N__38150));
    InMux I__6061 (
            .O(N__38176),
            .I(N__38150));
    InMux I__6060 (
            .O(N__38175),
            .I(N__38147));
    InMux I__6059 (
            .O(N__38174),
            .I(N__38144));
    LocalMux I__6058 (
            .O(N__38169),
            .I(N__38139));
    LocalMux I__6057 (
            .O(N__38166),
            .I(N__38139));
    InMux I__6056 (
            .O(N__38165),
            .I(N__38134));
    InMux I__6055 (
            .O(N__38164),
            .I(N__38134));
    LocalMux I__6054 (
            .O(N__38155),
            .I(N__38129));
    LocalMux I__6053 (
            .O(N__38150),
            .I(N__38129));
    LocalMux I__6052 (
            .O(N__38147),
            .I(N__38126));
    LocalMux I__6051 (
            .O(N__38144),
            .I(N__38123));
    Span4Mux_v I__6050 (
            .O(N__38139),
            .I(N__38115));
    LocalMux I__6049 (
            .O(N__38134),
            .I(N__38115));
    Span4Mux_v I__6048 (
            .O(N__38129),
            .I(N__38115));
    Span4Mux_v I__6047 (
            .O(N__38126),
            .I(N__38112));
    Span12Mux_s11_h I__6046 (
            .O(N__38123),
            .I(N__38109));
    InMux I__6045 (
            .O(N__38122),
            .I(N__38106));
    Span4Mux_v I__6044 (
            .O(N__38115),
            .I(N__38101));
    Span4Mux_v I__6043 (
            .O(N__38112),
            .I(N__38101));
    Odrv12 I__6042 (
            .O(N__38109),
            .I(\c0.n20333 ));
    LocalMux I__6041 (
            .O(N__38106),
            .I(\c0.n20333 ));
    Odrv4 I__6040 (
            .O(N__38101),
            .I(\c0.n20333 ));
    InMux I__6039 (
            .O(N__38094),
            .I(N__38084));
    InMux I__6038 (
            .O(N__38093),
            .I(N__38084));
    InMux I__6037 (
            .O(N__38092),
            .I(N__38077));
    InMux I__6036 (
            .O(N__38091),
            .I(N__38077));
    InMux I__6035 (
            .O(N__38090),
            .I(N__38072));
    InMux I__6034 (
            .O(N__38089),
            .I(N__38072));
    LocalMux I__6033 (
            .O(N__38084),
            .I(N__38069));
    InMux I__6032 (
            .O(N__38083),
            .I(N__38066));
    InMux I__6031 (
            .O(N__38082),
            .I(N__38063));
    LocalMux I__6030 (
            .O(N__38077),
            .I(N__38060));
    LocalMux I__6029 (
            .O(N__38072),
            .I(N__38052));
    Span4Mux_h I__6028 (
            .O(N__38069),
            .I(N__38052));
    LocalMux I__6027 (
            .O(N__38066),
            .I(N__38052));
    LocalMux I__6026 (
            .O(N__38063),
            .I(N__38049));
    Span4Mux_h I__6025 (
            .O(N__38060),
            .I(N__38046));
    InMux I__6024 (
            .O(N__38059),
            .I(N__38043));
    Span4Mux_v I__6023 (
            .O(N__38052),
            .I(N__38038));
    Span4Mux_v I__6022 (
            .O(N__38049),
            .I(N__38038));
    Odrv4 I__6021 (
            .O(N__38046),
            .I(\c0.data_out_frame_29__7__N_1148 ));
    LocalMux I__6020 (
            .O(N__38043),
            .I(\c0.data_out_frame_29__7__N_1148 ));
    Odrv4 I__6019 (
            .O(N__38038),
            .I(\c0.data_out_frame_29__7__N_1148 ));
    InMux I__6018 (
            .O(N__38031),
            .I(N__38026));
    InMux I__6017 (
            .O(N__38030),
            .I(N__38022));
    InMux I__6016 (
            .O(N__38029),
            .I(N__38018));
    LocalMux I__6015 (
            .O(N__38026),
            .I(N__38015));
    InMux I__6014 (
            .O(N__38025),
            .I(N__38012));
    LocalMux I__6013 (
            .O(N__38022),
            .I(N__38007));
    InMux I__6012 (
            .O(N__38021),
            .I(N__38003));
    LocalMux I__6011 (
            .O(N__38018),
            .I(N__38000));
    Span4Mux_v I__6010 (
            .O(N__38015),
            .I(N__37995));
    LocalMux I__6009 (
            .O(N__38012),
            .I(N__37995));
    InMux I__6008 (
            .O(N__38011),
            .I(N__37990));
    InMux I__6007 (
            .O(N__38010),
            .I(N__37990));
    Span4Mux_h I__6006 (
            .O(N__38007),
            .I(N__37987));
    InMux I__6005 (
            .O(N__38006),
            .I(N__37984));
    LocalMux I__6004 (
            .O(N__38003),
            .I(N__37979));
    Span4Mux_h I__6003 (
            .O(N__38000),
            .I(N__37979));
    Span4Mux_h I__6002 (
            .O(N__37995),
            .I(N__37976));
    LocalMux I__6001 (
            .O(N__37990),
            .I(N__37973));
    Odrv4 I__6000 (
            .O(N__37987),
            .I(\c0.n21464 ));
    LocalMux I__5999 (
            .O(N__37984),
            .I(\c0.n21464 ));
    Odrv4 I__5998 (
            .O(N__37979),
            .I(\c0.n21464 ));
    Odrv4 I__5997 (
            .O(N__37976),
            .I(\c0.n21464 ));
    Odrv12 I__5996 (
            .O(N__37973),
            .I(\c0.n21464 ));
    InMux I__5995 (
            .O(N__37962),
            .I(N__37959));
    LocalMux I__5994 (
            .O(N__37959),
            .I(N__37956));
    Span4Mux_v I__5993 (
            .O(N__37956),
            .I(N__37953));
    Odrv4 I__5992 (
            .O(N__37953),
            .I(n2267));
    CascadeMux I__5991 (
            .O(N__37950),
            .I(N__37947));
    InMux I__5990 (
            .O(N__37947),
            .I(N__37943));
    CascadeMux I__5989 (
            .O(N__37946),
            .I(N__37940));
    LocalMux I__5988 (
            .O(N__37943),
            .I(N__37935));
    InMux I__5987 (
            .O(N__37940),
            .I(N__37932));
    InMux I__5986 (
            .O(N__37939),
            .I(N__37927));
    InMux I__5985 (
            .O(N__37938),
            .I(N__37927));
    Span4Mux_h I__5984 (
            .O(N__37935),
            .I(N__37923));
    LocalMux I__5983 (
            .O(N__37932),
            .I(N__37920));
    LocalMux I__5982 (
            .O(N__37927),
            .I(N__37917));
    InMux I__5981 (
            .O(N__37926),
            .I(N__37914));
    Span4Mux_h I__5980 (
            .O(N__37923),
            .I(N__37911));
    Span4Mux_h I__5979 (
            .O(N__37920),
            .I(N__37906));
    Span4Mux_h I__5978 (
            .O(N__37917),
            .I(N__37906));
    LocalMux I__5977 (
            .O(N__37914),
            .I(encoder1_position_24));
    Odrv4 I__5976 (
            .O(N__37911),
            .I(encoder1_position_24));
    Odrv4 I__5975 (
            .O(N__37906),
            .I(encoder1_position_24));
    InMux I__5974 (
            .O(N__37899),
            .I(N__37896));
    LocalMux I__5973 (
            .O(N__37896),
            .I(N__37893));
    Span4Mux_h I__5972 (
            .O(N__37893),
            .I(N__37890));
    Span4Mux_v I__5971 (
            .O(N__37890),
            .I(N__37887));
    Odrv4 I__5970 (
            .O(N__37887),
            .I(\c0.n10_adj_4367 ));
    InMux I__5969 (
            .O(N__37884),
            .I(N__37881));
    LocalMux I__5968 (
            .O(N__37881),
            .I(\c0.n10_adj_4239 ));
    InMux I__5967 (
            .O(N__37878),
            .I(N__37875));
    LocalMux I__5966 (
            .O(N__37875),
            .I(\c0.n13049 ));
    InMux I__5965 (
            .O(N__37872),
            .I(N__37869));
    LocalMux I__5964 (
            .O(N__37869),
            .I(N__37866));
    Span4Mux_v I__5963 (
            .O(N__37866),
            .I(N__37862));
    InMux I__5962 (
            .O(N__37865),
            .I(N__37857));
    Span4Mux_h I__5961 (
            .O(N__37862),
            .I(N__37854));
    InMux I__5960 (
            .O(N__37861),
            .I(N__37851));
    InMux I__5959 (
            .O(N__37860),
            .I(N__37848));
    LocalMux I__5958 (
            .O(N__37857),
            .I(data_in_2_4));
    Odrv4 I__5957 (
            .O(N__37854),
            .I(data_in_2_4));
    LocalMux I__5956 (
            .O(N__37851),
            .I(data_in_2_4));
    LocalMux I__5955 (
            .O(N__37848),
            .I(data_in_2_4));
    CascadeMux I__5954 (
            .O(N__37839),
            .I(\c0.n13049_cascade_ ));
    CascadeMux I__5953 (
            .O(N__37836),
            .I(\c0.n18_adj_4236_cascade_ ));
    InMux I__5952 (
            .O(N__37833),
            .I(N__37830));
    LocalMux I__5951 (
            .O(N__37830),
            .I(\c0.n20_adj_4237 ));
    CascadeMux I__5950 (
            .O(N__37827),
            .I(N__37823));
    InMux I__5949 (
            .O(N__37826),
            .I(N__37819));
    InMux I__5948 (
            .O(N__37823),
            .I(N__37816));
    InMux I__5947 (
            .O(N__37822),
            .I(N__37813));
    LocalMux I__5946 (
            .O(N__37819),
            .I(N__37809));
    LocalMux I__5945 (
            .O(N__37816),
            .I(N__37804));
    LocalMux I__5944 (
            .O(N__37813),
            .I(N__37804));
    InMux I__5943 (
            .O(N__37812),
            .I(N__37801));
    Span4Mux_v I__5942 (
            .O(N__37809),
            .I(N__37796));
    Span4Mux_v I__5941 (
            .O(N__37804),
            .I(N__37796));
    LocalMux I__5940 (
            .O(N__37801),
            .I(data_in_1_4));
    Odrv4 I__5939 (
            .O(N__37796),
            .I(data_in_1_4));
    InMux I__5938 (
            .O(N__37791),
            .I(N__37788));
    LocalMux I__5937 (
            .O(N__37788),
            .I(\c0.n14_adj_4241 ));
    InMux I__5936 (
            .O(N__37785),
            .I(N__37782));
    LocalMux I__5935 (
            .O(N__37782),
            .I(\c0.n22489 ));
    InMux I__5934 (
            .O(N__37779),
            .I(N__37775));
    InMux I__5933 (
            .O(N__37778),
            .I(N__37772));
    LocalMux I__5932 (
            .O(N__37775),
            .I(N__37769));
    LocalMux I__5931 (
            .O(N__37772),
            .I(N__37766));
    Odrv4 I__5930 (
            .O(N__37769),
            .I(\c0.n21393 ));
    Odrv4 I__5929 (
            .O(N__37766),
            .I(\c0.n21393 ));
    CascadeMux I__5928 (
            .O(N__37761),
            .I(N__37758));
    InMux I__5927 (
            .O(N__37758),
            .I(N__37755));
    LocalMux I__5926 (
            .O(N__37755),
            .I(\c0.n22797 ));
    InMux I__5925 (
            .O(N__37752),
            .I(N__37749));
    LocalMux I__5924 (
            .O(N__37749),
            .I(N__37746));
    Odrv12 I__5923 (
            .O(N__37746),
            .I(\c0.n26_adj_4697 ));
    InMux I__5922 (
            .O(N__37743),
            .I(N__37739));
    InMux I__5921 (
            .O(N__37742),
            .I(N__37736));
    LocalMux I__5920 (
            .O(N__37739),
            .I(N__37733));
    LocalMux I__5919 (
            .O(N__37736),
            .I(N__37730));
    Odrv12 I__5918 (
            .O(N__37733),
            .I(\c0.n22475 ));
    Odrv4 I__5917 (
            .O(N__37730),
            .I(\c0.n22475 ));
    InMux I__5916 (
            .O(N__37725),
            .I(N__37722));
    LocalMux I__5915 (
            .O(N__37722),
            .I(N__37718));
    InMux I__5914 (
            .O(N__37721),
            .I(N__37715));
    Odrv12 I__5913 (
            .O(N__37718),
            .I(\c0.data_out_frame_29__7__N_1143 ));
    LocalMux I__5912 (
            .O(N__37715),
            .I(\c0.data_out_frame_29__7__N_1143 ));
    InMux I__5911 (
            .O(N__37710),
            .I(N__37707));
    LocalMux I__5910 (
            .O(N__37707),
            .I(N__37704));
    Span4Mux_h I__5909 (
            .O(N__37704),
            .I(N__37701));
    Odrv4 I__5908 (
            .O(N__37701),
            .I(\c0.n10_adj_4214 ));
    InMux I__5907 (
            .O(N__37698),
            .I(N__37695));
    LocalMux I__5906 (
            .O(N__37695),
            .I(N__37692));
    Span4Mux_h I__5905 (
            .O(N__37692),
            .I(N__37689));
    Span4Mux_h I__5904 (
            .O(N__37689),
            .I(N__37686));
    Odrv4 I__5903 (
            .O(N__37686),
            .I(\c0.data_out_frame_28_1 ));
    CascadeMux I__5902 (
            .O(N__37683),
            .I(N__37680));
    InMux I__5901 (
            .O(N__37680),
            .I(N__37677));
    LocalMux I__5900 (
            .O(N__37677),
            .I(N__37674));
    Odrv12 I__5899 (
            .O(N__37674),
            .I(\c0.n24033 ));
    InMux I__5898 (
            .O(N__37671),
            .I(N__37668));
    LocalMux I__5897 (
            .O(N__37668),
            .I(\c0.n27_adj_4696 ));
    InMux I__5896 (
            .O(N__37665),
            .I(N__37661));
    InMux I__5895 (
            .O(N__37664),
            .I(N__37658));
    LocalMux I__5894 (
            .O(N__37661),
            .I(data_in_0_0));
    LocalMux I__5893 (
            .O(N__37658),
            .I(data_in_0_0));
    CascadeMux I__5892 (
            .O(N__37653),
            .I(N__37649));
    InMux I__5891 (
            .O(N__37652),
            .I(N__37644));
    InMux I__5890 (
            .O(N__37649),
            .I(N__37644));
    LocalMux I__5889 (
            .O(N__37644),
            .I(data_in_0_4));
    CascadeMux I__5888 (
            .O(N__37641),
            .I(\c0.n15_adj_4242_cascade_ ));
    InMux I__5887 (
            .O(N__37638),
            .I(N__37634));
    InMux I__5886 (
            .O(N__37637),
            .I(N__37631));
    LocalMux I__5885 (
            .O(N__37634),
            .I(\c0.n20766 ));
    LocalMux I__5884 (
            .O(N__37631),
            .I(\c0.n20766 ));
    InMux I__5883 (
            .O(N__37626),
            .I(N__37623));
    LocalMux I__5882 (
            .O(N__37623),
            .I(N__37620));
    Odrv4 I__5881 (
            .O(N__37620),
            .I(n2335));
    CascadeMux I__5880 (
            .O(N__37617),
            .I(N__37614));
    InMux I__5879 (
            .O(N__37614),
            .I(N__37611));
    LocalMux I__5878 (
            .O(N__37611),
            .I(\c0.n10427 ));
    CascadeMux I__5877 (
            .O(N__37608),
            .I(\c0.n21360_cascade_ ));
    InMux I__5876 (
            .O(N__37605),
            .I(N__37602));
    LocalMux I__5875 (
            .O(N__37602),
            .I(N__37598));
    InMux I__5874 (
            .O(N__37601),
            .I(N__37594));
    Span4Mux_h I__5873 (
            .O(N__37598),
            .I(N__37591));
    InMux I__5872 (
            .O(N__37597),
            .I(N__37588));
    LocalMux I__5871 (
            .O(N__37594),
            .I(\c0.n10504 ));
    Odrv4 I__5870 (
            .O(N__37591),
            .I(\c0.n10504 ));
    LocalMux I__5869 (
            .O(N__37588),
            .I(\c0.n10504 ));
    InMux I__5868 (
            .O(N__37581),
            .I(N__37578));
    LocalMux I__5867 (
            .O(N__37578),
            .I(N__37574));
    InMux I__5866 (
            .O(N__37577),
            .I(N__37571));
    Span4Mux_h I__5865 (
            .O(N__37574),
            .I(N__37568));
    LocalMux I__5864 (
            .O(N__37571),
            .I(N__37565));
    Odrv4 I__5863 (
            .O(N__37568),
            .I(\c0.n22366 ));
    Odrv12 I__5862 (
            .O(N__37565),
            .I(\c0.n22366 ));
    CascadeMux I__5861 (
            .O(N__37560),
            .I(\c0.n10504_cascade_ ));
    InMux I__5860 (
            .O(N__37557),
            .I(N__37551));
    InMux I__5859 (
            .O(N__37556),
            .I(N__37551));
    LocalMux I__5858 (
            .O(N__37551),
            .I(N__37548));
    Odrv4 I__5857 (
            .O(N__37548),
            .I(\c0.n22327 ));
    InMux I__5856 (
            .O(N__37545),
            .I(N__37542));
    LocalMux I__5855 (
            .O(N__37542),
            .I(N__37539));
    Span4Mux_v I__5854 (
            .O(N__37539),
            .I(N__37536));
    Span4Mux_h I__5853 (
            .O(N__37536),
            .I(N__37532));
    InMux I__5852 (
            .O(N__37535),
            .I(N__37529));
    Sp12to4 I__5851 (
            .O(N__37532),
            .I(N__37524));
    LocalMux I__5850 (
            .O(N__37529),
            .I(N__37524));
    Odrv12 I__5849 (
            .O(N__37524),
            .I(n21484));
    InMux I__5848 (
            .O(N__37521),
            .I(N__37518));
    LocalMux I__5847 (
            .O(N__37518),
            .I(N__37515));
    Span4Mux_h I__5846 (
            .O(N__37515),
            .I(N__37512));
    Odrv4 I__5845 (
            .O(N__37512),
            .I(\c0.n28_adj_4698 ));
    CascadeMux I__5844 (
            .O(N__37509),
            .I(\c0.n25_adj_4695_cascade_ ));
    CascadeMux I__5843 (
            .O(N__37506),
            .I(N__37503));
    InMux I__5842 (
            .O(N__37503),
            .I(N__37500));
    LocalMux I__5841 (
            .O(N__37500),
            .I(N__37497));
    Span12Mux_v I__5840 (
            .O(N__37497),
            .I(N__37494));
    Odrv12 I__5839 (
            .O(N__37494),
            .I(\c0.data_out_frame_29_1 ));
    CascadeMux I__5838 (
            .O(N__37491),
            .I(N__37480));
    CascadeMux I__5837 (
            .O(N__37490),
            .I(N__37475));
    CascadeMux I__5836 (
            .O(N__37489),
            .I(N__37471));
    CascadeMux I__5835 (
            .O(N__37488),
            .I(N__37467));
    CascadeMux I__5834 (
            .O(N__37487),
            .I(N__37463));
    CascadeMux I__5833 (
            .O(N__37486),
            .I(N__37459));
    CascadeMux I__5832 (
            .O(N__37485),
            .I(N__37455));
    CascadeMux I__5831 (
            .O(N__37484),
            .I(N__37451));
    InMux I__5830 (
            .O(N__37483),
            .I(N__37441));
    InMux I__5829 (
            .O(N__37480),
            .I(N__37436));
    InMux I__5828 (
            .O(N__37479),
            .I(N__37436));
    InMux I__5827 (
            .O(N__37478),
            .I(N__37423));
    InMux I__5826 (
            .O(N__37475),
            .I(N__37423));
    InMux I__5825 (
            .O(N__37474),
            .I(N__37423));
    InMux I__5824 (
            .O(N__37471),
            .I(N__37423));
    InMux I__5823 (
            .O(N__37470),
            .I(N__37423));
    InMux I__5822 (
            .O(N__37467),
            .I(N__37423));
    InMux I__5821 (
            .O(N__37466),
            .I(N__37406));
    InMux I__5820 (
            .O(N__37463),
            .I(N__37406));
    InMux I__5819 (
            .O(N__37462),
            .I(N__37406));
    InMux I__5818 (
            .O(N__37459),
            .I(N__37406));
    InMux I__5817 (
            .O(N__37458),
            .I(N__37406));
    InMux I__5816 (
            .O(N__37455),
            .I(N__37406));
    InMux I__5815 (
            .O(N__37454),
            .I(N__37406));
    InMux I__5814 (
            .O(N__37451),
            .I(N__37406));
    CascadeMux I__5813 (
            .O(N__37450),
            .I(N__37403));
    CascadeMux I__5812 (
            .O(N__37449),
            .I(N__37400));
    CascadeMux I__5811 (
            .O(N__37448),
            .I(N__37397));
    CascadeMux I__5810 (
            .O(N__37447),
            .I(N__37394));
    CascadeMux I__5809 (
            .O(N__37446),
            .I(N__37391));
    CascadeMux I__5808 (
            .O(N__37445),
            .I(N__37388));
    CascadeMux I__5807 (
            .O(N__37444),
            .I(N__37385));
    LocalMux I__5806 (
            .O(N__37441),
            .I(N__37371));
    LocalMux I__5805 (
            .O(N__37436),
            .I(N__37371));
    LocalMux I__5804 (
            .O(N__37423),
            .I(N__37371));
    LocalMux I__5803 (
            .O(N__37406),
            .I(N__37371));
    InMux I__5802 (
            .O(N__37403),
            .I(N__37362));
    InMux I__5801 (
            .O(N__37400),
            .I(N__37362));
    InMux I__5800 (
            .O(N__37397),
            .I(N__37362));
    InMux I__5799 (
            .O(N__37394),
            .I(N__37362));
    InMux I__5798 (
            .O(N__37391),
            .I(N__37353));
    InMux I__5797 (
            .O(N__37388),
            .I(N__37353));
    InMux I__5796 (
            .O(N__37385),
            .I(N__37353));
    InMux I__5795 (
            .O(N__37384),
            .I(N__37353));
    CascadeMux I__5794 (
            .O(N__37383),
            .I(N__37350));
    CascadeMux I__5793 (
            .O(N__37382),
            .I(N__37346));
    CascadeMux I__5792 (
            .O(N__37381),
            .I(N__37342));
    CascadeMux I__5791 (
            .O(N__37380),
            .I(N__37338));
    Span4Mux_v I__5790 (
            .O(N__37371),
            .I(N__37334));
    LocalMux I__5789 (
            .O(N__37362),
            .I(N__37331));
    LocalMux I__5788 (
            .O(N__37353),
            .I(N__37328));
    InMux I__5787 (
            .O(N__37350),
            .I(N__37311));
    InMux I__5786 (
            .O(N__37349),
            .I(N__37311));
    InMux I__5785 (
            .O(N__37346),
            .I(N__37311));
    InMux I__5784 (
            .O(N__37345),
            .I(N__37311));
    InMux I__5783 (
            .O(N__37342),
            .I(N__37311));
    InMux I__5782 (
            .O(N__37341),
            .I(N__37311));
    InMux I__5781 (
            .O(N__37338),
            .I(N__37311));
    InMux I__5780 (
            .O(N__37337),
            .I(N__37311));
    Span4Mux_h I__5779 (
            .O(N__37334),
            .I(N__37304));
    Span4Mux_h I__5778 (
            .O(N__37331),
            .I(N__37304));
    Span4Mux_h I__5777 (
            .O(N__37328),
            .I(N__37304));
    LocalMux I__5776 (
            .O(N__37311),
            .I(N__37301));
    Span4Mux_h I__5775 (
            .O(N__37304),
            .I(N__37298));
    Odrv12 I__5774 (
            .O(N__37301),
            .I(\quad_counter0.n2313 ));
    Odrv4 I__5773 (
            .O(N__37298),
            .I(\quad_counter0.n2313 ));
    InMux I__5772 (
            .O(N__37293),
            .I(bfn_14_13_0_));
    CascadeMux I__5771 (
            .O(N__37290),
            .I(n2326_cascade_));
    InMux I__5770 (
            .O(N__37287),
            .I(N__37284));
    LocalMux I__5769 (
            .O(N__37284),
            .I(N__37280));
    InMux I__5768 (
            .O(N__37283),
            .I(N__37277));
    Span12Mux_s10_h I__5767 (
            .O(N__37280),
            .I(N__37272));
    LocalMux I__5766 (
            .O(N__37277),
            .I(N__37272));
    Span12Mux_h I__5765 (
            .O(N__37272),
            .I(N__37269));
    Odrv12 I__5764 (
            .O(N__37269),
            .I(\c0.n22218 ));
    CascadeMux I__5763 (
            .O(N__37266),
            .I(N__37262));
    InMux I__5762 (
            .O(N__37265),
            .I(N__37259));
    InMux I__5761 (
            .O(N__37262),
            .I(N__37255));
    LocalMux I__5760 (
            .O(N__37259),
            .I(N__37252));
    InMux I__5759 (
            .O(N__37258),
            .I(N__37249));
    LocalMux I__5758 (
            .O(N__37255),
            .I(N__37246));
    Span4Mux_v I__5757 (
            .O(N__37252),
            .I(N__37243));
    LocalMux I__5756 (
            .O(N__37249),
            .I(N__37240));
    Span4Mux_v I__5755 (
            .O(N__37246),
            .I(N__37235));
    Span4Mux_h I__5754 (
            .O(N__37243),
            .I(N__37235));
    Span4Mux_v I__5753 (
            .O(N__37240),
            .I(N__37232));
    Odrv4 I__5752 (
            .O(N__37235),
            .I(\c0.n21323 ));
    Odrv4 I__5751 (
            .O(N__37232),
            .I(\c0.n21323 ));
    InMux I__5750 (
            .O(N__37227),
            .I(N__37224));
    LocalMux I__5749 (
            .O(N__37224),
            .I(N__37221));
    Odrv4 I__5748 (
            .O(N__37221),
            .I(\c0.n22671 ));
    InMux I__5747 (
            .O(N__37218),
            .I(N__37215));
    LocalMux I__5746 (
            .O(N__37215),
            .I(N__37212));
    Odrv12 I__5745 (
            .O(N__37212),
            .I(\c0.n20_adj_4694 ));
    InMux I__5744 (
            .O(N__37209),
            .I(N__37205));
    InMux I__5743 (
            .O(N__37208),
            .I(N__37202));
    LocalMux I__5742 (
            .O(N__37205),
            .I(N__37198));
    LocalMux I__5741 (
            .O(N__37202),
            .I(N__37195));
    InMux I__5740 (
            .O(N__37201),
            .I(N__37192));
    Span4Mux_h I__5739 (
            .O(N__37198),
            .I(N__37189));
    Span4Mux_h I__5738 (
            .O(N__37195),
            .I(N__37183));
    LocalMux I__5737 (
            .O(N__37192),
            .I(N__37183));
    Span4Mux_v I__5736 (
            .O(N__37189),
            .I(N__37180));
    InMux I__5735 (
            .O(N__37188),
            .I(N__37177));
    Odrv4 I__5734 (
            .O(N__37183),
            .I(\c0.n20348 ));
    Odrv4 I__5733 (
            .O(N__37180),
            .I(\c0.n20348 ));
    LocalMux I__5732 (
            .O(N__37177),
            .I(\c0.n20348 ));
    CascadeMux I__5731 (
            .O(N__37170),
            .I(N__37165));
    InMux I__5730 (
            .O(N__37169),
            .I(N__37161));
    InMux I__5729 (
            .O(N__37168),
            .I(N__37158));
    InMux I__5728 (
            .O(N__37165),
            .I(N__37153));
    InMux I__5727 (
            .O(N__37164),
            .I(N__37153));
    LocalMux I__5726 (
            .O(N__37161),
            .I(\c0.n21330 ));
    LocalMux I__5725 (
            .O(N__37158),
            .I(\c0.n21330 ));
    LocalMux I__5724 (
            .O(N__37153),
            .I(\c0.n21330 ));
    CascadeMux I__5723 (
            .O(N__37146),
            .I(\c0.n21355_cascade_ ));
    InMux I__5722 (
            .O(N__37143),
            .I(N__37140));
    LocalMux I__5721 (
            .O(N__37140),
            .I(N__37134));
    InMux I__5720 (
            .O(N__37139),
            .I(N__37131));
    CascadeMux I__5719 (
            .O(N__37138),
            .I(N__37128));
    InMux I__5718 (
            .O(N__37137),
            .I(N__37125));
    Span4Mux_v I__5717 (
            .O(N__37134),
            .I(N__37120));
    LocalMux I__5716 (
            .O(N__37131),
            .I(N__37120));
    InMux I__5715 (
            .O(N__37128),
            .I(N__37117));
    LocalMux I__5714 (
            .O(N__37125),
            .I(N__37112));
    Span4Mux_h I__5713 (
            .O(N__37120),
            .I(N__37107));
    LocalMux I__5712 (
            .O(N__37117),
            .I(N__37107));
    InMux I__5711 (
            .O(N__37116),
            .I(N__37104));
    InMux I__5710 (
            .O(N__37115),
            .I(N__37101));
    Odrv4 I__5709 (
            .O(N__37112),
            .I(\c0.n12464 ));
    Odrv4 I__5708 (
            .O(N__37107),
            .I(\c0.n12464 ));
    LocalMux I__5707 (
            .O(N__37104),
            .I(\c0.n12464 ));
    LocalMux I__5706 (
            .O(N__37101),
            .I(\c0.n12464 ));
    InMux I__5705 (
            .O(N__37092),
            .I(N__37088));
    InMux I__5704 (
            .O(N__37091),
            .I(N__37085));
    LocalMux I__5703 (
            .O(N__37088),
            .I(\c0.n20404 ));
    LocalMux I__5702 (
            .O(N__37085),
            .I(\c0.n20404 ));
    InMux I__5701 (
            .O(N__37080),
            .I(\quad_counter0.n19785 ));
    InMux I__5700 (
            .O(N__37077),
            .I(bfn_14_12_0_));
    InMux I__5699 (
            .O(N__37074),
            .I(N__37071));
    LocalMux I__5698 (
            .O(N__37071),
            .I(n2333));
    InMux I__5697 (
            .O(N__37068),
            .I(\quad_counter0.n19787 ));
    InMux I__5696 (
            .O(N__37065),
            .I(N__37062));
    LocalMux I__5695 (
            .O(N__37062),
            .I(n2332));
    InMux I__5694 (
            .O(N__37059),
            .I(\quad_counter0.n19788 ));
    CascadeMux I__5693 (
            .O(N__37056),
            .I(N__37053));
    InMux I__5692 (
            .O(N__37053),
            .I(N__37049));
    InMux I__5691 (
            .O(N__37052),
            .I(N__37046));
    LocalMux I__5690 (
            .O(N__37049),
            .I(N__37042));
    LocalMux I__5689 (
            .O(N__37046),
            .I(N__37039));
    CascadeMux I__5688 (
            .O(N__37045),
            .I(N__37036));
    Span12Mux_v I__5687 (
            .O(N__37042),
            .I(N__37030));
    Span4Mux_h I__5686 (
            .O(N__37039),
            .I(N__37027));
    InMux I__5685 (
            .O(N__37036),
            .I(N__37022));
    InMux I__5684 (
            .O(N__37035),
            .I(N__37022));
    InMux I__5683 (
            .O(N__37034),
            .I(N__37017));
    InMux I__5682 (
            .O(N__37033),
            .I(N__37017));
    Odrv12 I__5681 (
            .O(N__37030),
            .I(encoder0_position_26));
    Odrv4 I__5680 (
            .O(N__37027),
            .I(encoder0_position_26));
    LocalMux I__5679 (
            .O(N__37022),
            .I(encoder0_position_26));
    LocalMux I__5678 (
            .O(N__37017),
            .I(encoder0_position_26));
    InMux I__5677 (
            .O(N__37008),
            .I(N__37005));
    LocalMux I__5676 (
            .O(N__37005),
            .I(N__37002));
    Span4Mux_v I__5675 (
            .O(N__37002),
            .I(N__36999));
    Odrv4 I__5674 (
            .O(N__36999),
            .I(n2331));
    InMux I__5673 (
            .O(N__36996),
            .I(\quad_counter0.n19789 ));
    InMux I__5672 (
            .O(N__36993),
            .I(N__36990));
    LocalMux I__5671 (
            .O(N__36990),
            .I(n2330));
    InMux I__5670 (
            .O(N__36987),
            .I(\quad_counter0.n19790 ));
    InMux I__5669 (
            .O(N__36984),
            .I(N__36981));
    LocalMux I__5668 (
            .O(N__36981),
            .I(N__36978));
    Span4Mux_v I__5667 (
            .O(N__36978),
            .I(N__36971));
    InMux I__5666 (
            .O(N__36977),
            .I(N__36968));
    InMux I__5665 (
            .O(N__36976),
            .I(N__36965));
    CascadeMux I__5664 (
            .O(N__36975),
            .I(N__36961));
    CascadeMux I__5663 (
            .O(N__36974),
            .I(N__36958));
    Span4Mux_v I__5662 (
            .O(N__36971),
            .I(N__36952));
    LocalMux I__5661 (
            .O(N__36968),
            .I(N__36952));
    LocalMux I__5660 (
            .O(N__36965),
            .I(N__36948));
    InMux I__5659 (
            .O(N__36964),
            .I(N__36945));
    InMux I__5658 (
            .O(N__36961),
            .I(N__36940));
    InMux I__5657 (
            .O(N__36958),
            .I(N__36940));
    InMux I__5656 (
            .O(N__36957),
            .I(N__36937));
    Span4Mux_v I__5655 (
            .O(N__36952),
            .I(N__36934));
    InMux I__5654 (
            .O(N__36951),
            .I(N__36931));
    Span4Mux_v I__5653 (
            .O(N__36948),
            .I(N__36928));
    LocalMux I__5652 (
            .O(N__36945),
            .I(N__36923));
    LocalMux I__5651 (
            .O(N__36940),
            .I(N__36923));
    LocalMux I__5650 (
            .O(N__36937),
            .I(encoder0_position_28));
    Odrv4 I__5649 (
            .O(N__36934),
            .I(encoder0_position_28));
    LocalMux I__5648 (
            .O(N__36931),
            .I(encoder0_position_28));
    Odrv4 I__5647 (
            .O(N__36928),
            .I(encoder0_position_28));
    Odrv4 I__5646 (
            .O(N__36923),
            .I(encoder0_position_28));
    InMux I__5645 (
            .O(N__36912),
            .I(N__36909));
    LocalMux I__5644 (
            .O(N__36909),
            .I(N__36906));
    Span4Mux_h I__5643 (
            .O(N__36906),
            .I(N__36903));
    Odrv4 I__5642 (
            .O(N__36903),
            .I(n2329));
    InMux I__5641 (
            .O(N__36900),
            .I(\quad_counter0.n19791 ));
    InMux I__5640 (
            .O(N__36897),
            .I(N__36894));
    LocalMux I__5639 (
            .O(N__36894),
            .I(N__36890));
    CascadeMux I__5638 (
            .O(N__36893),
            .I(N__36887));
    Span4Mux_v I__5637 (
            .O(N__36890),
            .I(N__36884));
    InMux I__5636 (
            .O(N__36887),
            .I(N__36881));
    Span4Mux_v I__5635 (
            .O(N__36884),
            .I(N__36878));
    LocalMux I__5634 (
            .O(N__36881),
            .I(N__36875));
    Span4Mux_v I__5633 (
            .O(N__36878),
            .I(N__36867));
    Span4Mux_h I__5632 (
            .O(N__36875),
            .I(N__36864));
    InMux I__5631 (
            .O(N__36874),
            .I(N__36857));
    InMux I__5630 (
            .O(N__36873),
            .I(N__36857));
    InMux I__5629 (
            .O(N__36872),
            .I(N__36857));
    InMux I__5628 (
            .O(N__36871),
            .I(N__36852));
    InMux I__5627 (
            .O(N__36870),
            .I(N__36852));
    Odrv4 I__5626 (
            .O(N__36867),
            .I(encoder0_position_29));
    Odrv4 I__5625 (
            .O(N__36864),
            .I(encoder0_position_29));
    LocalMux I__5624 (
            .O(N__36857),
            .I(encoder0_position_29));
    LocalMux I__5623 (
            .O(N__36852),
            .I(encoder0_position_29));
    InMux I__5622 (
            .O(N__36843),
            .I(N__36840));
    LocalMux I__5621 (
            .O(N__36840),
            .I(N__36837));
    Span4Mux_v I__5620 (
            .O(N__36837),
            .I(N__36834));
    Span4Mux_h I__5619 (
            .O(N__36834),
            .I(N__36831));
    Odrv4 I__5618 (
            .O(N__36831),
            .I(n2328));
    InMux I__5617 (
            .O(N__36828),
            .I(\quad_counter0.n19792 ));
    InMux I__5616 (
            .O(N__36825),
            .I(N__36822));
    LocalMux I__5615 (
            .O(N__36822),
            .I(N__36819));
    Odrv12 I__5614 (
            .O(N__36819),
            .I(n2327));
    InMux I__5613 (
            .O(N__36816),
            .I(\quad_counter0.n19793 ));
    InMux I__5612 (
            .O(N__36813),
            .I(\quad_counter0.n19776 ));
    InMux I__5611 (
            .O(N__36810),
            .I(\quad_counter0.n19777 ));
    InMux I__5610 (
            .O(N__36807),
            .I(bfn_14_11_0_));
    CascadeMux I__5609 (
            .O(N__36804),
            .I(N__36798));
    CascadeMux I__5608 (
            .O(N__36803),
            .I(N__36795));
    InMux I__5607 (
            .O(N__36802),
            .I(N__36792));
    InMux I__5606 (
            .O(N__36801),
            .I(N__36789));
    InMux I__5605 (
            .O(N__36798),
            .I(N__36785));
    InMux I__5604 (
            .O(N__36795),
            .I(N__36781));
    LocalMux I__5603 (
            .O(N__36792),
            .I(N__36776));
    LocalMux I__5602 (
            .O(N__36789),
            .I(N__36776));
    InMux I__5601 (
            .O(N__36788),
            .I(N__36773));
    LocalMux I__5600 (
            .O(N__36785),
            .I(N__36770));
    InMux I__5599 (
            .O(N__36784),
            .I(N__36767));
    LocalMux I__5598 (
            .O(N__36781),
            .I(N__36760));
    Span4Mux_v I__5597 (
            .O(N__36776),
            .I(N__36760));
    LocalMux I__5596 (
            .O(N__36773),
            .I(N__36760));
    Odrv4 I__5595 (
            .O(N__36770),
            .I(encoder0_position_16));
    LocalMux I__5594 (
            .O(N__36767),
            .I(encoder0_position_16));
    Odrv4 I__5593 (
            .O(N__36760),
            .I(encoder0_position_16));
    InMux I__5592 (
            .O(N__36753),
            .I(N__36750));
    LocalMux I__5591 (
            .O(N__36750),
            .I(N__36747));
    Odrv4 I__5590 (
            .O(N__36747),
            .I(n2341));
    InMux I__5589 (
            .O(N__36744),
            .I(\quad_counter0.n19779 ));
    InMux I__5588 (
            .O(N__36741),
            .I(\quad_counter0.n19780 ));
    InMux I__5587 (
            .O(N__36738),
            .I(\quad_counter0.n19781 ));
    InMux I__5586 (
            .O(N__36735),
            .I(\quad_counter0.n19782 ));
    InMux I__5585 (
            .O(N__36732),
            .I(\quad_counter0.n19783 ));
    InMux I__5584 (
            .O(N__36729),
            .I(\quad_counter0.n19784 ));
    InMux I__5583 (
            .O(N__36726),
            .I(\quad_counter0.n19768 ));
    InMux I__5582 (
            .O(N__36723),
            .I(N__36720));
    LocalMux I__5581 (
            .O(N__36720),
            .I(N__36717));
    Odrv4 I__5580 (
            .O(N__36717),
            .I(n2351));
    InMux I__5579 (
            .O(N__36714),
            .I(\quad_counter0.n19769 ));
    CascadeMux I__5578 (
            .O(N__36711),
            .I(N__36708));
    InMux I__5577 (
            .O(N__36708),
            .I(N__36703));
    InMux I__5576 (
            .O(N__36707),
            .I(N__36698));
    InMux I__5575 (
            .O(N__36706),
            .I(N__36698));
    LocalMux I__5574 (
            .O(N__36703),
            .I(N__36694));
    LocalMux I__5573 (
            .O(N__36698),
            .I(N__36690));
    InMux I__5572 (
            .O(N__36697),
            .I(N__36685));
    Span12Mux_v I__5571 (
            .O(N__36694),
            .I(N__36682));
    InMux I__5570 (
            .O(N__36693),
            .I(N__36679));
    Span4Mux_v I__5569 (
            .O(N__36690),
            .I(N__36676));
    InMux I__5568 (
            .O(N__36689),
            .I(N__36673));
    InMux I__5567 (
            .O(N__36688),
            .I(N__36670));
    LocalMux I__5566 (
            .O(N__36685),
            .I(N__36667));
    Span12Mux_v I__5565 (
            .O(N__36682),
            .I(N__36664));
    LocalMux I__5564 (
            .O(N__36679),
            .I(N__36659));
    Span4Mux_h I__5563 (
            .O(N__36676),
            .I(N__36659));
    LocalMux I__5562 (
            .O(N__36673),
            .I(N__36652));
    LocalMux I__5561 (
            .O(N__36670),
            .I(N__36652));
    Span4Mux_v I__5560 (
            .O(N__36667),
            .I(N__36652));
    Odrv12 I__5559 (
            .O(N__36664),
            .I(encoder0_position_7));
    Odrv4 I__5558 (
            .O(N__36659),
            .I(encoder0_position_7));
    Odrv4 I__5557 (
            .O(N__36652),
            .I(encoder0_position_7));
    InMux I__5556 (
            .O(N__36645),
            .I(N__36642));
    LocalMux I__5555 (
            .O(N__36642),
            .I(N__36639));
    Odrv4 I__5554 (
            .O(N__36639),
            .I(n2350));
    InMux I__5553 (
            .O(N__36636),
            .I(bfn_14_10_0_));
    InMux I__5552 (
            .O(N__36633),
            .I(\quad_counter0.n19771 ));
    InMux I__5551 (
            .O(N__36630),
            .I(\quad_counter0.n19772 ));
    CascadeMux I__5550 (
            .O(N__36627),
            .I(N__36624));
    InMux I__5549 (
            .O(N__36624),
            .I(N__36619));
    CascadeMux I__5548 (
            .O(N__36623),
            .I(N__36616));
    CascadeMux I__5547 (
            .O(N__36622),
            .I(N__36613));
    LocalMux I__5546 (
            .O(N__36619),
            .I(N__36610));
    InMux I__5545 (
            .O(N__36616),
            .I(N__36607));
    InMux I__5544 (
            .O(N__36613),
            .I(N__36604));
    Span4Mux_v I__5543 (
            .O(N__36610),
            .I(N__36599));
    LocalMux I__5542 (
            .O(N__36607),
            .I(N__36599));
    LocalMux I__5541 (
            .O(N__36604),
            .I(N__36594));
    Span4Mux_h I__5540 (
            .O(N__36599),
            .I(N__36591));
    InMux I__5539 (
            .O(N__36598),
            .I(N__36586));
    InMux I__5538 (
            .O(N__36597),
            .I(N__36586));
    Odrv12 I__5537 (
            .O(N__36594),
            .I(encoder0_position_10));
    Odrv4 I__5536 (
            .O(N__36591),
            .I(encoder0_position_10));
    LocalMux I__5535 (
            .O(N__36586),
            .I(encoder0_position_10));
    InMux I__5534 (
            .O(N__36579),
            .I(N__36576));
    LocalMux I__5533 (
            .O(N__36576),
            .I(N__36573));
    Span4Mux_h I__5532 (
            .O(N__36573),
            .I(N__36570));
    Odrv4 I__5531 (
            .O(N__36570),
            .I(n2347));
    InMux I__5530 (
            .O(N__36567),
            .I(\quad_counter0.n19773 ));
    CascadeMux I__5529 (
            .O(N__36564),
            .I(N__36561));
    InMux I__5528 (
            .O(N__36561),
            .I(N__36558));
    LocalMux I__5527 (
            .O(N__36558),
            .I(N__36555));
    Span4Mux_h I__5526 (
            .O(N__36555),
            .I(N__36551));
    InMux I__5525 (
            .O(N__36554),
            .I(N__36548));
    Span4Mux_v I__5524 (
            .O(N__36551),
            .I(N__36544));
    LocalMux I__5523 (
            .O(N__36548),
            .I(N__36541));
    InMux I__5522 (
            .O(N__36547),
            .I(N__36537));
    Span4Mux_h I__5521 (
            .O(N__36544),
            .I(N__36532));
    Span4Mux_h I__5520 (
            .O(N__36541),
            .I(N__36532));
    InMux I__5519 (
            .O(N__36540),
            .I(N__36529));
    LocalMux I__5518 (
            .O(N__36537),
            .I(encoder0_position_11));
    Odrv4 I__5517 (
            .O(N__36532),
            .I(encoder0_position_11));
    LocalMux I__5516 (
            .O(N__36529),
            .I(encoder0_position_11));
    InMux I__5515 (
            .O(N__36522),
            .I(N__36519));
    LocalMux I__5514 (
            .O(N__36519),
            .I(N__36516));
    Span4Mux_v I__5513 (
            .O(N__36516),
            .I(N__36513));
    Sp12to4 I__5512 (
            .O(N__36513),
            .I(N__36510));
    Odrv12 I__5511 (
            .O(N__36510),
            .I(n2346));
    InMux I__5510 (
            .O(N__36507),
            .I(\quad_counter0.n19774 ));
    CascadeMux I__5509 (
            .O(N__36504),
            .I(N__36501));
    InMux I__5508 (
            .O(N__36501),
            .I(N__36497));
    CascadeMux I__5507 (
            .O(N__36500),
            .I(N__36494));
    LocalMux I__5506 (
            .O(N__36497),
            .I(N__36491));
    InMux I__5505 (
            .O(N__36494),
            .I(N__36484));
    Span4Mux_h I__5504 (
            .O(N__36491),
            .I(N__36481));
    InMux I__5503 (
            .O(N__36490),
            .I(N__36476));
    InMux I__5502 (
            .O(N__36489),
            .I(N__36476));
    InMux I__5501 (
            .O(N__36488),
            .I(N__36473));
    InMux I__5500 (
            .O(N__36487),
            .I(N__36470));
    LocalMux I__5499 (
            .O(N__36484),
            .I(N__36467));
    Sp12to4 I__5498 (
            .O(N__36481),
            .I(N__36460));
    LocalMux I__5497 (
            .O(N__36476),
            .I(N__36460));
    LocalMux I__5496 (
            .O(N__36473),
            .I(N__36460));
    LocalMux I__5495 (
            .O(N__36470),
            .I(encoder0_position_12));
    Odrv12 I__5494 (
            .O(N__36467),
            .I(encoder0_position_12));
    Odrv12 I__5493 (
            .O(N__36460),
            .I(encoder0_position_12));
    InMux I__5492 (
            .O(N__36453),
            .I(N__36450));
    LocalMux I__5491 (
            .O(N__36450),
            .I(N__36447));
    Span4Mux_v I__5490 (
            .O(N__36447),
            .I(N__36444));
    Span4Mux_v I__5489 (
            .O(N__36444),
            .I(N__36441));
    Span4Mux_v I__5488 (
            .O(N__36441),
            .I(N__36438));
    Odrv4 I__5487 (
            .O(N__36438),
            .I(n2345));
    InMux I__5486 (
            .O(N__36435),
            .I(\quad_counter0.n19775 ));
    CascadeMux I__5485 (
            .O(N__36432),
            .I(N__36429));
    InMux I__5484 (
            .O(N__36429),
            .I(N__36426));
    LocalMux I__5483 (
            .O(N__36426),
            .I(N__36423));
    Span4Mux_h I__5482 (
            .O(N__36423),
            .I(N__36418));
    InMux I__5481 (
            .O(N__36422),
            .I(N__36415));
    InMux I__5480 (
            .O(N__36421),
            .I(N__36410));
    Span4Mux_v I__5479 (
            .O(N__36418),
            .I(N__36405));
    LocalMux I__5478 (
            .O(N__36415),
            .I(N__36405));
    InMux I__5477 (
            .O(N__36414),
            .I(N__36402));
    InMux I__5476 (
            .O(N__36413),
            .I(N__36399));
    LocalMux I__5475 (
            .O(N__36410),
            .I(N__36394));
    Span4Mux_v I__5474 (
            .O(N__36405),
            .I(N__36394));
    LocalMux I__5473 (
            .O(N__36402),
            .I(encoder0_position_0));
    LocalMux I__5472 (
            .O(N__36399),
            .I(encoder0_position_0));
    Odrv4 I__5471 (
            .O(N__36394),
            .I(encoder0_position_0));
    CascadeMux I__5470 (
            .O(N__36387),
            .I(N__36384));
    InMux I__5469 (
            .O(N__36384),
            .I(N__36381));
    LocalMux I__5468 (
            .O(N__36381),
            .I(N__36378));
    Span12Mux_s11_v I__5467 (
            .O(N__36378),
            .I(N__36375));
    Odrv12 I__5466 (
            .O(N__36375),
            .I(\quad_counter0.count_direction ));
    InMux I__5465 (
            .O(N__36372),
            .I(N__36369));
    LocalMux I__5464 (
            .O(N__36369),
            .I(n2357));
    InMux I__5463 (
            .O(N__36366),
            .I(\quad_counter0.n19763 ));
    CascadeMux I__5462 (
            .O(N__36363),
            .I(N__36360));
    InMux I__5461 (
            .O(N__36360),
            .I(N__36357));
    LocalMux I__5460 (
            .O(N__36357),
            .I(N__36353));
    InMux I__5459 (
            .O(N__36356),
            .I(N__36350));
    Sp12to4 I__5458 (
            .O(N__36353),
            .I(N__36346));
    LocalMux I__5457 (
            .O(N__36350),
            .I(N__36343));
    InMux I__5456 (
            .O(N__36349),
            .I(N__36338));
    Span12Mux_v I__5455 (
            .O(N__36346),
            .I(N__36335));
    Span4Mux_h I__5454 (
            .O(N__36343),
            .I(N__36332));
    InMux I__5453 (
            .O(N__36342),
            .I(N__36329));
    InMux I__5452 (
            .O(N__36341),
            .I(N__36326));
    LocalMux I__5451 (
            .O(N__36338),
            .I(encoder0_position_1));
    Odrv12 I__5450 (
            .O(N__36335),
            .I(encoder0_position_1));
    Odrv4 I__5449 (
            .O(N__36332),
            .I(encoder0_position_1));
    LocalMux I__5448 (
            .O(N__36329),
            .I(encoder0_position_1));
    LocalMux I__5447 (
            .O(N__36326),
            .I(encoder0_position_1));
    InMux I__5446 (
            .O(N__36315),
            .I(N__36312));
    LocalMux I__5445 (
            .O(N__36312),
            .I(N__36309));
    Span4Mux_h I__5444 (
            .O(N__36309),
            .I(N__36306));
    Odrv4 I__5443 (
            .O(N__36306),
            .I(n2356));
    InMux I__5442 (
            .O(N__36303),
            .I(\quad_counter0.n19764 ));
    InMux I__5441 (
            .O(N__36300),
            .I(N__36297));
    LocalMux I__5440 (
            .O(N__36297),
            .I(n2355));
    InMux I__5439 (
            .O(N__36294),
            .I(\quad_counter0.n19765 ));
    InMux I__5438 (
            .O(N__36291),
            .I(N__36288));
    LocalMux I__5437 (
            .O(N__36288),
            .I(n2354));
    InMux I__5436 (
            .O(N__36285),
            .I(\quad_counter0.n19766 ));
    InMux I__5435 (
            .O(N__36282),
            .I(N__36279));
    LocalMux I__5434 (
            .O(N__36279),
            .I(N__36276));
    Span4Mux_h I__5433 (
            .O(N__36276),
            .I(N__36273));
    Odrv4 I__5432 (
            .O(N__36273),
            .I(n2353));
    InMux I__5431 (
            .O(N__36270),
            .I(\quad_counter0.n19767 ));
    InMux I__5430 (
            .O(N__36267),
            .I(N__36260));
    InMux I__5429 (
            .O(N__36266),
            .I(N__36260));
    InMux I__5428 (
            .O(N__36265),
            .I(N__36256));
    LocalMux I__5427 (
            .O(N__36260),
            .I(N__36253));
    InMux I__5426 (
            .O(N__36259),
            .I(N__36250));
    LocalMux I__5425 (
            .O(N__36256),
            .I(N__36246));
    Span4Mux_v I__5424 (
            .O(N__36253),
            .I(N__36241));
    LocalMux I__5423 (
            .O(N__36250),
            .I(N__36241));
    InMux I__5422 (
            .O(N__36249),
            .I(N__36238));
    Span4Mux_h I__5421 (
            .O(N__36246),
            .I(N__36235));
    Span4Mux_h I__5420 (
            .O(N__36241),
            .I(N__36232));
    LocalMux I__5419 (
            .O(N__36238),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__5418 (
            .O(N__36235),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__5417 (
            .O(N__36232),
            .I(\c0.FRAME_MATCHER_state_25 ));
    SRMux I__5416 (
            .O(N__36225),
            .I(N__36222));
    LocalMux I__5415 (
            .O(N__36222),
            .I(N__36219));
    Span4Mux_h I__5414 (
            .O(N__36219),
            .I(N__36216));
    Odrv4 I__5413 (
            .O(N__36216),
            .I(\c0.n21653 ));
    InMux I__5412 (
            .O(N__36213),
            .I(N__36209));
    InMux I__5411 (
            .O(N__36212),
            .I(N__36206));
    LocalMux I__5410 (
            .O(N__36209),
            .I(N__36202));
    LocalMux I__5409 (
            .O(N__36206),
            .I(N__36199));
    InMux I__5408 (
            .O(N__36205),
            .I(N__36196));
    Span4Mux_h I__5407 (
            .O(N__36202),
            .I(N__36193));
    Span4Mux_h I__5406 (
            .O(N__36199),
            .I(N__36190));
    LocalMux I__5405 (
            .O(N__36196),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv4 I__5404 (
            .O(N__36193),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv4 I__5403 (
            .O(N__36190),
            .I(\c0.FRAME_MATCHER_state_29 ));
    SRMux I__5402 (
            .O(N__36183),
            .I(N__36180));
    LocalMux I__5401 (
            .O(N__36180),
            .I(N__36177));
    Span4Mux_v I__5400 (
            .O(N__36177),
            .I(N__36174));
    Odrv4 I__5399 (
            .O(N__36174),
            .I(\c0.n21649 ));
    CascadeMux I__5398 (
            .O(N__36171),
            .I(N__36167));
    InMux I__5397 (
            .O(N__36170),
            .I(N__36163));
    InMux I__5396 (
            .O(N__36167),
            .I(N__36160));
    CascadeMux I__5395 (
            .O(N__36166),
            .I(N__36156));
    LocalMux I__5394 (
            .O(N__36163),
            .I(N__36152));
    LocalMux I__5393 (
            .O(N__36160),
            .I(N__36149));
    InMux I__5392 (
            .O(N__36159),
            .I(N__36144));
    InMux I__5391 (
            .O(N__36156),
            .I(N__36144));
    InMux I__5390 (
            .O(N__36155),
            .I(N__36141));
    Span4Mux_h I__5389 (
            .O(N__36152),
            .I(N__36138));
    Span4Mux_h I__5388 (
            .O(N__36149),
            .I(N__36133));
    LocalMux I__5387 (
            .O(N__36144),
            .I(N__36133));
    LocalMux I__5386 (
            .O(N__36141),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__5385 (
            .O(N__36138),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__5384 (
            .O(N__36133),
            .I(\c0.FRAME_MATCHER_state_24 ));
    SRMux I__5383 (
            .O(N__36126),
            .I(N__36123));
    LocalMux I__5382 (
            .O(N__36123),
            .I(N__36120));
    Span4Mux_v I__5381 (
            .O(N__36120),
            .I(N__36117));
    Span4Mux_h I__5380 (
            .O(N__36117),
            .I(N__36114));
    Odrv4 I__5379 (
            .O(N__36114),
            .I(\c0.n21595 ));
    SRMux I__5378 (
            .O(N__36111),
            .I(N__36108));
    LocalMux I__5377 (
            .O(N__36108),
            .I(N__36105));
    Span4Mux_v I__5376 (
            .O(N__36105),
            .I(N__36102));
    Odrv4 I__5375 (
            .O(N__36102),
            .I(\c0.n21643 ));
    CascadeMux I__5374 (
            .O(N__36099),
            .I(N__36096));
    InMux I__5373 (
            .O(N__36096),
            .I(N__36093));
    LocalMux I__5372 (
            .O(N__36093),
            .I(N__36090));
    Span4Mux_v I__5371 (
            .O(N__36090),
            .I(N__36087));
    Sp12to4 I__5370 (
            .O(N__36087),
            .I(N__36084));
    Odrv12 I__5369 (
            .O(N__36084),
            .I(\c0.n6_adj_4583 ));
    InMux I__5368 (
            .O(N__36081),
            .I(N__36077));
    InMux I__5367 (
            .O(N__36080),
            .I(N__36073));
    LocalMux I__5366 (
            .O(N__36077),
            .I(N__36070));
    InMux I__5365 (
            .O(N__36076),
            .I(N__36067));
    LocalMux I__5364 (
            .O(N__36073),
            .I(N__36064));
    Span4Mux_h I__5363 (
            .O(N__36070),
            .I(N__36061));
    LocalMux I__5362 (
            .O(N__36067),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv4 I__5361 (
            .O(N__36064),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv4 I__5360 (
            .O(N__36061),
            .I(\c0.FRAME_MATCHER_state_6 ));
    InMux I__5359 (
            .O(N__36054),
            .I(N__36051));
    LocalMux I__5358 (
            .O(N__36051),
            .I(N__36048));
    Span4Mux_v I__5357 (
            .O(N__36048),
            .I(N__36045));
    Odrv4 I__5356 (
            .O(N__36045),
            .I(\c0.n14_adj_4520 ));
    CascadeMux I__5355 (
            .O(N__36042),
            .I(N__36038));
    InMux I__5354 (
            .O(N__36041),
            .I(N__36035));
    InMux I__5353 (
            .O(N__36038),
            .I(N__36032));
    LocalMux I__5352 (
            .O(N__36035),
            .I(N__36026));
    LocalMux I__5351 (
            .O(N__36032),
            .I(N__36026));
    InMux I__5350 (
            .O(N__36031),
            .I(N__36023));
    Span4Mux_h I__5349 (
            .O(N__36026),
            .I(N__36020));
    LocalMux I__5348 (
            .O(N__36023),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__5347 (
            .O(N__36020),
            .I(\c0.FRAME_MATCHER_state_4 ));
    InMux I__5346 (
            .O(N__36015),
            .I(N__36012));
    LocalMux I__5345 (
            .O(N__36012),
            .I(\c0.n9_adj_4522 ));
    InMux I__5344 (
            .O(N__36009),
            .I(N__36006));
    LocalMux I__5343 (
            .O(N__36006),
            .I(\c0.n20_adj_4265 ));
    InMux I__5342 (
            .O(N__36003),
            .I(N__36000));
    LocalMux I__5341 (
            .O(N__36000),
            .I(N__35996));
    InMux I__5340 (
            .O(N__35999),
            .I(N__35993));
    Span4Mux_h I__5339 (
            .O(N__35996),
            .I(N__35990));
    LocalMux I__5338 (
            .O(N__35993),
            .I(\c0.n16919 ));
    Odrv4 I__5337 (
            .O(N__35990),
            .I(\c0.n16919 ));
    CascadeMux I__5336 (
            .O(N__35985),
            .I(\c0.n20_adj_4265_cascade_ ));
    InMux I__5335 (
            .O(N__35982),
            .I(N__35979));
    LocalMux I__5334 (
            .O(N__35979),
            .I(N__35976));
    Span4Mux_h I__5333 (
            .O(N__35976),
            .I(N__35972));
    InMux I__5332 (
            .O(N__35975),
            .I(N__35969));
    Odrv4 I__5331 (
            .O(N__35972),
            .I(\c0.n22148 ));
    LocalMux I__5330 (
            .O(N__35969),
            .I(\c0.n22148 ));
    InMux I__5329 (
            .O(N__35964),
            .I(N__35960));
    InMux I__5328 (
            .O(N__35963),
            .I(N__35957));
    LocalMux I__5327 (
            .O(N__35960),
            .I(N__35954));
    LocalMux I__5326 (
            .O(N__35957),
            .I(N__35950));
    Span4Mux_v I__5325 (
            .O(N__35954),
            .I(N__35947));
    InMux I__5324 (
            .O(N__35953),
            .I(N__35944));
    Span4Mux_v I__5323 (
            .O(N__35950),
            .I(N__35940));
    Sp12to4 I__5322 (
            .O(N__35947),
            .I(N__35937));
    LocalMux I__5321 (
            .O(N__35944),
            .I(N__35934));
    InMux I__5320 (
            .O(N__35943),
            .I(N__35931));
    Odrv4 I__5319 (
            .O(N__35940),
            .I(\c0.n22145 ));
    Odrv12 I__5318 (
            .O(N__35937),
            .I(\c0.n22145 ));
    Odrv4 I__5317 (
            .O(N__35934),
            .I(\c0.n22145 ));
    LocalMux I__5316 (
            .O(N__35931),
            .I(\c0.n22145 ));
    InMux I__5315 (
            .O(N__35922),
            .I(N__35919));
    LocalMux I__5314 (
            .O(N__35919),
            .I(\c0.n6_adj_4264 ));
    InMux I__5313 (
            .O(N__35916),
            .I(N__35912));
    CascadeMux I__5312 (
            .O(N__35915),
            .I(N__35909));
    LocalMux I__5311 (
            .O(N__35912),
            .I(N__35905));
    InMux I__5310 (
            .O(N__35909),
            .I(N__35902));
    CascadeMux I__5309 (
            .O(N__35908),
            .I(N__35898));
    Span4Mux_v I__5308 (
            .O(N__35905),
            .I(N__35892));
    LocalMux I__5307 (
            .O(N__35902),
            .I(N__35892));
    InMux I__5306 (
            .O(N__35901),
            .I(N__35889));
    InMux I__5305 (
            .O(N__35898),
            .I(N__35886));
    InMux I__5304 (
            .O(N__35897),
            .I(N__35883));
    Span4Mux_h I__5303 (
            .O(N__35892),
            .I(N__35880));
    LocalMux I__5302 (
            .O(N__35889),
            .I(\c0.FRAME_MATCHER_state_22 ));
    LocalMux I__5301 (
            .O(N__35886),
            .I(\c0.FRAME_MATCHER_state_22 ));
    LocalMux I__5300 (
            .O(N__35883),
            .I(\c0.FRAME_MATCHER_state_22 ));
    Odrv4 I__5299 (
            .O(N__35880),
            .I(\c0.FRAME_MATCHER_state_22 ));
    CascadeMux I__5298 (
            .O(N__35871),
            .I(N__35868));
    InMux I__5297 (
            .O(N__35868),
            .I(N__35865));
    LocalMux I__5296 (
            .O(N__35865),
            .I(N__35862));
    Span4Mux_h I__5295 (
            .O(N__35862),
            .I(N__35859));
    Span4Mux_h I__5294 (
            .O(N__35859),
            .I(N__35856));
    Odrv4 I__5293 (
            .O(N__35856),
            .I(\c0.n14721 ));
    InMux I__5292 (
            .O(N__35853),
            .I(N__35850));
    LocalMux I__5291 (
            .O(N__35850),
            .I(N__35846));
    InMux I__5290 (
            .O(N__35849),
            .I(N__35843));
    Span4Mux_h I__5289 (
            .O(N__35846),
            .I(N__35840));
    LocalMux I__5288 (
            .O(N__35843),
            .I(N__35837));
    Sp12to4 I__5287 (
            .O(N__35840),
            .I(N__35834));
    Span4Mux_h I__5286 (
            .O(N__35837),
            .I(N__35831));
    Odrv12 I__5285 (
            .O(N__35834),
            .I(\c0.n14530 ));
    Odrv4 I__5284 (
            .O(N__35831),
            .I(\c0.n14530 ));
    InMux I__5283 (
            .O(N__35826),
            .I(N__35823));
    LocalMux I__5282 (
            .O(N__35823),
            .I(N__35820));
    Span12Mux_h I__5281 (
            .O(N__35820),
            .I(N__35817));
    Odrv12 I__5280 (
            .O(N__35817),
            .I(\c0.n7_adj_4741 ));
    CascadeMux I__5279 (
            .O(N__35814),
            .I(N__35810));
    InMux I__5278 (
            .O(N__35813),
            .I(N__35805));
    InMux I__5277 (
            .O(N__35810),
            .I(N__35805));
    LocalMux I__5276 (
            .O(N__35805),
            .I(N__35802));
    Odrv4 I__5275 (
            .O(N__35802),
            .I(\c0.n9683 ));
    InMux I__5274 (
            .O(N__35799),
            .I(N__35796));
    LocalMux I__5273 (
            .O(N__35796),
            .I(N__35793));
    Odrv4 I__5272 (
            .O(N__35793),
            .I(\c0.n9587 ));
    CascadeMux I__5271 (
            .O(N__35790),
            .I(\c0.n9683_cascade_ ));
    InMux I__5270 (
            .O(N__35787),
            .I(N__35770));
    InMux I__5269 (
            .O(N__35786),
            .I(N__35770));
    InMux I__5268 (
            .O(N__35785),
            .I(N__35770));
    InMux I__5267 (
            .O(N__35784),
            .I(N__35770));
    InMux I__5266 (
            .O(N__35783),
            .I(N__35761));
    InMux I__5265 (
            .O(N__35782),
            .I(N__35761));
    InMux I__5264 (
            .O(N__35781),
            .I(N__35761));
    InMux I__5263 (
            .O(N__35780),
            .I(N__35761));
    InMux I__5262 (
            .O(N__35779),
            .I(N__35758));
    LocalMux I__5261 (
            .O(N__35770),
            .I(N__35751));
    LocalMux I__5260 (
            .O(N__35761),
            .I(N__35751));
    LocalMux I__5259 (
            .O(N__35758),
            .I(N__35748));
    InMux I__5258 (
            .O(N__35757),
            .I(N__35745));
    InMux I__5257 (
            .O(N__35756),
            .I(N__35742));
    Span4Mux_v I__5256 (
            .O(N__35751),
            .I(N__35739));
    Span4Mux_v I__5255 (
            .O(N__35748),
            .I(N__35736));
    LocalMux I__5254 (
            .O(N__35745),
            .I(N__35733));
    LocalMux I__5253 (
            .O(N__35742),
            .I(N__35730));
    Odrv4 I__5252 (
            .O(N__35739),
            .I(\c0.n10 ));
    Odrv4 I__5251 (
            .O(N__35736),
            .I(\c0.n10 ));
    Odrv12 I__5250 (
            .O(N__35733),
            .I(\c0.n10 ));
    Odrv4 I__5249 (
            .O(N__35730),
            .I(\c0.n10 ));
    InMux I__5248 (
            .O(N__35721),
            .I(N__35716));
    InMux I__5247 (
            .O(N__35720),
            .I(N__35711));
    InMux I__5246 (
            .O(N__35719),
            .I(N__35711));
    LocalMux I__5245 (
            .O(N__35716),
            .I(N__35708));
    LocalMux I__5244 (
            .O(N__35711),
            .I(N__35705));
    Span4Mux_v I__5243 (
            .O(N__35708),
            .I(N__35702));
    Span4Mux_h I__5242 (
            .O(N__35705),
            .I(N__35699));
    Odrv4 I__5241 (
            .O(N__35702),
            .I(\c0.data_out_frame_29_7_N_1482_2 ));
    Odrv4 I__5240 (
            .O(N__35699),
            .I(\c0.data_out_frame_29_7_N_1482_2 ));
    CascadeMux I__5239 (
            .O(N__35694),
            .I(\c0.n14_adj_4727_cascade_ ));
    CascadeMux I__5238 (
            .O(N__35691),
            .I(N__35686));
    InMux I__5237 (
            .O(N__35690),
            .I(N__35683));
    InMux I__5236 (
            .O(N__35689),
            .I(N__35680));
    InMux I__5235 (
            .O(N__35686),
            .I(N__35677));
    LocalMux I__5234 (
            .O(N__35683),
            .I(N__35674));
    LocalMux I__5233 (
            .O(N__35680),
            .I(N__35669));
    LocalMux I__5232 (
            .O(N__35677),
            .I(N__35669));
    Odrv4 I__5231 (
            .O(N__35674),
            .I(\c0.n13056 ));
    Odrv12 I__5230 (
            .O(N__35669),
            .I(\c0.n13056 ));
    InMux I__5229 (
            .O(N__35664),
            .I(N__35659));
    InMux I__5228 (
            .O(N__35663),
            .I(N__35654));
    InMux I__5227 (
            .O(N__35662),
            .I(N__35654));
    LocalMux I__5226 (
            .O(N__35659),
            .I(N__35646));
    LocalMux I__5225 (
            .O(N__35654),
            .I(N__35646));
    InMux I__5224 (
            .O(N__35653),
            .I(N__35641));
    InMux I__5223 (
            .O(N__35652),
            .I(N__35641));
    InMux I__5222 (
            .O(N__35651),
            .I(N__35638));
    Span4Mux_v I__5221 (
            .O(N__35646),
            .I(N__35634));
    LocalMux I__5220 (
            .O(N__35641),
            .I(N__35631));
    LocalMux I__5219 (
            .O(N__35638),
            .I(N__35628));
    InMux I__5218 (
            .O(N__35637),
            .I(N__35625));
    Odrv4 I__5217 (
            .O(N__35634),
            .I(\c0.n63_adj_4235 ));
    Odrv12 I__5216 (
            .O(N__35631),
            .I(\c0.n63_adj_4235 ));
    Odrv4 I__5215 (
            .O(N__35628),
            .I(\c0.n63_adj_4235 ));
    LocalMux I__5214 (
            .O(N__35625),
            .I(\c0.n63_adj_4235 ));
    InMux I__5213 (
            .O(N__35616),
            .I(N__35611));
    InMux I__5212 (
            .O(N__35615),
            .I(N__35606));
    InMux I__5211 (
            .O(N__35614),
            .I(N__35606));
    LocalMux I__5210 (
            .O(N__35611),
            .I(N__35597));
    LocalMux I__5209 (
            .O(N__35606),
            .I(N__35597));
    InMux I__5208 (
            .O(N__35605),
            .I(N__35592));
    InMux I__5207 (
            .O(N__35604),
            .I(N__35592));
    InMux I__5206 (
            .O(N__35603),
            .I(N__35589));
    InMux I__5205 (
            .O(N__35602),
            .I(N__35586));
    Sp12to4 I__5204 (
            .O(N__35597),
            .I(N__35577));
    LocalMux I__5203 (
            .O(N__35592),
            .I(N__35577));
    LocalMux I__5202 (
            .O(N__35589),
            .I(N__35577));
    LocalMux I__5201 (
            .O(N__35586),
            .I(N__35577));
    Odrv12 I__5200 (
            .O(N__35577),
            .I(\c0.n63_adj_4238 ));
    CascadeMux I__5199 (
            .O(N__35574),
            .I(\c0.n2004_cascade_ ));
    CascadeMux I__5198 (
            .O(N__35571),
            .I(N__35568));
    InMux I__5197 (
            .O(N__35568),
            .I(N__35565));
    LocalMux I__5196 (
            .O(N__35565),
            .I(\c0.n28_adj_4565 ));
    CascadeMux I__5195 (
            .O(N__35562),
            .I(N__35558));
    CascadeMux I__5194 (
            .O(N__35561),
            .I(N__35555));
    InMux I__5193 (
            .O(N__35558),
            .I(N__35551));
    InMux I__5192 (
            .O(N__35555),
            .I(N__35546));
    InMux I__5191 (
            .O(N__35554),
            .I(N__35546));
    LocalMux I__5190 (
            .O(N__35551),
            .I(N__35539));
    LocalMux I__5189 (
            .O(N__35546),
            .I(N__35539));
    InMux I__5188 (
            .O(N__35545),
            .I(N__35536));
    InMux I__5187 (
            .O(N__35544),
            .I(N__35533));
    Span4Mux_v I__5186 (
            .O(N__35539),
            .I(N__35530));
    LocalMux I__5185 (
            .O(N__35536),
            .I(\c0.FRAME_MATCHER_state_16 ));
    LocalMux I__5184 (
            .O(N__35533),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv4 I__5183 (
            .O(N__35530),
            .I(\c0.FRAME_MATCHER_state_16 ));
    CascadeMux I__5182 (
            .O(N__35523),
            .I(\c0.n7570_cascade_ ));
    InMux I__5181 (
            .O(N__35520),
            .I(N__35514));
    InMux I__5180 (
            .O(N__35519),
            .I(N__35514));
    LocalMux I__5179 (
            .O(N__35514),
            .I(data_out_frame_6_4));
    InMux I__5178 (
            .O(N__35511),
            .I(N__35508));
    LocalMux I__5177 (
            .O(N__35508),
            .I(N__35504));
    InMux I__5176 (
            .O(N__35507),
            .I(N__35501));
    Span4Mux_v I__5175 (
            .O(N__35504),
            .I(N__35498));
    LocalMux I__5174 (
            .O(N__35501),
            .I(data_out_frame_7_4));
    Odrv4 I__5173 (
            .O(N__35498),
            .I(data_out_frame_7_4));
    CascadeMux I__5172 (
            .O(N__35493),
            .I(\c0.n13055_cascade_ ));
    CascadeMux I__5171 (
            .O(N__35490),
            .I(n13058_cascade_));
    InMux I__5170 (
            .O(N__35487),
            .I(N__35483));
    InMux I__5169 (
            .O(N__35486),
            .I(N__35480));
    LocalMux I__5168 (
            .O(N__35483),
            .I(N__35477));
    LocalMux I__5167 (
            .O(N__35480),
            .I(data_out_frame_7_6));
    Odrv4 I__5166 (
            .O(N__35477),
            .I(data_out_frame_7_6));
    InMux I__5165 (
            .O(N__35472),
            .I(N__35467));
    InMux I__5164 (
            .O(N__35471),
            .I(N__35464));
    InMux I__5163 (
            .O(N__35470),
            .I(N__35460));
    LocalMux I__5162 (
            .O(N__35467),
            .I(N__35457));
    LocalMux I__5161 (
            .O(N__35464),
            .I(N__35454));
    CascadeMux I__5160 (
            .O(N__35463),
            .I(N__35450));
    LocalMux I__5159 (
            .O(N__35460),
            .I(N__35443));
    Span4Mux_v I__5158 (
            .O(N__35457),
            .I(N__35443));
    Span4Mux_h I__5157 (
            .O(N__35454),
            .I(N__35443));
    InMux I__5156 (
            .O(N__35453),
            .I(N__35438));
    InMux I__5155 (
            .O(N__35450),
            .I(N__35438));
    Span4Mux_h I__5154 (
            .O(N__35443),
            .I(N__35435));
    LocalMux I__5153 (
            .O(N__35438),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__5152 (
            .O(N__35435),
            .I(\c0.FRAME_MATCHER_state_3 ));
    CascadeMux I__5151 (
            .O(N__35430),
            .I(N__35427));
    InMux I__5150 (
            .O(N__35427),
            .I(N__35424));
    LocalMux I__5149 (
            .O(N__35424),
            .I(N__35421));
    Odrv4 I__5148 (
            .O(N__35421),
            .I(\c0.n5_adj_4477 ));
    InMux I__5147 (
            .O(N__35418),
            .I(N__35412));
    InMux I__5146 (
            .O(N__35417),
            .I(N__35412));
    LocalMux I__5145 (
            .O(N__35412),
            .I(data_out_frame_13_4));
    InMux I__5144 (
            .O(N__35409),
            .I(N__35406));
    LocalMux I__5143 (
            .O(N__35406),
            .I(\c0.n11_adj_4669 ));
    InMux I__5142 (
            .O(N__35403),
            .I(N__35400));
    LocalMux I__5141 (
            .O(N__35400),
            .I(N__35396));
    InMux I__5140 (
            .O(N__35399),
            .I(N__35393));
    Span4Mux_h I__5139 (
            .O(N__35396),
            .I(N__35390));
    LocalMux I__5138 (
            .O(N__35393),
            .I(data_out_frame_8_5));
    Odrv4 I__5137 (
            .O(N__35390),
            .I(data_out_frame_8_5));
    InMux I__5136 (
            .O(N__35385),
            .I(N__35382));
    LocalMux I__5135 (
            .O(N__35382),
            .I(N__35378));
    InMux I__5134 (
            .O(N__35381),
            .I(N__35375));
    Span4Mux_v I__5133 (
            .O(N__35378),
            .I(N__35372));
    LocalMux I__5132 (
            .O(N__35375),
            .I(data_out_frame_7_5));
    Odrv4 I__5131 (
            .O(N__35372),
            .I(data_out_frame_7_5));
    CascadeMux I__5130 (
            .O(N__35367),
            .I(N__35364));
    InMux I__5129 (
            .O(N__35364),
            .I(N__35361));
    LocalMux I__5128 (
            .O(N__35361),
            .I(N__35357));
    InMux I__5127 (
            .O(N__35360),
            .I(N__35354));
    Span4Mux_v I__5126 (
            .O(N__35357),
            .I(N__35348));
    LocalMux I__5125 (
            .O(N__35354),
            .I(N__35348));
    InMux I__5124 (
            .O(N__35353),
            .I(N__35345));
    Span4Mux_h I__5123 (
            .O(N__35348),
            .I(N__35341));
    LocalMux I__5122 (
            .O(N__35345),
            .I(N__35338));
    InMux I__5121 (
            .O(N__35344),
            .I(N__35335));
    Span4Mux_v I__5120 (
            .O(N__35341),
            .I(N__35330));
    Span4Mux_h I__5119 (
            .O(N__35338),
            .I(N__35330));
    LocalMux I__5118 (
            .O(N__35335),
            .I(encoder1_position_25));
    Odrv4 I__5117 (
            .O(N__35330),
            .I(encoder1_position_25));
    InMux I__5116 (
            .O(N__35325),
            .I(N__35322));
    LocalMux I__5115 (
            .O(N__35322),
            .I(n2262));
    InMux I__5114 (
            .O(N__35319),
            .I(N__35315));
    CascadeMux I__5113 (
            .O(N__35318),
            .I(N__35312));
    LocalMux I__5112 (
            .O(N__35315),
            .I(N__35309));
    InMux I__5111 (
            .O(N__35312),
            .I(N__35306));
    Span4Mux_h I__5110 (
            .O(N__35309),
            .I(N__35303));
    LocalMux I__5109 (
            .O(N__35306),
            .I(data_out_frame_10_6));
    Odrv4 I__5108 (
            .O(N__35303),
            .I(data_out_frame_10_6));
    CascadeMux I__5107 (
            .O(N__35298),
            .I(N__35294));
    CascadeMux I__5106 (
            .O(N__35297),
            .I(N__35291));
    InMux I__5105 (
            .O(N__35294),
            .I(N__35288));
    InMux I__5104 (
            .O(N__35291),
            .I(N__35280));
    LocalMux I__5103 (
            .O(N__35288),
            .I(N__35277));
    InMux I__5102 (
            .O(N__35287),
            .I(N__35274));
    InMux I__5101 (
            .O(N__35286),
            .I(N__35269));
    InMux I__5100 (
            .O(N__35285),
            .I(N__35269));
    InMux I__5099 (
            .O(N__35284),
            .I(N__35265));
    CascadeMux I__5098 (
            .O(N__35283),
            .I(N__35262));
    LocalMux I__5097 (
            .O(N__35280),
            .I(N__35258));
    Span4Mux_v I__5096 (
            .O(N__35277),
            .I(N__35251));
    LocalMux I__5095 (
            .O(N__35274),
            .I(N__35251));
    LocalMux I__5094 (
            .O(N__35269),
            .I(N__35251));
    InMux I__5093 (
            .O(N__35268),
            .I(N__35248));
    LocalMux I__5092 (
            .O(N__35265),
            .I(N__35245));
    InMux I__5091 (
            .O(N__35262),
            .I(N__35240));
    InMux I__5090 (
            .O(N__35261),
            .I(N__35240));
    Span4Mux_v I__5089 (
            .O(N__35258),
            .I(N__35235));
    Span4Mux_v I__5088 (
            .O(N__35251),
            .I(N__35235));
    LocalMux I__5087 (
            .O(N__35248),
            .I(encoder1_position_4));
    Odrv12 I__5086 (
            .O(N__35245),
            .I(encoder1_position_4));
    LocalMux I__5085 (
            .O(N__35240),
            .I(encoder1_position_4));
    Odrv4 I__5084 (
            .O(N__35235),
            .I(encoder1_position_4));
    InMux I__5083 (
            .O(N__35226),
            .I(N__35222));
    InMux I__5082 (
            .O(N__35225),
            .I(N__35219));
    LocalMux I__5081 (
            .O(N__35222),
            .I(N__35216));
    LocalMux I__5080 (
            .O(N__35219),
            .I(data_out_frame_8_0));
    Odrv4 I__5079 (
            .O(N__35216),
            .I(data_out_frame_8_0));
    CascadeMux I__5078 (
            .O(N__35211),
            .I(N__35208));
    InMux I__5077 (
            .O(N__35208),
            .I(N__35204));
    InMux I__5076 (
            .O(N__35207),
            .I(N__35201));
    LocalMux I__5075 (
            .O(N__35204),
            .I(N__35198));
    LocalMux I__5074 (
            .O(N__35201),
            .I(N__35195));
    Span4Mux_v I__5073 (
            .O(N__35198),
            .I(N__35189));
    Span4Mux_h I__5072 (
            .O(N__35195),
            .I(N__35189));
    InMux I__5071 (
            .O(N__35194),
            .I(N__35185));
    Span4Mux_v I__5070 (
            .O(N__35189),
            .I(N__35182));
    InMux I__5069 (
            .O(N__35188),
            .I(N__35179));
    LocalMux I__5068 (
            .O(N__35185),
            .I(encoder1_position_17));
    Odrv4 I__5067 (
            .O(N__35182),
            .I(encoder1_position_17));
    LocalMux I__5066 (
            .O(N__35179),
            .I(encoder1_position_17));
    InMux I__5065 (
            .O(N__35172),
            .I(N__35169));
    LocalMux I__5064 (
            .O(N__35169),
            .I(\c0.n16_adj_4233 ));
    CascadeMux I__5063 (
            .O(N__35166),
            .I(N__35163));
    InMux I__5062 (
            .O(N__35163),
            .I(N__35159));
    InMux I__5061 (
            .O(N__35162),
            .I(N__35156));
    LocalMux I__5060 (
            .O(N__35159),
            .I(N__35153));
    LocalMux I__5059 (
            .O(N__35156),
            .I(data_out_frame_11_7));
    Odrv12 I__5058 (
            .O(N__35153),
            .I(data_out_frame_11_7));
    InMux I__5057 (
            .O(N__35148),
            .I(N__35144));
    InMux I__5056 (
            .O(N__35147),
            .I(N__35141));
    LocalMux I__5055 (
            .O(N__35144),
            .I(N__35138));
    LocalMux I__5054 (
            .O(N__35141),
            .I(data_out_frame_13_5));
    Odrv12 I__5053 (
            .O(N__35138),
            .I(data_out_frame_13_5));
    InMux I__5052 (
            .O(N__35133),
            .I(N__35129));
    InMux I__5051 (
            .O(N__35132),
            .I(N__35126));
    LocalMux I__5050 (
            .O(N__35129),
            .I(N__35123));
    LocalMux I__5049 (
            .O(N__35126),
            .I(N__35120));
    Span4Mux_v I__5048 (
            .O(N__35123),
            .I(N__35117));
    Span4Mux_v I__5047 (
            .O(N__35120),
            .I(N__35113));
    Span4Mux_v I__5046 (
            .O(N__35117),
            .I(N__35108));
    InMux I__5045 (
            .O(N__35116),
            .I(N__35105));
    Span4Mux_v I__5044 (
            .O(N__35113),
            .I(N__35102));
    InMux I__5043 (
            .O(N__35112),
            .I(N__35099));
    InMux I__5042 (
            .O(N__35111),
            .I(N__35096));
    Odrv4 I__5041 (
            .O(N__35108),
            .I(encoder1_position_11));
    LocalMux I__5040 (
            .O(N__35105),
            .I(encoder1_position_11));
    Odrv4 I__5039 (
            .O(N__35102),
            .I(encoder1_position_11));
    LocalMux I__5038 (
            .O(N__35099),
            .I(encoder1_position_11));
    LocalMux I__5037 (
            .O(N__35096),
            .I(encoder1_position_11));
    InMux I__5036 (
            .O(N__35085),
            .I(N__35082));
    LocalMux I__5035 (
            .O(N__35082),
            .I(N__35079));
    Span4Mux_v I__5034 (
            .O(N__35079),
            .I(N__35075));
    InMux I__5033 (
            .O(N__35078),
            .I(N__35072));
    Span4Mux_h I__5032 (
            .O(N__35075),
            .I(N__35069));
    LocalMux I__5031 (
            .O(N__35072),
            .I(data_out_frame_12_3));
    Odrv4 I__5030 (
            .O(N__35069),
            .I(data_out_frame_12_3));
    CascadeMux I__5029 (
            .O(N__35064),
            .I(N__35061));
    InMux I__5028 (
            .O(N__35061),
            .I(N__35057));
    InMux I__5027 (
            .O(N__35060),
            .I(N__35054));
    LocalMux I__5026 (
            .O(N__35057),
            .I(N__35051));
    LocalMux I__5025 (
            .O(N__35054),
            .I(data_out_frame_12_2));
    Odrv4 I__5024 (
            .O(N__35051),
            .I(data_out_frame_12_2));
    InMux I__5023 (
            .O(N__35046),
            .I(N__35043));
    LocalMux I__5022 (
            .O(N__35043),
            .I(n2281));
    InMux I__5021 (
            .O(N__35040),
            .I(N__35035));
    CascadeMux I__5020 (
            .O(N__35039),
            .I(N__35029));
    CascadeMux I__5019 (
            .O(N__35038),
            .I(N__35026));
    LocalMux I__5018 (
            .O(N__35035),
            .I(N__35023));
    InMux I__5017 (
            .O(N__35034),
            .I(N__35018));
    InMux I__5016 (
            .O(N__35033),
            .I(N__35018));
    InMux I__5015 (
            .O(N__35032),
            .I(N__35013));
    InMux I__5014 (
            .O(N__35029),
            .I(N__35013));
    InMux I__5013 (
            .O(N__35026),
            .I(N__35010));
    Span4Mux_h I__5012 (
            .O(N__35023),
            .I(N__35007));
    LocalMux I__5011 (
            .O(N__35018),
            .I(N__35004));
    LocalMux I__5010 (
            .O(N__35013),
            .I(encoder1_position_10));
    LocalMux I__5009 (
            .O(N__35010),
            .I(encoder1_position_10));
    Odrv4 I__5008 (
            .O(N__35007),
            .I(encoder1_position_10));
    Odrv12 I__5007 (
            .O(N__35004),
            .I(encoder1_position_10));
    InMux I__5006 (
            .O(N__34995),
            .I(N__34992));
    LocalMux I__5005 (
            .O(N__34992),
            .I(N__34988));
    InMux I__5004 (
            .O(N__34991),
            .I(N__34985));
    Span4Mux_h I__5003 (
            .O(N__34988),
            .I(N__34982));
    LocalMux I__5002 (
            .O(N__34985),
            .I(data_out_frame_5_6));
    Odrv4 I__5001 (
            .O(N__34982),
            .I(data_out_frame_5_6));
    InMux I__5000 (
            .O(N__34977),
            .I(N__34970));
    InMux I__4999 (
            .O(N__34976),
            .I(N__34970));
    CascadeMux I__4998 (
            .O(N__34975),
            .I(N__34967));
    LocalMux I__4997 (
            .O(N__34970),
            .I(N__34964));
    InMux I__4996 (
            .O(N__34967),
            .I(N__34960));
    Span4Mux_h I__4995 (
            .O(N__34964),
            .I(N__34956));
    InMux I__4994 (
            .O(N__34963),
            .I(N__34953));
    LocalMux I__4993 (
            .O(N__34960),
            .I(N__34950));
    InMux I__4992 (
            .O(N__34959),
            .I(N__34947));
    Span4Mux_v I__4991 (
            .O(N__34956),
            .I(N__34944));
    LocalMux I__4990 (
            .O(N__34953),
            .I(encoder1_position_15));
    Odrv4 I__4989 (
            .O(N__34950),
            .I(encoder1_position_15));
    LocalMux I__4988 (
            .O(N__34947),
            .I(encoder1_position_15));
    Odrv4 I__4987 (
            .O(N__34944),
            .I(encoder1_position_15));
    InMux I__4986 (
            .O(N__34935),
            .I(N__34932));
    LocalMux I__4985 (
            .O(N__34932),
            .I(N__34929));
    Span4Mux_v I__4984 (
            .O(N__34929),
            .I(N__34925));
    InMux I__4983 (
            .O(N__34928),
            .I(N__34922));
    Span4Mux_h I__4982 (
            .O(N__34925),
            .I(N__34919));
    LocalMux I__4981 (
            .O(N__34922),
            .I(data_out_frame_12_7));
    Odrv4 I__4980 (
            .O(N__34919),
            .I(data_out_frame_12_7));
    InMux I__4979 (
            .O(N__34914),
            .I(N__34911));
    LocalMux I__4978 (
            .O(N__34911),
            .I(n2263));
    CascadeMux I__4977 (
            .O(N__34908),
            .I(N__34905));
    InMux I__4976 (
            .O(N__34905),
            .I(N__34902));
    LocalMux I__4975 (
            .O(N__34902),
            .I(n2264));
    CascadeMux I__4974 (
            .O(N__34899),
            .I(N__34896));
    InMux I__4973 (
            .O(N__34896),
            .I(N__34892));
    InMux I__4972 (
            .O(N__34895),
            .I(N__34889));
    LocalMux I__4971 (
            .O(N__34892),
            .I(N__34885));
    LocalMux I__4970 (
            .O(N__34889),
            .I(N__34881));
    InMux I__4969 (
            .O(N__34888),
            .I(N__34878));
    Span4Mux_v I__4968 (
            .O(N__34885),
            .I(N__34875));
    InMux I__4967 (
            .O(N__34884),
            .I(N__34872));
    Span4Mux_v I__4966 (
            .O(N__34881),
            .I(N__34869));
    LocalMux I__4965 (
            .O(N__34878),
            .I(encoder1_position_27));
    Odrv4 I__4964 (
            .O(N__34875),
            .I(encoder1_position_27));
    LocalMux I__4963 (
            .O(N__34872),
            .I(encoder1_position_27));
    Odrv4 I__4962 (
            .O(N__34869),
            .I(encoder1_position_27));
    CascadeMux I__4961 (
            .O(N__34860),
            .I(N__34857));
    InMux I__4960 (
            .O(N__34857),
            .I(N__34853));
    InMux I__4959 (
            .O(N__34856),
            .I(N__34850));
    LocalMux I__4958 (
            .O(N__34853),
            .I(N__34847));
    LocalMux I__4957 (
            .O(N__34850),
            .I(data_out_frame_5_3));
    Odrv4 I__4956 (
            .O(N__34847),
            .I(data_out_frame_5_3));
    InMux I__4955 (
            .O(N__34842),
            .I(N__34838));
    InMux I__4954 (
            .O(N__34841),
            .I(N__34835));
    LocalMux I__4953 (
            .O(N__34838),
            .I(N__34832));
    LocalMux I__4952 (
            .O(N__34835),
            .I(data_out_frame_7_1));
    Odrv4 I__4951 (
            .O(N__34832),
            .I(data_out_frame_7_1));
    InMux I__4950 (
            .O(N__34827),
            .I(N__34824));
    LocalMux I__4949 (
            .O(N__34824),
            .I(n2270));
    InMux I__4948 (
            .O(N__34821),
            .I(N__34818));
    LocalMux I__4947 (
            .O(N__34818),
            .I(N__34811));
    InMux I__4946 (
            .O(N__34817),
            .I(N__34806));
    InMux I__4945 (
            .O(N__34816),
            .I(N__34806));
    InMux I__4944 (
            .O(N__34815),
            .I(N__34800));
    InMux I__4943 (
            .O(N__34814),
            .I(N__34800));
    Span4Mux_v I__4942 (
            .O(N__34811),
            .I(N__34795));
    LocalMux I__4941 (
            .O(N__34806),
            .I(N__34795));
    InMux I__4940 (
            .O(N__34805),
            .I(N__34792));
    LocalMux I__4939 (
            .O(N__34800),
            .I(\c0.n13395 ));
    Odrv4 I__4938 (
            .O(N__34795),
            .I(\c0.n13395 ));
    LocalMux I__4937 (
            .O(N__34792),
            .I(\c0.n13395 ));
    CascadeMux I__4936 (
            .O(N__34785),
            .I(N__34782));
    InMux I__4935 (
            .O(N__34782),
            .I(N__34777));
    InMux I__4934 (
            .O(N__34781),
            .I(N__34772));
    CascadeMux I__4933 (
            .O(N__34780),
            .I(N__34769));
    LocalMux I__4932 (
            .O(N__34777),
            .I(N__34766));
    InMux I__4931 (
            .O(N__34776),
            .I(N__34762));
    InMux I__4930 (
            .O(N__34775),
            .I(N__34759));
    LocalMux I__4929 (
            .O(N__34772),
            .I(N__34756));
    InMux I__4928 (
            .O(N__34769),
            .I(N__34753));
    Span4Mux_h I__4927 (
            .O(N__34766),
            .I(N__34750));
    InMux I__4926 (
            .O(N__34765),
            .I(N__34747));
    LocalMux I__4925 (
            .O(N__34762),
            .I(N__34741));
    LocalMux I__4924 (
            .O(N__34759),
            .I(N__34741));
    Span4Mux_v I__4923 (
            .O(N__34756),
            .I(N__34738));
    LocalMux I__4922 (
            .O(N__34753),
            .I(N__34734));
    Span4Mux_v I__4921 (
            .O(N__34750),
            .I(N__34729));
    LocalMux I__4920 (
            .O(N__34747),
            .I(N__34729));
    InMux I__4919 (
            .O(N__34746),
            .I(N__34726));
    Span4Mux_v I__4918 (
            .O(N__34741),
            .I(N__34721));
    Span4Mux_h I__4917 (
            .O(N__34738),
            .I(N__34721));
    InMux I__4916 (
            .O(N__34737),
            .I(N__34718));
    Span4Mux_h I__4915 (
            .O(N__34734),
            .I(N__34715));
    Span4Mux_v I__4914 (
            .O(N__34729),
            .I(N__34712));
    LocalMux I__4913 (
            .O(N__34726),
            .I(N__34709));
    Span4Mux_h I__4912 (
            .O(N__34721),
            .I(N__34706));
    LocalMux I__4911 (
            .O(N__34718),
            .I(encoder1_position_1));
    Odrv4 I__4910 (
            .O(N__34715),
            .I(encoder1_position_1));
    Odrv4 I__4909 (
            .O(N__34712),
            .I(encoder1_position_1));
    Odrv4 I__4908 (
            .O(N__34709),
            .I(encoder1_position_1));
    Odrv4 I__4907 (
            .O(N__34706),
            .I(encoder1_position_1));
    InMux I__4906 (
            .O(N__34695),
            .I(N__34692));
    LocalMux I__4905 (
            .O(N__34692),
            .I(N__34688));
    InMux I__4904 (
            .O(N__34691),
            .I(N__34685));
    Span4Mux_h I__4903 (
            .O(N__34688),
            .I(N__34682));
    LocalMux I__4902 (
            .O(N__34685),
            .I(data_out_frame_9_0));
    Odrv4 I__4901 (
            .O(N__34682),
            .I(data_out_frame_9_0));
    InMux I__4900 (
            .O(N__34677),
            .I(N__34674));
    LocalMux I__4899 (
            .O(N__34674),
            .I(N__34670));
    InMux I__4898 (
            .O(N__34673),
            .I(N__34667));
    Span4Mux_v I__4897 (
            .O(N__34670),
            .I(N__34664));
    LocalMux I__4896 (
            .O(N__34667),
            .I(data_out_frame_5_4));
    Odrv4 I__4895 (
            .O(N__34664),
            .I(data_out_frame_5_4));
    CascadeMux I__4894 (
            .O(N__34659),
            .I(N__34656));
    InMux I__4893 (
            .O(N__34656),
            .I(N__34651));
    CascadeMux I__4892 (
            .O(N__34655),
            .I(N__34646));
    InMux I__4891 (
            .O(N__34654),
            .I(N__34643));
    LocalMux I__4890 (
            .O(N__34651),
            .I(N__34640));
    InMux I__4889 (
            .O(N__34650),
            .I(N__34637));
    InMux I__4888 (
            .O(N__34649),
            .I(N__34634));
    InMux I__4887 (
            .O(N__34646),
            .I(N__34631));
    LocalMux I__4886 (
            .O(N__34643),
            .I(N__34628));
    Span4Mux_h I__4885 (
            .O(N__34640),
            .I(N__34623));
    LocalMux I__4884 (
            .O(N__34637),
            .I(N__34623));
    LocalMux I__4883 (
            .O(N__34634),
            .I(encoder1_position_22));
    LocalMux I__4882 (
            .O(N__34631),
            .I(encoder1_position_22));
    Odrv4 I__4881 (
            .O(N__34628),
            .I(encoder1_position_22));
    Odrv4 I__4880 (
            .O(N__34623),
            .I(encoder1_position_22));
    CascadeMux I__4879 (
            .O(N__34614),
            .I(N__34611));
    InMux I__4878 (
            .O(N__34611),
            .I(N__34606));
    InMux I__4877 (
            .O(N__34610),
            .I(N__34603));
    InMux I__4876 (
            .O(N__34609),
            .I(N__34599));
    LocalMux I__4875 (
            .O(N__34606),
            .I(N__34596));
    LocalMux I__4874 (
            .O(N__34603),
            .I(N__34590));
    InMux I__4873 (
            .O(N__34602),
            .I(N__34587));
    LocalMux I__4872 (
            .O(N__34599),
            .I(N__34584));
    Span4Mux_h I__4871 (
            .O(N__34596),
            .I(N__34581));
    InMux I__4870 (
            .O(N__34595),
            .I(N__34578));
    InMux I__4869 (
            .O(N__34594),
            .I(N__34575));
    InMux I__4868 (
            .O(N__34593),
            .I(N__34572));
    Span12Mux_s7_v I__4867 (
            .O(N__34590),
            .I(N__34569));
    LocalMux I__4866 (
            .O(N__34587),
            .I(N__34566));
    Span4Mux_h I__4865 (
            .O(N__34584),
            .I(N__34561));
    Span4Mux_h I__4864 (
            .O(N__34581),
            .I(N__34561));
    LocalMux I__4863 (
            .O(N__34578),
            .I(encoder1_position_7));
    LocalMux I__4862 (
            .O(N__34575),
            .I(encoder1_position_7));
    LocalMux I__4861 (
            .O(N__34572),
            .I(encoder1_position_7));
    Odrv12 I__4860 (
            .O(N__34569),
            .I(encoder1_position_7));
    Odrv4 I__4859 (
            .O(N__34566),
            .I(encoder1_position_7));
    Odrv4 I__4858 (
            .O(N__34561),
            .I(encoder1_position_7));
    InMux I__4857 (
            .O(N__34548),
            .I(N__34545));
    LocalMux I__4856 (
            .O(N__34545),
            .I(N__34541));
    InMux I__4855 (
            .O(N__34544),
            .I(N__34538));
    Span4Mux_h I__4854 (
            .O(N__34541),
            .I(N__34535));
    LocalMux I__4853 (
            .O(N__34538),
            .I(data_out_frame_7_2));
    Odrv4 I__4852 (
            .O(N__34535),
            .I(data_out_frame_7_2));
    InMux I__4851 (
            .O(N__34530),
            .I(N__34527));
    LocalMux I__4850 (
            .O(N__34527),
            .I(N__34524));
    Span4Mux_v I__4849 (
            .O(N__34524),
            .I(N__34521));
    Odrv4 I__4848 (
            .O(N__34521),
            .I(\c0.data_out_frame_29_0 ));
    InMux I__4847 (
            .O(N__34518),
            .I(N__34515));
    LocalMux I__4846 (
            .O(N__34515),
            .I(\c0.data_out_frame_28_0 ));
    InMux I__4845 (
            .O(N__34512),
            .I(N__34509));
    LocalMux I__4844 (
            .O(N__34509),
            .I(N__34506));
    Span12Mux_v I__4843 (
            .O(N__34506),
            .I(N__34503));
    Odrv12 I__4842 (
            .O(N__34503),
            .I(\c0.n26_adj_4570 ));
    CascadeMux I__4841 (
            .O(N__34500),
            .I(\c0.n10529_cascade_ ));
    CascadeMux I__4840 (
            .O(N__34497),
            .I(\c0.n22489_cascade_ ));
    CascadeMux I__4839 (
            .O(N__34494),
            .I(\c0.n21416_cascade_ ));
    InMux I__4838 (
            .O(N__34491),
            .I(N__34488));
    LocalMux I__4837 (
            .O(N__34488),
            .I(N__34485));
    Span4Mux_v I__4836 (
            .O(N__34485),
            .I(N__34482));
    Odrv4 I__4835 (
            .O(N__34482),
            .I(\c0.n24530 ));
    CascadeMux I__4834 (
            .O(N__34479),
            .I(\c0.n22671_cascade_ ));
    InMux I__4833 (
            .O(N__34476),
            .I(N__34473));
    LocalMux I__4832 (
            .O(N__34473),
            .I(\c0.n20230 ));
    CascadeMux I__4831 (
            .O(N__34470),
            .I(\c0.n20230_cascade_ ));
    InMux I__4830 (
            .O(N__34467),
            .I(N__34464));
    LocalMux I__4829 (
            .O(N__34464),
            .I(N__34461));
    Sp12to4 I__4828 (
            .O(N__34461),
            .I(N__34458));
    Odrv12 I__4827 (
            .O(N__34458),
            .I(\c0.data_out_frame_29_5 ));
    InMux I__4826 (
            .O(N__34455),
            .I(N__34452));
    LocalMux I__4825 (
            .O(N__34452),
            .I(\c0.n21457 ));
    InMux I__4824 (
            .O(N__34449),
            .I(N__34445));
    InMux I__4823 (
            .O(N__34448),
            .I(N__34442));
    LocalMux I__4822 (
            .O(N__34445),
            .I(\c0.n21489 ));
    LocalMux I__4821 (
            .O(N__34442),
            .I(\c0.n21489 ));
    InMux I__4820 (
            .O(N__34437),
            .I(N__34434));
    LocalMux I__4819 (
            .O(N__34434),
            .I(N__34429));
    InMux I__4818 (
            .O(N__34433),
            .I(N__34426));
    CascadeMux I__4817 (
            .O(N__34432),
            .I(N__34422));
    Span4Mux_v I__4816 (
            .O(N__34429),
            .I(N__34416));
    LocalMux I__4815 (
            .O(N__34426),
            .I(N__34416));
    InMux I__4814 (
            .O(N__34425),
            .I(N__34413));
    InMux I__4813 (
            .O(N__34422),
            .I(N__34410));
    InMux I__4812 (
            .O(N__34421),
            .I(N__34407));
    Span4Mux_v I__4811 (
            .O(N__34416),
            .I(N__34404));
    LocalMux I__4810 (
            .O(N__34413),
            .I(N__34401));
    LocalMux I__4809 (
            .O(N__34410),
            .I(N__34398));
    LocalMux I__4808 (
            .O(N__34407),
            .I(encoder1_position_6));
    Odrv4 I__4807 (
            .O(N__34404),
            .I(encoder1_position_6));
    Odrv4 I__4806 (
            .O(N__34401),
            .I(encoder1_position_6));
    Odrv4 I__4805 (
            .O(N__34398),
            .I(encoder1_position_6));
    InMux I__4804 (
            .O(N__34389),
            .I(N__34386));
    LocalMux I__4803 (
            .O(N__34386),
            .I(N__34383));
    Odrv4 I__4802 (
            .O(N__34383),
            .I(\c0.n20461 ));
    CascadeMux I__4801 (
            .O(N__34380),
            .I(\c0.n21330_cascade_ ));
    InMux I__4800 (
            .O(N__34377),
            .I(N__34374));
    LocalMux I__4799 (
            .O(N__34374),
            .I(\c0.n6_adj_4331 ));
    InMux I__4798 (
            .O(N__34371),
            .I(N__34368));
    LocalMux I__4797 (
            .O(N__34368),
            .I(N__34364));
    InMux I__4796 (
            .O(N__34367),
            .I(N__34361));
    Odrv4 I__4795 (
            .O(N__34364),
            .I(\c0.n22414 ));
    LocalMux I__4794 (
            .O(N__34361),
            .I(\c0.n22414 ));
    InMux I__4793 (
            .O(N__34356),
            .I(N__34353));
    LocalMux I__4792 (
            .O(N__34353),
            .I(N__34349));
    InMux I__4791 (
            .O(N__34352),
            .I(N__34346));
    Span4Mux_v I__4790 (
            .O(N__34349),
            .I(N__34339));
    LocalMux I__4789 (
            .O(N__34346),
            .I(N__34339));
    InMux I__4788 (
            .O(N__34345),
            .I(N__34336));
    InMux I__4787 (
            .O(N__34344),
            .I(N__34333));
    Span4Mux_h I__4786 (
            .O(N__34339),
            .I(N__34330));
    LocalMux I__4785 (
            .O(N__34336),
            .I(n21307));
    LocalMux I__4784 (
            .O(N__34333),
            .I(n21307));
    Odrv4 I__4783 (
            .O(N__34330),
            .I(n21307));
    CascadeMux I__4782 (
            .O(N__34323),
            .I(\c0.n6_adj_4215_cascade_ ));
    InMux I__4781 (
            .O(N__34320),
            .I(N__34317));
    LocalMux I__4780 (
            .O(N__34317),
            .I(N__34313));
    InMux I__4779 (
            .O(N__34316),
            .I(N__34310));
    Odrv4 I__4778 (
            .O(N__34313),
            .I(\c0.n22268 ));
    LocalMux I__4777 (
            .O(N__34310),
            .I(\c0.n22268 ));
    CascadeMux I__4776 (
            .O(N__34305),
            .I(N__34302));
    InMux I__4775 (
            .O(N__34302),
            .I(N__34299));
    LocalMux I__4774 (
            .O(N__34299),
            .I(N__34296));
    Span4Mux_h I__4773 (
            .O(N__34296),
            .I(N__34293));
    Span4Mux_h I__4772 (
            .O(N__34293),
            .I(N__34290));
    Odrv4 I__4771 (
            .O(N__34290),
            .I(\c0.n5_adj_4660 ));
    InMux I__4770 (
            .O(N__34287),
            .I(N__34284));
    LocalMux I__4769 (
            .O(N__34284),
            .I(N__34281));
    Span12Mux_v I__4768 (
            .O(N__34281),
            .I(N__34278));
    Odrv12 I__4767 (
            .O(N__34278),
            .I(\c0.n6_adj_4659 ));
    InMux I__4766 (
            .O(N__34275),
            .I(N__34272));
    LocalMux I__4765 (
            .O(N__34272),
            .I(N__34269));
    Span4Mux_v I__4764 (
            .O(N__34269),
            .I(N__34266));
    Odrv4 I__4763 (
            .O(N__34266),
            .I(\c0.n24755 ));
    InMux I__4762 (
            .O(N__34263),
            .I(N__34259));
    InMux I__4761 (
            .O(N__34262),
            .I(N__34256));
    LocalMux I__4760 (
            .O(N__34259),
            .I(N__34251));
    LocalMux I__4759 (
            .O(N__34256),
            .I(N__34251));
    Span4Mux_h I__4758 (
            .O(N__34251),
            .I(N__34248));
    Odrv4 I__4757 (
            .O(N__34248),
            .I(\c0.n22330 ));
    CascadeMux I__4756 (
            .O(N__34245),
            .I(\c0.n19_adj_4693_cascade_ ));
    CascadeMux I__4755 (
            .O(N__34242),
            .I(\c0.n6_adj_4691_cascade_ ));
    InMux I__4754 (
            .O(N__34239),
            .I(N__34236));
    LocalMux I__4753 (
            .O(N__34236),
            .I(\c0.n21_adj_4692 ));
    InMux I__4752 (
            .O(N__34233),
            .I(N__34230));
    LocalMux I__4751 (
            .O(N__34230),
            .I(N__34227));
    Span4Mux_h I__4750 (
            .O(N__34227),
            .I(N__34224));
    Span4Mux_v I__4749 (
            .O(N__34224),
            .I(N__34221));
    Odrv4 I__4748 (
            .O(N__34221),
            .I(n2274));
    InMux I__4747 (
            .O(N__34218),
            .I(N__34215));
    LocalMux I__4746 (
            .O(N__34215),
            .I(N__34212));
    Span4Mux_v I__4745 (
            .O(N__34212),
            .I(N__34209));
    Odrv4 I__4744 (
            .O(N__34209),
            .I(n2283));
    InMux I__4743 (
            .O(N__34206),
            .I(N__34202));
    InMux I__4742 (
            .O(N__34205),
            .I(N__34199));
    LocalMux I__4741 (
            .O(N__34202),
            .I(N__34196));
    LocalMux I__4740 (
            .O(N__34199),
            .I(\c0.n22656 ));
    Odrv4 I__4739 (
            .O(N__34196),
            .I(\c0.n22656 ));
    CascadeMux I__4738 (
            .O(N__34191),
            .I(N__34188));
    InMux I__4737 (
            .O(N__34188),
            .I(N__34185));
    LocalMux I__4736 (
            .O(N__34185),
            .I(N__34182));
    Span4Mux_h I__4735 (
            .O(N__34182),
            .I(N__34178));
    InMux I__4734 (
            .O(N__34181),
            .I(N__34175));
    Odrv4 I__4733 (
            .O(N__34178),
            .I(\c0.n22800 ));
    LocalMux I__4732 (
            .O(N__34175),
            .I(\c0.n22800 ));
    InMux I__4731 (
            .O(N__34170),
            .I(N__34167));
    LocalMux I__4730 (
            .O(N__34167),
            .I(N__34164));
    Odrv12 I__4729 (
            .O(N__34164),
            .I(\c0.n10_adj_4339 ));
    CascadeMux I__4728 (
            .O(N__34161),
            .I(\c0.n14_adj_4338_cascade_ ));
    CascadeMux I__4727 (
            .O(N__34158),
            .I(\c0.n20461_cascade_ ));
    InMux I__4726 (
            .O(N__34155),
            .I(N__34151));
    InMux I__4725 (
            .O(N__34154),
            .I(N__34147));
    LocalMux I__4724 (
            .O(N__34151),
            .I(N__34144));
    InMux I__4723 (
            .O(N__34150),
            .I(N__34141));
    LocalMux I__4722 (
            .O(N__34147),
            .I(N__34138));
    Span4Mux_v I__4721 (
            .O(N__34144),
            .I(N__34133));
    LocalMux I__4720 (
            .O(N__34141),
            .I(N__34130));
    Span4Mux_h I__4719 (
            .O(N__34138),
            .I(N__34127));
    InMux I__4718 (
            .O(N__34137),
            .I(N__34122));
    InMux I__4717 (
            .O(N__34136),
            .I(N__34122));
    Odrv4 I__4716 (
            .O(N__34133),
            .I(\c0.n20388 ));
    Odrv4 I__4715 (
            .O(N__34130),
            .I(\c0.n20388 ));
    Odrv4 I__4714 (
            .O(N__34127),
            .I(\c0.n20388 ));
    LocalMux I__4713 (
            .O(N__34122),
            .I(\c0.n20388 ));
    InMux I__4712 (
            .O(N__34113),
            .I(N__34110));
    LocalMux I__4711 (
            .O(N__34110),
            .I(N__34106));
    InMux I__4710 (
            .O(N__34109),
            .I(N__34103));
    Odrv4 I__4709 (
            .O(N__34106),
            .I(\c0.n22408 ));
    LocalMux I__4708 (
            .O(N__34103),
            .I(\c0.n22408 ));
    CascadeMux I__4707 (
            .O(N__34098),
            .I(N__34095));
    InMux I__4706 (
            .O(N__34095),
            .I(N__34092));
    LocalMux I__4705 (
            .O(N__34092),
            .I(N__34087));
    InMux I__4704 (
            .O(N__34091),
            .I(N__34084));
    InMux I__4703 (
            .O(N__34090),
            .I(N__34080));
    Span4Mux_v I__4702 (
            .O(N__34087),
            .I(N__34075));
    LocalMux I__4701 (
            .O(N__34084),
            .I(N__34075));
    CascadeMux I__4700 (
            .O(N__34083),
            .I(N__34070));
    LocalMux I__4699 (
            .O(N__34080),
            .I(N__34067));
    Span4Mux_h I__4698 (
            .O(N__34075),
            .I(N__34064));
    InMux I__4697 (
            .O(N__34074),
            .I(N__34061));
    CascadeMux I__4696 (
            .O(N__34073),
            .I(N__34058));
    InMux I__4695 (
            .O(N__34070),
            .I(N__34055));
    Sp12to4 I__4694 (
            .O(N__34067),
            .I(N__34050));
    Sp12to4 I__4693 (
            .O(N__34064),
            .I(N__34050));
    LocalMux I__4692 (
            .O(N__34061),
            .I(N__34047));
    InMux I__4691 (
            .O(N__34058),
            .I(N__34044));
    LocalMux I__4690 (
            .O(N__34055),
            .I(N__34041));
    Span12Mux_v I__4689 (
            .O(N__34050),
            .I(N__34038));
    Odrv4 I__4688 (
            .O(N__34047),
            .I(encoder1_position_16));
    LocalMux I__4687 (
            .O(N__34044),
            .I(encoder1_position_16));
    Odrv4 I__4686 (
            .O(N__34041),
            .I(encoder1_position_16));
    Odrv12 I__4685 (
            .O(N__34038),
            .I(encoder1_position_16));
    InMux I__4684 (
            .O(N__34029),
            .I(N__34024));
    InMux I__4683 (
            .O(N__34028),
            .I(N__34021));
    InMux I__4682 (
            .O(N__34027),
            .I(N__34018));
    LocalMux I__4681 (
            .O(N__34024),
            .I(\c0.n20449 ));
    LocalMux I__4680 (
            .O(N__34021),
            .I(\c0.n20449 ));
    LocalMux I__4679 (
            .O(N__34018),
            .I(\c0.n20449 ));
    InMux I__4678 (
            .O(N__34011),
            .I(N__34008));
    LocalMux I__4677 (
            .O(N__34008),
            .I(N__34005));
    Odrv4 I__4676 (
            .O(N__34005),
            .I(\c0.n10_adj_4374 ));
    InMux I__4675 (
            .O(N__34002),
            .I(N__33999));
    LocalMux I__4674 (
            .O(N__33999),
            .I(\c0.data_out_frame_29__7__N_855 ));
    CascadeMux I__4673 (
            .O(N__33996),
            .I(N__33990));
    CascadeMux I__4672 (
            .O(N__33995),
            .I(N__33987));
    CascadeMux I__4671 (
            .O(N__33994),
            .I(N__33984));
    InMux I__4670 (
            .O(N__33993),
            .I(N__33981));
    InMux I__4669 (
            .O(N__33990),
            .I(N__33978));
    InMux I__4668 (
            .O(N__33987),
            .I(N__33973));
    InMux I__4667 (
            .O(N__33984),
            .I(N__33973));
    LocalMux I__4666 (
            .O(N__33981),
            .I(N__33970));
    LocalMux I__4665 (
            .O(N__33978),
            .I(N__33967));
    LocalMux I__4664 (
            .O(N__33973),
            .I(N__33964));
    Span4Mux_h I__4663 (
            .O(N__33970),
            .I(N__33961));
    Odrv4 I__4662 (
            .O(N__33967),
            .I(\c0.n13384 ));
    Odrv4 I__4661 (
            .O(N__33964),
            .I(\c0.n13384 ));
    Odrv4 I__4660 (
            .O(N__33961),
            .I(\c0.n13384 ));
    CascadeMux I__4659 (
            .O(N__33954),
            .I(N__33950));
    InMux I__4658 (
            .O(N__33953),
            .I(N__33947));
    InMux I__4657 (
            .O(N__33950),
            .I(N__33943));
    LocalMux I__4656 (
            .O(N__33947),
            .I(N__33939));
    InMux I__4655 (
            .O(N__33946),
            .I(N__33936));
    LocalMux I__4654 (
            .O(N__33943),
            .I(N__33933));
    InMux I__4653 (
            .O(N__33942),
            .I(N__33930));
    Span4Mux_v I__4652 (
            .O(N__33939),
            .I(N__33925));
    LocalMux I__4651 (
            .O(N__33936),
            .I(N__33925));
    Span4Mux_h I__4650 (
            .O(N__33933),
            .I(N__33922));
    LocalMux I__4649 (
            .O(N__33930),
            .I(encoder1_position_0));
    Odrv4 I__4648 (
            .O(N__33925),
            .I(encoder1_position_0));
    Odrv4 I__4647 (
            .O(N__33922),
            .I(encoder1_position_0));
    InMux I__4646 (
            .O(N__33915),
            .I(N__33912));
    LocalMux I__4645 (
            .O(N__33912),
            .I(N__33908));
    CascadeMux I__4644 (
            .O(N__33911),
            .I(N__33905));
    Span4Mux_v I__4643 (
            .O(N__33908),
            .I(N__33902));
    InMux I__4642 (
            .O(N__33905),
            .I(N__33899));
    Sp12to4 I__4641 (
            .O(N__33902),
            .I(N__33896));
    LocalMux I__4640 (
            .O(N__33899),
            .I(\c0.n22611 ));
    Odrv12 I__4639 (
            .O(N__33896),
            .I(\c0.n22611 ));
    InMux I__4638 (
            .O(N__33891),
            .I(N__33888));
    LocalMux I__4637 (
            .O(N__33888),
            .I(\c0.n10_adj_4274 ));
    CascadeMux I__4636 (
            .O(N__33885),
            .I(N__33881));
    InMux I__4635 (
            .O(N__33884),
            .I(N__33878));
    InMux I__4634 (
            .O(N__33881),
            .I(N__33875));
    LocalMux I__4633 (
            .O(N__33878),
            .I(\c0.n22791 ));
    LocalMux I__4632 (
            .O(N__33875),
            .I(\c0.n22791 ));
    InMux I__4631 (
            .O(N__33870),
            .I(N__33866));
    InMux I__4630 (
            .O(N__33869),
            .I(N__33863));
    LocalMux I__4629 (
            .O(N__33866),
            .I(N__33860));
    LocalMux I__4628 (
            .O(N__33863),
            .I(\c0.n22466 ));
    Odrv4 I__4627 (
            .O(N__33860),
            .I(\c0.n22466 ));
    InMux I__4626 (
            .O(N__33855),
            .I(N__33847));
    InMux I__4625 (
            .O(N__33854),
            .I(N__33847));
    InMux I__4624 (
            .O(N__33853),
            .I(N__33844));
    InMux I__4623 (
            .O(N__33852),
            .I(N__33841));
    LocalMux I__4622 (
            .O(N__33847),
            .I(N__33838));
    LocalMux I__4621 (
            .O(N__33844),
            .I(N__33835));
    LocalMux I__4620 (
            .O(N__33841),
            .I(\c0.n13121 ));
    Odrv4 I__4619 (
            .O(N__33838),
            .I(\c0.n13121 ));
    Odrv4 I__4618 (
            .O(N__33835),
            .I(\c0.n13121 ));
    InMux I__4617 (
            .O(N__33828),
            .I(N__33825));
    LocalMux I__4616 (
            .O(N__33825),
            .I(N__33822));
    Odrv4 I__4615 (
            .O(N__33822),
            .I(\c0.n34_adj_4328 ));
    CascadeMux I__4614 (
            .O(N__33819),
            .I(\c0.n30_adj_4326_cascade_ ));
    InMux I__4613 (
            .O(N__33816),
            .I(N__33813));
    LocalMux I__4612 (
            .O(N__33813),
            .I(\c0.n29_adj_4329 ));
    CascadeMux I__4611 (
            .O(N__33810),
            .I(N__33807));
    InMux I__4610 (
            .O(N__33807),
            .I(N__33803));
    CascadeMux I__4609 (
            .O(N__33806),
            .I(N__33800));
    LocalMux I__4608 (
            .O(N__33803),
            .I(N__33795));
    InMux I__4607 (
            .O(N__33800),
            .I(N__33792));
    InMux I__4606 (
            .O(N__33799),
            .I(N__33789));
    InMux I__4605 (
            .O(N__33798),
            .I(N__33786));
    Span12Mux_v I__4604 (
            .O(N__33795),
            .I(N__33781));
    LocalMux I__4603 (
            .O(N__33792),
            .I(N__33781));
    LocalMux I__4602 (
            .O(N__33789),
            .I(N__33778));
    LocalMux I__4601 (
            .O(N__33786),
            .I(encoder1_position_20));
    Odrv12 I__4600 (
            .O(N__33781),
            .I(encoder1_position_20));
    Odrv4 I__4599 (
            .O(N__33778),
            .I(encoder1_position_20));
    CascadeMux I__4598 (
            .O(N__33771),
            .I(N__33768));
    InMux I__4597 (
            .O(N__33768),
            .I(N__33765));
    LocalMux I__4596 (
            .O(N__33765),
            .I(\c0.n22788 ));
    CascadeMux I__4595 (
            .O(N__33762),
            .I(\c0.n22788_cascade_ ));
    SRMux I__4594 (
            .O(N__33759),
            .I(N__33756));
    LocalMux I__4593 (
            .O(N__33756),
            .I(N__33753));
    Span4Mux_h I__4592 (
            .O(N__33753),
            .I(N__33750));
    Odrv4 I__4591 (
            .O(N__33750),
            .I(\c0.n21637 ));
    InMux I__4590 (
            .O(N__33747),
            .I(N__33744));
    LocalMux I__4589 (
            .O(N__33744),
            .I(\c0.n22638 ));
    CascadeMux I__4588 (
            .O(N__33741),
            .I(\c0.n22831_cascade_ ));
    InMux I__4587 (
            .O(N__33738),
            .I(N__33735));
    LocalMux I__4586 (
            .O(N__33735),
            .I(N__33732));
    Odrv4 I__4585 (
            .O(N__33732),
            .I(\c0.n20_adj_4321 ));
    CascadeMux I__4584 (
            .O(N__33729),
            .I(\c0.n13_adj_4320_cascade_ ));
    InMux I__4583 (
            .O(N__33726),
            .I(N__33723));
    LocalMux I__4582 (
            .O(N__33723),
            .I(\c0.n14_adj_4319 ));
    CascadeMux I__4581 (
            .O(N__33720),
            .I(\c0.n28_adj_4322_cascade_ ));
    InMux I__4580 (
            .O(N__33717),
            .I(N__33712));
    InMux I__4579 (
            .O(N__33716),
            .I(N__33707));
    InMux I__4578 (
            .O(N__33715),
            .I(N__33707));
    LocalMux I__4577 (
            .O(N__33712),
            .I(\c0.n12488 ));
    LocalMux I__4576 (
            .O(N__33707),
            .I(\c0.n12488 ));
    InMux I__4575 (
            .O(N__33702),
            .I(N__33697));
    CascadeMux I__4574 (
            .O(N__33701),
            .I(N__33694));
    CascadeMux I__4573 (
            .O(N__33700),
            .I(N__33690));
    LocalMux I__4572 (
            .O(N__33697),
            .I(N__33687));
    InMux I__4571 (
            .O(N__33694),
            .I(N__33683));
    InMux I__4570 (
            .O(N__33693),
            .I(N__33678));
    InMux I__4569 (
            .O(N__33690),
            .I(N__33678));
    Span4Mux_v I__4568 (
            .O(N__33687),
            .I(N__33675));
    InMux I__4567 (
            .O(N__33686),
            .I(N__33672));
    LocalMux I__4566 (
            .O(N__33683),
            .I(N__33668));
    LocalMux I__4565 (
            .O(N__33678),
            .I(N__33665));
    Span4Mux_v I__4564 (
            .O(N__33675),
            .I(N__33662));
    LocalMux I__4563 (
            .O(N__33672),
            .I(N__33659));
    InMux I__4562 (
            .O(N__33671),
            .I(N__33656));
    Span4Mux_v I__4561 (
            .O(N__33668),
            .I(N__33653));
    Span4Mux_h I__4560 (
            .O(N__33665),
            .I(N__33650));
    Span4Mux_v I__4559 (
            .O(N__33662),
            .I(N__33645));
    Span4Mux_v I__4558 (
            .O(N__33659),
            .I(N__33645));
    LocalMux I__4557 (
            .O(N__33656),
            .I(encoder1_position_14));
    Odrv4 I__4556 (
            .O(N__33653),
            .I(encoder1_position_14));
    Odrv4 I__4555 (
            .O(N__33650),
            .I(encoder1_position_14));
    Odrv4 I__4554 (
            .O(N__33645),
            .I(encoder1_position_14));
    CascadeMux I__4553 (
            .O(N__33636),
            .I(\c0.n20318_cascade_ ));
    SRMux I__4552 (
            .O(N__33633),
            .I(N__33630));
    LocalMux I__4551 (
            .O(N__33630),
            .I(N__33627));
    Span4Mux_h I__4550 (
            .O(N__33627),
            .I(N__33624));
    Odrv4 I__4549 (
            .O(N__33624),
            .I(\c0.n21579 ));
    InMux I__4548 (
            .O(N__33621),
            .I(N__33615));
    InMux I__4547 (
            .O(N__33620),
            .I(N__33615));
    LocalMux I__4546 (
            .O(N__33615),
            .I(\c0.n4_adj_4678 ));
    InMux I__4545 (
            .O(N__33612),
            .I(N__33607));
    CascadeMux I__4544 (
            .O(N__33611),
            .I(N__33604));
    CascadeMux I__4543 (
            .O(N__33610),
            .I(N__33601));
    LocalMux I__4542 (
            .O(N__33607),
            .I(N__33597));
    InMux I__4541 (
            .O(N__33604),
            .I(N__33594));
    InMux I__4540 (
            .O(N__33601),
            .I(N__33589));
    InMux I__4539 (
            .O(N__33600),
            .I(N__33586));
    Span4Mux_h I__4538 (
            .O(N__33597),
            .I(N__33581));
    LocalMux I__4537 (
            .O(N__33594),
            .I(N__33581));
    InMux I__4536 (
            .O(N__33593),
            .I(N__33578));
    InMux I__4535 (
            .O(N__33592),
            .I(N__33575));
    LocalMux I__4534 (
            .O(N__33589),
            .I(N__33572));
    LocalMux I__4533 (
            .O(N__33586),
            .I(N__33569));
    Span4Mux_v I__4532 (
            .O(N__33581),
            .I(N__33566));
    LocalMux I__4531 (
            .O(N__33578),
            .I(N__33563));
    LocalMux I__4530 (
            .O(N__33575),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv12 I__4529 (
            .O(N__33572),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv12 I__4528 (
            .O(N__33569),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv4 I__4527 (
            .O(N__33566),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv4 I__4526 (
            .O(N__33563),
            .I(\c0.FRAME_MATCHER_state_28 ));
    InMux I__4525 (
            .O(N__33552),
            .I(N__33548));
    InMux I__4524 (
            .O(N__33551),
            .I(N__33545));
    LocalMux I__4523 (
            .O(N__33548),
            .I(N__33538));
    LocalMux I__4522 (
            .O(N__33545),
            .I(N__33538));
    InMux I__4521 (
            .O(N__33544),
            .I(N__33535));
    InMux I__4520 (
            .O(N__33543),
            .I(N__33532));
    Odrv4 I__4519 (
            .O(N__33538),
            .I(\c0.n22131 ));
    LocalMux I__4518 (
            .O(N__33535),
            .I(\c0.n22131 ));
    LocalMux I__4517 (
            .O(N__33532),
            .I(\c0.n22131 ));
    CascadeMux I__4516 (
            .O(N__33525),
            .I(N__33520));
    InMux I__4515 (
            .O(N__33524),
            .I(N__33517));
    InMux I__4514 (
            .O(N__33523),
            .I(N__33514));
    InMux I__4513 (
            .O(N__33520),
            .I(N__33511));
    LocalMux I__4512 (
            .O(N__33517),
            .I(N__33508));
    LocalMux I__4511 (
            .O(N__33514),
            .I(\c0.FRAME_MATCHER_state_9 ));
    LocalMux I__4510 (
            .O(N__33511),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__4509 (
            .O(N__33508),
            .I(\c0.FRAME_MATCHER_state_9 ));
    InMux I__4508 (
            .O(N__33501),
            .I(N__33496));
    InMux I__4507 (
            .O(N__33500),
            .I(N__33491));
    InMux I__4506 (
            .O(N__33499),
            .I(N__33491));
    LocalMux I__4505 (
            .O(N__33496),
            .I(\c0.FRAME_MATCHER_state_5 ));
    LocalMux I__4504 (
            .O(N__33491),
            .I(\c0.FRAME_MATCHER_state_5 ));
    SRMux I__4503 (
            .O(N__33486),
            .I(N__33483));
    LocalMux I__4502 (
            .O(N__33483),
            .I(\c0.n21625 ));
    SRMux I__4501 (
            .O(N__33480),
            .I(N__33477));
    LocalMux I__4500 (
            .O(N__33477),
            .I(N__33474));
    Odrv4 I__4499 (
            .O(N__33474),
            .I(\c0.n8_adj_4561 ));
    InMux I__4498 (
            .O(N__33471),
            .I(N__33467));
    InMux I__4497 (
            .O(N__33470),
            .I(N__33463));
    LocalMux I__4496 (
            .O(N__33467),
            .I(N__33460));
    InMux I__4495 (
            .O(N__33466),
            .I(N__33457));
    LocalMux I__4494 (
            .O(N__33463),
            .I(N__33454));
    Span4Mux_h I__4493 (
            .O(N__33460),
            .I(N__33451));
    LocalMux I__4492 (
            .O(N__33457),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv12 I__4491 (
            .O(N__33454),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__4490 (
            .O(N__33451),
            .I(\c0.FRAME_MATCHER_state_8 ));
    SRMux I__4489 (
            .O(N__33444),
            .I(N__33441));
    LocalMux I__4488 (
            .O(N__33441),
            .I(N__33438));
    Odrv12 I__4487 (
            .O(N__33438),
            .I(\c0.n8_adj_4558 ));
    CascadeMux I__4486 (
            .O(N__33435),
            .I(\c0.data_out_frame_29_7_N_1482_0_cascade_ ));
    InMux I__4485 (
            .O(N__33432),
            .I(N__33429));
    LocalMux I__4484 (
            .O(N__33429),
            .I(\c0.n6_adj_4495 ));
    InMux I__4483 (
            .O(N__33426),
            .I(N__33423));
    LocalMux I__4482 (
            .O(N__33423),
            .I(\c0.n14784 ));
    CascadeMux I__4481 (
            .O(N__33420),
            .I(\c0.n9706_cascade_ ));
    CascadeMux I__4480 (
            .O(N__33417),
            .I(\c0.n6_cascade_ ));
    InMux I__4479 (
            .O(N__33414),
            .I(N__33410));
    InMux I__4478 (
            .O(N__33413),
            .I(N__33407));
    LocalMux I__4477 (
            .O(N__33410),
            .I(N__33402));
    LocalMux I__4476 (
            .O(N__33407),
            .I(N__33402));
    Odrv4 I__4475 (
            .O(N__33402),
            .I(data_out_frame_9_6));
    InMux I__4474 (
            .O(N__33399),
            .I(N__33395));
    InMux I__4473 (
            .O(N__33398),
            .I(N__33392));
    LocalMux I__4472 (
            .O(N__33395),
            .I(data_out_frame_6_6));
    LocalMux I__4471 (
            .O(N__33392),
            .I(data_out_frame_6_6));
    InMux I__4470 (
            .O(N__33387),
            .I(N__33384));
    LocalMux I__4469 (
            .O(N__33384),
            .I(N__33381));
    Span4Mux_h I__4468 (
            .O(N__33381),
            .I(N__33377));
    InMux I__4467 (
            .O(N__33380),
            .I(N__33374));
    Odrv4 I__4466 (
            .O(N__33377),
            .I(n14247));
    LocalMux I__4465 (
            .O(N__33374),
            .I(n14247));
    CascadeMux I__4464 (
            .O(N__33369),
            .I(N__33366));
    InMux I__4463 (
            .O(N__33366),
            .I(N__33363));
    LocalMux I__4462 (
            .O(N__33363),
            .I(N__33359));
    CascadeMux I__4461 (
            .O(N__33362),
            .I(N__33356));
    Span4Mux_v I__4460 (
            .O(N__33359),
            .I(N__33353));
    InMux I__4459 (
            .O(N__33356),
            .I(N__33350));
    Span4Mux_v I__4458 (
            .O(N__33353),
            .I(N__33347));
    LocalMux I__4457 (
            .O(N__33350),
            .I(data_out_frame_0_4));
    Odrv4 I__4456 (
            .O(N__33347),
            .I(data_out_frame_0_4));
    InMux I__4455 (
            .O(N__33342),
            .I(N__33338));
    InMux I__4454 (
            .O(N__33341),
            .I(N__33335));
    LocalMux I__4453 (
            .O(N__33338),
            .I(N__33332));
    LocalMux I__4452 (
            .O(N__33335),
            .I(data_out_frame_9_2));
    Odrv4 I__4451 (
            .O(N__33332),
            .I(data_out_frame_9_2));
    InMux I__4450 (
            .O(N__33327),
            .I(N__33323));
    InMux I__4449 (
            .O(N__33326),
            .I(N__33320));
    LocalMux I__4448 (
            .O(N__33323),
            .I(data_out_frame_11_4));
    LocalMux I__4447 (
            .O(N__33320),
            .I(data_out_frame_11_4));
    InMux I__4446 (
            .O(N__33315),
            .I(N__33312));
    LocalMux I__4445 (
            .O(N__33312),
            .I(N__33308));
    CascadeMux I__4444 (
            .O(N__33311),
            .I(N__33305));
    Span4Mux_v I__4443 (
            .O(N__33308),
            .I(N__33302));
    InMux I__4442 (
            .O(N__33305),
            .I(N__33299));
    Span4Mux_v I__4441 (
            .O(N__33302),
            .I(N__33296));
    LocalMux I__4440 (
            .O(N__33299),
            .I(data_out_frame_13_2));
    Odrv4 I__4439 (
            .O(N__33296),
            .I(data_out_frame_13_2));
    InMux I__4438 (
            .O(N__33291),
            .I(N__33288));
    LocalMux I__4437 (
            .O(N__33288),
            .I(\c0.n12976 ));
    CascadeMux I__4436 (
            .O(N__33285),
            .I(\c0.n12976_cascade_ ));
    InMux I__4435 (
            .O(N__33282),
            .I(N__33279));
    LocalMux I__4434 (
            .O(N__33279),
            .I(N__33276));
    Span4Mux_h I__4433 (
            .O(N__33276),
            .I(N__33273));
    Odrv4 I__4432 (
            .O(N__33273),
            .I(n2275));
    InMux I__4431 (
            .O(N__33270),
            .I(N__33266));
    InMux I__4430 (
            .O(N__33269),
            .I(N__33263));
    LocalMux I__4429 (
            .O(N__33266),
            .I(data_out_frame_10_0));
    LocalMux I__4428 (
            .O(N__33263),
            .I(data_out_frame_10_0));
    InMux I__4427 (
            .O(N__33258),
            .I(N__33255));
    LocalMux I__4426 (
            .O(N__33255),
            .I(N__33251));
    InMux I__4425 (
            .O(N__33254),
            .I(N__33248));
    Span4Mux_h I__4424 (
            .O(N__33251),
            .I(N__33245));
    LocalMux I__4423 (
            .O(N__33248),
            .I(data_out_frame_10_4));
    Odrv4 I__4422 (
            .O(N__33245),
            .I(data_out_frame_10_4));
    InMux I__4421 (
            .O(N__33240),
            .I(N__33237));
    LocalMux I__4420 (
            .O(N__33237),
            .I(\c0.n24783 ));
    InMux I__4419 (
            .O(N__33234),
            .I(N__33230));
    InMux I__4418 (
            .O(N__33233),
            .I(N__33227));
    LocalMux I__4417 (
            .O(N__33230),
            .I(N__33224));
    LocalMux I__4416 (
            .O(N__33227),
            .I(data_out_frame_6_0));
    Odrv12 I__4415 (
            .O(N__33224),
            .I(data_out_frame_6_0));
    CascadeMux I__4414 (
            .O(N__33219),
            .I(N__33216));
    InMux I__4413 (
            .O(N__33216),
            .I(N__33212));
    CascadeMux I__4412 (
            .O(N__33215),
            .I(N__33209));
    LocalMux I__4411 (
            .O(N__33212),
            .I(N__33206));
    InMux I__4410 (
            .O(N__33209),
            .I(N__33203));
    Odrv12 I__4409 (
            .O(N__33206),
            .I(\c0.tx_transmit_N_3650 ));
    LocalMux I__4408 (
            .O(N__33203),
            .I(\c0.tx_transmit_N_3650 ));
    InMux I__4407 (
            .O(N__33198),
            .I(N__33195));
    LocalMux I__4406 (
            .O(N__33195),
            .I(N__33192));
    Span4Mux_v I__4405 (
            .O(N__33192),
            .I(N__33189));
    Odrv4 I__4404 (
            .O(N__33189),
            .I(\c0.n24888 ));
    InMux I__4403 (
            .O(N__33186),
            .I(N__33182));
    InMux I__4402 (
            .O(N__33185),
            .I(N__33179));
    LocalMux I__4401 (
            .O(N__33182),
            .I(N__33174));
    LocalMux I__4400 (
            .O(N__33179),
            .I(N__33174));
    Odrv4 I__4399 (
            .O(N__33174),
            .I(data_out_frame_12_0));
    InMux I__4398 (
            .O(N__33171),
            .I(N__33168));
    LocalMux I__4397 (
            .O(N__33168),
            .I(N__33165));
    Span4Mux_v I__4396 (
            .O(N__33165),
            .I(N__33161));
    InMux I__4395 (
            .O(N__33164),
            .I(N__33158));
    Span4Mux_h I__4394 (
            .O(N__33161),
            .I(N__33155));
    LocalMux I__4393 (
            .O(N__33158),
            .I(data_out_frame_12_1));
    Odrv4 I__4392 (
            .O(N__33155),
            .I(data_out_frame_12_1));
    InMux I__4391 (
            .O(N__33150),
            .I(\quad_counter1.n19759 ));
    InMux I__4390 (
            .O(N__33147),
            .I(\quad_counter1.n19760 ));
    InMux I__4389 (
            .O(N__33144),
            .I(\quad_counter1.n19761 ));
    InMux I__4388 (
            .O(N__33141),
            .I(N__33126));
    CascadeMux I__4387 (
            .O(N__33140),
            .I(N__33122));
    CascadeMux I__4386 (
            .O(N__33139),
            .I(N__33118));
    CascadeMux I__4385 (
            .O(N__33138),
            .I(N__33114));
    CascadeMux I__4384 (
            .O(N__33137),
            .I(N__33110));
    CascadeMux I__4383 (
            .O(N__33136),
            .I(N__33106));
    CascadeMux I__4382 (
            .O(N__33135),
            .I(N__33102));
    CascadeMux I__4381 (
            .O(N__33134),
            .I(N__33098));
    CascadeMux I__4380 (
            .O(N__33133),
            .I(N__33094));
    CascadeMux I__4379 (
            .O(N__33132),
            .I(N__33090));
    CascadeMux I__4378 (
            .O(N__33131),
            .I(N__33086));
    CascadeMux I__4377 (
            .O(N__33130),
            .I(N__33082));
    CascadeMux I__4376 (
            .O(N__33129),
            .I(N__33078));
    LocalMux I__4375 (
            .O(N__33126),
            .I(N__33068));
    InMux I__4374 (
            .O(N__33125),
            .I(N__33051));
    InMux I__4373 (
            .O(N__33122),
            .I(N__33051));
    InMux I__4372 (
            .O(N__33121),
            .I(N__33051));
    InMux I__4371 (
            .O(N__33118),
            .I(N__33051));
    InMux I__4370 (
            .O(N__33117),
            .I(N__33051));
    InMux I__4369 (
            .O(N__33114),
            .I(N__33051));
    InMux I__4368 (
            .O(N__33113),
            .I(N__33051));
    InMux I__4367 (
            .O(N__33110),
            .I(N__33051));
    InMux I__4366 (
            .O(N__33109),
            .I(N__33034));
    InMux I__4365 (
            .O(N__33106),
            .I(N__33034));
    InMux I__4364 (
            .O(N__33105),
            .I(N__33034));
    InMux I__4363 (
            .O(N__33102),
            .I(N__33034));
    InMux I__4362 (
            .O(N__33101),
            .I(N__33034));
    InMux I__4361 (
            .O(N__33098),
            .I(N__33034));
    InMux I__4360 (
            .O(N__33097),
            .I(N__33034));
    InMux I__4359 (
            .O(N__33094),
            .I(N__33034));
    InMux I__4358 (
            .O(N__33093),
            .I(N__33017));
    InMux I__4357 (
            .O(N__33090),
            .I(N__33017));
    InMux I__4356 (
            .O(N__33089),
            .I(N__33017));
    InMux I__4355 (
            .O(N__33086),
            .I(N__33017));
    InMux I__4354 (
            .O(N__33085),
            .I(N__33017));
    InMux I__4353 (
            .O(N__33082),
            .I(N__33017));
    InMux I__4352 (
            .O(N__33081),
            .I(N__33017));
    InMux I__4351 (
            .O(N__33078),
            .I(N__33017));
    CascadeMux I__4350 (
            .O(N__33077),
            .I(N__33014));
    CascadeMux I__4349 (
            .O(N__33076),
            .I(N__33011));
    CascadeMux I__4348 (
            .O(N__33075),
            .I(N__33008));
    CascadeMux I__4347 (
            .O(N__33074),
            .I(N__33005));
    CascadeMux I__4346 (
            .O(N__33073),
            .I(N__33002));
    CascadeMux I__4345 (
            .O(N__33072),
            .I(N__32999));
    CascadeMux I__4344 (
            .O(N__33071),
            .I(N__32996));
    Span4Mux_v I__4343 (
            .O(N__33068),
            .I(N__32990));
    LocalMux I__4342 (
            .O(N__33051),
            .I(N__32990));
    LocalMux I__4341 (
            .O(N__33034),
            .I(N__32987));
    LocalMux I__4340 (
            .O(N__33017),
            .I(N__32984));
    InMux I__4339 (
            .O(N__33014),
            .I(N__32975));
    InMux I__4338 (
            .O(N__33011),
            .I(N__32975));
    InMux I__4337 (
            .O(N__33008),
            .I(N__32975));
    InMux I__4336 (
            .O(N__33005),
            .I(N__32975));
    InMux I__4335 (
            .O(N__33002),
            .I(N__32966));
    InMux I__4334 (
            .O(N__32999),
            .I(N__32966));
    InMux I__4333 (
            .O(N__32996),
            .I(N__32966));
    InMux I__4332 (
            .O(N__32995),
            .I(N__32966));
    Span4Mux_v I__4331 (
            .O(N__32990),
            .I(N__32963));
    Span4Mux_h I__4330 (
            .O(N__32987),
            .I(N__32960));
    Span4Mux_h I__4329 (
            .O(N__32984),
            .I(N__32957));
    LocalMux I__4328 (
            .O(N__32975),
            .I(N__32952));
    LocalMux I__4327 (
            .O(N__32966),
            .I(N__32952));
    Span4Mux_v I__4326 (
            .O(N__32963),
            .I(N__32949));
    Span4Mux_v I__4325 (
            .O(N__32960),
            .I(N__32946));
    Sp12to4 I__4324 (
            .O(N__32957),
            .I(N__32941));
    Span12Mux_h I__4323 (
            .O(N__32952),
            .I(N__32941));
    Odrv4 I__4322 (
            .O(N__32949),
            .I(\quad_counter1.n2226 ));
    Odrv4 I__4321 (
            .O(N__32946),
            .I(\quad_counter1.n2226 ));
    Odrv12 I__4320 (
            .O(N__32941),
            .I(\quad_counter1.n2226 ));
    InMux I__4319 (
            .O(N__32934),
            .I(bfn_12_19_0_));
    CascadeMux I__4318 (
            .O(N__32931),
            .I(\c0.n24784_cascade_ ));
    InMux I__4317 (
            .O(N__32928),
            .I(N__32925));
    LocalMux I__4316 (
            .O(N__32925),
            .I(N__32922));
    Span4Mux_v I__4315 (
            .O(N__32922),
            .I(N__32919));
    Span4Mux_v I__4314 (
            .O(N__32919),
            .I(N__32916));
    Odrv4 I__4313 (
            .O(N__32916),
            .I(n25019));
    CascadeMux I__4312 (
            .O(N__32913),
            .I(N__32909));
    InMux I__4311 (
            .O(N__32912),
            .I(N__32906));
    InMux I__4310 (
            .O(N__32909),
            .I(N__32903));
    LocalMux I__4309 (
            .O(N__32906),
            .I(data_out_frame_11_2));
    LocalMux I__4308 (
            .O(N__32903),
            .I(data_out_frame_11_2));
    InMux I__4307 (
            .O(N__32898),
            .I(N__32895));
    LocalMux I__4306 (
            .O(N__32895),
            .I(N__32892));
    Odrv4 I__4305 (
            .O(N__32892),
            .I(n2273));
    CascadeMux I__4304 (
            .O(N__32889),
            .I(N__32885));
    CascadeMux I__4303 (
            .O(N__32888),
            .I(N__32881));
    InMux I__4302 (
            .O(N__32885),
            .I(N__32878));
    CascadeMux I__4301 (
            .O(N__32884),
            .I(N__32874));
    InMux I__4300 (
            .O(N__32881),
            .I(N__32871));
    LocalMux I__4299 (
            .O(N__32878),
            .I(N__32868));
    InMux I__4298 (
            .O(N__32877),
            .I(N__32863));
    InMux I__4297 (
            .O(N__32874),
            .I(N__32863));
    LocalMux I__4296 (
            .O(N__32871),
            .I(N__32858));
    Span4Mux_v I__4295 (
            .O(N__32868),
            .I(N__32858));
    LocalMux I__4294 (
            .O(N__32863),
            .I(encoder1_position_18));
    Odrv4 I__4293 (
            .O(N__32858),
            .I(encoder1_position_18));
    InMux I__4292 (
            .O(N__32853),
            .I(N__32850));
    LocalMux I__4291 (
            .O(N__32850),
            .I(N__32844));
    InMux I__4290 (
            .O(N__32849),
            .I(N__32841));
    InMux I__4289 (
            .O(N__32848),
            .I(N__32838));
    InMux I__4288 (
            .O(N__32847),
            .I(N__32835));
    Sp12to4 I__4287 (
            .O(N__32844),
            .I(N__32830));
    LocalMux I__4286 (
            .O(N__32841),
            .I(N__32830));
    LocalMux I__4285 (
            .O(N__32838),
            .I(N__32827));
    LocalMux I__4284 (
            .O(N__32835),
            .I(encoder1_position_19));
    Odrv12 I__4283 (
            .O(N__32830),
            .I(encoder1_position_19));
    Odrv4 I__4282 (
            .O(N__32827),
            .I(encoder1_position_19));
    InMux I__4281 (
            .O(N__32820),
            .I(N__32817));
    LocalMux I__4280 (
            .O(N__32817),
            .I(N__32814));
    Span4Mux_v I__4279 (
            .O(N__32814),
            .I(N__32811));
    Odrv4 I__4278 (
            .O(N__32811),
            .I(n2272));
    InMux I__4277 (
            .O(N__32808),
            .I(\quad_counter1.n19750 ));
    InMux I__4276 (
            .O(N__32805),
            .I(N__32802));
    LocalMux I__4275 (
            .O(N__32802),
            .I(N__32799));
    Odrv12 I__4274 (
            .O(N__32799),
            .I(n2271));
    InMux I__4273 (
            .O(N__32796),
            .I(\quad_counter1.n19751 ));
    InMux I__4272 (
            .O(N__32793),
            .I(\quad_counter1.n19752 ));
    InMux I__4271 (
            .O(N__32790),
            .I(N__32787));
    LocalMux I__4270 (
            .O(N__32787),
            .I(N__32784));
    Span4Mux_h I__4269 (
            .O(N__32784),
            .I(N__32781));
    Odrv4 I__4268 (
            .O(N__32781),
            .I(n2269));
    InMux I__4267 (
            .O(N__32778),
            .I(\quad_counter1.n19753 ));
    InMux I__4266 (
            .O(N__32775),
            .I(bfn_12_18_0_));
    InMux I__4265 (
            .O(N__32772),
            .I(\quad_counter1.n19755 ));
    InMux I__4264 (
            .O(N__32769),
            .I(N__32766));
    LocalMux I__4263 (
            .O(N__32766),
            .I(N__32763));
    Span4Mux_h I__4262 (
            .O(N__32763),
            .I(N__32760));
    Span4Mux_v I__4261 (
            .O(N__32760),
            .I(N__32757));
    Odrv4 I__4260 (
            .O(N__32757),
            .I(n2266));
    InMux I__4259 (
            .O(N__32754),
            .I(\quad_counter1.n19756 ));
    InMux I__4258 (
            .O(N__32751),
            .I(\quad_counter1.n19757 ));
    InMux I__4257 (
            .O(N__32748),
            .I(\quad_counter1.n19758 ));
    InMux I__4256 (
            .O(N__32745),
            .I(N__32742));
    LocalMux I__4255 (
            .O(N__32742),
            .I(N__32739));
    Span4Mux_v I__4254 (
            .O(N__32739),
            .I(N__32736));
    Odrv4 I__4253 (
            .O(N__32736),
            .I(n2280));
    InMux I__4252 (
            .O(N__32733),
            .I(\quad_counter1.n19742 ));
    InMux I__4251 (
            .O(N__32730),
            .I(N__32727));
    LocalMux I__4250 (
            .O(N__32727),
            .I(N__32724));
    Span4Mux_v I__4249 (
            .O(N__32724),
            .I(N__32721));
    Odrv4 I__4248 (
            .O(N__32721),
            .I(n2279));
    InMux I__4247 (
            .O(N__32718),
            .I(\quad_counter1.n19743 ));
    CascadeMux I__4246 (
            .O(N__32715),
            .I(N__32712));
    InMux I__4245 (
            .O(N__32712),
            .I(N__32708));
    InMux I__4244 (
            .O(N__32711),
            .I(N__32703));
    LocalMux I__4243 (
            .O(N__32708),
            .I(N__32700));
    InMux I__4242 (
            .O(N__32707),
            .I(N__32695));
    InMux I__4241 (
            .O(N__32706),
            .I(N__32695));
    LocalMux I__4240 (
            .O(N__32703),
            .I(N__32691));
    Span4Mux_v I__4239 (
            .O(N__32700),
            .I(N__32688));
    LocalMux I__4238 (
            .O(N__32695),
            .I(N__32685));
    InMux I__4237 (
            .O(N__32694),
            .I(N__32681));
    Span12Mux_h I__4236 (
            .O(N__32691),
            .I(N__32678));
    Span4Mux_v I__4235 (
            .O(N__32688),
            .I(N__32673));
    Span4Mux_h I__4234 (
            .O(N__32685),
            .I(N__32673));
    InMux I__4233 (
            .O(N__32684),
            .I(N__32670));
    LocalMux I__4232 (
            .O(N__32681),
            .I(encoder1_position_13));
    Odrv12 I__4231 (
            .O(N__32678),
            .I(encoder1_position_13));
    Odrv4 I__4230 (
            .O(N__32673),
            .I(encoder1_position_13));
    LocalMux I__4229 (
            .O(N__32670),
            .I(encoder1_position_13));
    InMux I__4228 (
            .O(N__32661),
            .I(N__32658));
    LocalMux I__4227 (
            .O(N__32658),
            .I(N__32655));
    Span4Mux_v I__4226 (
            .O(N__32655),
            .I(N__32652));
    Span4Mux_v I__4225 (
            .O(N__32652),
            .I(N__32649));
    Odrv4 I__4224 (
            .O(N__32649),
            .I(n2278));
    InMux I__4223 (
            .O(N__32646),
            .I(\quad_counter1.n19744 ));
    InMux I__4222 (
            .O(N__32643),
            .I(N__32640));
    LocalMux I__4221 (
            .O(N__32640),
            .I(N__32637));
    Span4Mux_h I__4220 (
            .O(N__32637),
            .I(N__32634));
    Span4Mux_v I__4219 (
            .O(N__32634),
            .I(N__32631));
    Odrv4 I__4218 (
            .O(N__32631),
            .I(n2277));
    InMux I__4217 (
            .O(N__32628),
            .I(\quad_counter1.n19745 ));
    InMux I__4216 (
            .O(N__32625),
            .I(N__32622));
    LocalMux I__4215 (
            .O(N__32622),
            .I(n2276));
    InMux I__4214 (
            .O(N__32619),
            .I(bfn_12_17_0_));
    InMux I__4213 (
            .O(N__32616),
            .I(\quad_counter1.n19747 ));
    InMux I__4212 (
            .O(N__32613),
            .I(\quad_counter1.n19748 ));
    InMux I__4211 (
            .O(N__32610),
            .I(\quad_counter1.n19749 ));
    InMux I__4210 (
            .O(N__32607),
            .I(N__32604));
    LocalMux I__4209 (
            .O(N__32604),
            .I(N__32601));
    Odrv4 I__4208 (
            .O(N__32601),
            .I(n2289));
    InMux I__4207 (
            .O(N__32598),
            .I(\quad_counter1.n19733 ));
    InMux I__4206 (
            .O(N__32595),
            .I(N__32592));
    LocalMux I__4205 (
            .O(N__32592),
            .I(N__32589));
    Sp12to4 I__4204 (
            .O(N__32589),
            .I(N__32586));
    Odrv12 I__4203 (
            .O(N__32586),
            .I(n2288));
    InMux I__4202 (
            .O(N__32583),
            .I(\quad_counter1.n19734 ));
    InMux I__4201 (
            .O(N__32580),
            .I(N__32577));
    LocalMux I__4200 (
            .O(N__32577),
            .I(N__32574));
    Odrv12 I__4199 (
            .O(N__32574),
            .I(n2287));
    InMux I__4198 (
            .O(N__32571),
            .I(\quad_counter1.n19735 ));
    InMux I__4197 (
            .O(N__32568),
            .I(N__32565));
    LocalMux I__4196 (
            .O(N__32565),
            .I(N__32562));
    Span4Mux_h I__4195 (
            .O(N__32562),
            .I(N__32559));
    Span4Mux_v I__4194 (
            .O(N__32559),
            .I(N__32556));
    Odrv4 I__4193 (
            .O(N__32556),
            .I(n2286));
    InMux I__4192 (
            .O(N__32553),
            .I(\quad_counter1.n19736 ));
    InMux I__4191 (
            .O(N__32550),
            .I(N__32547));
    LocalMux I__4190 (
            .O(N__32547),
            .I(N__32544));
    Span4Mux_h I__4189 (
            .O(N__32544),
            .I(N__32541));
    Odrv4 I__4188 (
            .O(N__32541),
            .I(n2285));
    InMux I__4187 (
            .O(N__32538),
            .I(\quad_counter1.n19737 ));
    InMux I__4186 (
            .O(N__32535),
            .I(N__32532));
    LocalMux I__4185 (
            .O(N__32532),
            .I(n2284));
    InMux I__4184 (
            .O(N__32529),
            .I(bfn_12_16_0_));
    InMux I__4183 (
            .O(N__32526),
            .I(\quad_counter1.n19739 ));
    InMux I__4182 (
            .O(N__32523),
            .I(N__32520));
    LocalMux I__4181 (
            .O(N__32520),
            .I(N__32517));
    Span4Mux_h I__4180 (
            .O(N__32517),
            .I(N__32514));
    Span4Mux_v I__4179 (
            .O(N__32514),
            .I(N__32511));
    Odrv4 I__4178 (
            .O(N__32511),
            .I(n2282));
    InMux I__4177 (
            .O(N__32508),
            .I(\quad_counter1.n19740 ));
    InMux I__4176 (
            .O(N__32505),
            .I(\quad_counter1.n19741 ));
    CascadeMux I__4175 (
            .O(N__32502),
            .I(N__32499));
    InMux I__4174 (
            .O(N__32499),
            .I(N__32495));
    InMux I__4173 (
            .O(N__32498),
            .I(N__32492));
    LocalMux I__4172 (
            .O(N__32495),
            .I(data_out_frame_7_0));
    LocalMux I__4171 (
            .O(N__32492),
            .I(data_out_frame_7_0));
    InMux I__4170 (
            .O(N__32487),
            .I(N__32484));
    LocalMux I__4169 (
            .O(N__32484),
            .I(N__32481));
    Span4Mux_v I__4168 (
            .O(N__32481),
            .I(N__32478));
    Odrv4 I__4167 (
            .O(N__32478),
            .I(\c0.n5_adj_4567 ));
    InMux I__4166 (
            .O(N__32475),
            .I(N__32472));
    LocalMux I__4165 (
            .O(N__32472),
            .I(N__32469));
    Span4Mux_v I__4164 (
            .O(N__32469),
            .I(N__32465));
    InMux I__4163 (
            .O(N__32468),
            .I(N__32462));
    Span4Mux_h I__4162 (
            .O(N__32465),
            .I(N__32459));
    LocalMux I__4161 (
            .O(N__32462),
            .I(data_out_frame_13_1));
    Odrv4 I__4160 (
            .O(N__32459),
            .I(data_out_frame_13_1));
    CascadeMux I__4159 (
            .O(N__32454),
            .I(N__32451));
    InMux I__4158 (
            .O(N__32451),
            .I(N__32448));
    LocalMux I__4157 (
            .O(N__32448),
            .I(N__32445));
    Span4Mux_v I__4156 (
            .O(N__32445),
            .I(N__32442));
    Span4Mux_h I__4155 (
            .O(N__32442),
            .I(N__32439));
    Odrv4 I__4154 (
            .O(N__32439),
            .I(\c0.n11_adj_4646 ));
    InMux I__4153 (
            .O(N__32436),
            .I(N__32433));
    LocalMux I__4152 (
            .O(N__32433),
            .I(N__32430));
    Odrv4 I__4151 (
            .O(N__32430),
            .I(\c0.n5_adj_4644 ));
    InMux I__4150 (
            .O(N__32427),
            .I(N__32424));
    LocalMux I__4149 (
            .O(N__32424),
            .I(N__32421));
    Span4Mux_v I__4148 (
            .O(N__32421),
            .I(N__32418));
    Odrv4 I__4147 (
            .O(N__32418),
            .I(\c0.n11_adj_4652 ));
    InMux I__4146 (
            .O(N__32415),
            .I(N__32412));
    LocalMux I__4145 (
            .O(N__32412),
            .I(\c0.data_out_frame_28_2 ));
    InMux I__4144 (
            .O(N__32409),
            .I(N__32406));
    LocalMux I__4143 (
            .O(N__32406),
            .I(N__32403));
    Span4Mux_v I__4142 (
            .O(N__32403),
            .I(N__32400));
    Span4Mux_v I__4141 (
            .O(N__32400),
            .I(N__32397));
    Odrv4 I__4140 (
            .O(N__32397),
            .I(\c0.n26_adj_4651 ));
    CascadeMux I__4139 (
            .O(N__32394),
            .I(N__32391));
    InMux I__4138 (
            .O(N__32391),
            .I(N__32388));
    LocalMux I__4137 (
            .O(N__32388),
            .I(N__32385));
    Odrv4 I__4136 (
            .O(N__32385),
            .I(\quad_counter1.count_direction ));
    InMux I__4135 (
            .O(N__32382),
            .I(N__32379));
    LocalMux I__4134 (
            .O(N__32379),
            .I(N__32376));
    Span4Mux_h I__4133 (
            .O(N__32376),
            .I(N__32373));
    Odrv4 I__4132 (
            .O(N__32373),
            .I(n2291));
    InMux I__4131 (
            .O(N__32370),
            .I(\quad_counter1.n19731 ));
    InMux I__4130 (
            .O(N__32367),
            .I(N__32364));
    LocalMux I__4129 (
            .O(N__32364),
            .I(N__32361));
    Span4Mux_v I__4128 (
            .O(N__32361),
            .I(N__32358));
    Span4Mux_h I__4127 (
            .O(N__32358),
            .I(N__32355));
    Odrv4 I__4126 (
            .O(N__32355),
            .I(n2290));
    InMux I__4125 (
            .O(N__32352),
            .I(\quad_counter1.n19732 ));
    InMux I__4124 (
            .O(N__32349),
            .I(N__32346));
    LocalMux I__4123 (
            .O(N__32346),
            .I(N__32341));
    InMux I__4122 (
            .O(N__32345),
            .I(N__32338));
    InMux I__4121 (
            .O(N__32344),
            .I(N__32335));
    Span4Mux_h I__4120 (
            .O(N__32341),
            .I(N__32330));
    LocalMux I__4119 (
            .O(N__32338),
            .I(N__32330));
    LocalMux I__4118 (
            .O(N__32335),
            .I(N__32327));
    Span4Mux_v I__4117 (
            .O(N__32330),
            .I(N__32324));
    Odrv12 I__4116 (
            .O(N__32327),
            .I(\c0.n13531 ));
    Odrv4 I__4115 (
            .O(N__32324),
            .I(\c0.n13531 ));
    CascadeMux I__4114 (
            .O(N__32319),
            .I(N__32315));
    CascadeMux I__4113 (
            .O(N__32318),
            .I(N__32312));
    InMux I__4112 (
            .O(N__32315),
            .I(N__32309));
    InMux I__4111 (
            .O(N__32312),
            .I(N__32306));
    LocalMux I__4110 (
            .O(N__32309),
            .I(\c0.n20415 ));
    LocalMux I__4109 (
            .O(N__32306),
            .I(\c0.n20415 ));
    InMux I__4108 (
            .O(N__32301),
            .I(N__32298));
    LocalMux I__4107 (
            .O(N__32298),
            .I(N__32294));
    InMux I__4106 (
            .O(N__32297),
            .I(N__32291));
    Odrv4 I__4105 (
            .O(N__32294),
            .I(\c0.n22452 ));
    LocalMux I__4104 (
            .O(N__32291),
            .I(\c0.n22452 ));
    InMux I__4103 (
            .O(N__32286),
            .I(N__32283));
    LocalMux I__4102 (
            .O(N__32283),
            .I(N__32280));
    Odrv4 I__4101 (
            .O(N__32280),
            .I(\c0.n9_adj_4562 ));
    CascadeMux I__4100 (
            .O(N__32277),
            .I(\c0.n10_adj_4690_cascade_ ));
    InMux I__4099 (
            .O(N__32274),
            .I(N__32271));
    LocalMux I__4098 (
            .O(N__32271),
            .I(\c0.n22710 ));
    CascadeMux I__4097 (
            .O(N__32268),
            .I(\c0.n22710_cascade_ ));
    InMux I__4096 (
            .O(N__32265),
            .I(N__32262));
    LocalMux I__4095 (
            .O(N__32262),
            .I(N__32256));
    InMux I__4094 (
            .O(N__32261),
            .I(N__32253));
    InMux I__4093 (
            .O(N__32260),
            .I(N__32248));
    InMux I__4092 (
            .O(N__32259),
            .I(N__32248));
    Span4Mux_h I__4091 (
            .O(N__32256),
            .I(N__32245));
    LocalMux I__4090 (
            .O(N__32253),
            .I(N__32240));
    LocalMux I__4089 (
            .O(N__32248),
            .I(N__32240));
    Odrv4 I__4088 (
            .O(N__32245),
            .I(\c0.n12539 ));
    Odrv12 I__4087 (
            .O(N__32240),
            .I(\c0.n12539 ));
    InMux I__4086 (
            .O(N__32235),
            .I(N__32227));
    InMux I__4085 (
            .O(N__32234),
            .I(N__32227));
    InMux I__4084 (
            .O(N__32233),
            .I(N__32224));
    InMux I__4083 (
            .O(N__32232),
            .I(N__32221));
    LocalMux I__4082 (
            .O(N__32227),
            .I(N__32218));
    LocalMux I__4081 (
            .O(N__32224),
            .I(N__32215));
    LocalMux I__4080 (
            .O(N__32221),
            .I(\c0.n21309 ));
    Odrv12 I__4079 (
            .O(N__32218),
            .I(\c0.n21309 ));
    Odrv4 I__4078 (
            .O(N__32215),
            .I(\c0.n21309 ));
    CascadeMux I__4077 (
            .O(N__32208),
            .I(\c0.n6_adj_4683_cascade_ ));
    CascadeMux I__4076 (
            .O(N__32205),
            .I(N__32202));
    InMux I__4075 (
            .O(N__32202),
            .I(N__32197));
    InMux I__4074 (
            .O(N__32201),
            .I(N__32192));
    InMux I__4073 (
            .O(N__32200),
            .I(N__32192));
    LocalMux I__4072 (
            .O(N__32197),
            .I(N__32189));
    LocalMux I__4071 (
            .O(N__32192),
            .I(N__32186));
    Odrv4 I__4070 (
            .O(N__32189),
            .I(\c0.n13938 ));
    Odrv4 I__4069 (
            .O(N__32186),
            .I(\c0.n13938 ));
    InMux I__4068 (
            .O(N__32181),
            .I(N__32178));
    LocalMux I__4067 (
            .O(N__32178),
            .I(\c0.n12_adj_4688 ));
    InMux I__4066 (
            .O(N__32175),
            .I(N__32172));
    LocalMux I__4065 (
            .O(N__32172),
            .I(\c0.n20360 ));
    InMux I__4064 (
            .O(N__32169),
            .I(N__32163));
    InMux I__4063 (
            .O(N__32168),
            .I(N__32163));
    LocalMux I__4062 (
            .O(N__32163),
            .I(\c0.n22668 ));
    CascadeMux I__4061 (
            .O(N__32160),
            .I(\c0.n20360_cascade_ ));
    InMux I__4060 (
            .O(N__32157),
            .I(N__32154));
    LocalMux I__4059 (
            .O(N__32154),
            .I(\c0.data_out_frame_29_7 ));
    InMux I__4058 (
            .O(N__32151),
            .I(N__32148));
    LocalMux I__4057 (
            .O(N__32148),
            .I(N__32145));
    Odrv12 I__4056 (
            .O(N__32145),
            .I(\c0.n26_adj_4713 ));
    InMux I__4055 (
            .O(N__32142),
            .I(N__32131));
    InMux I__4054 (
            .O(N__32141),
            .I(N__32131));
    InMux I__4053 (
            .O(N__32140),
            .I(N__32131));
    InMux I__4052 (
            .O(N__32139),
            .I(N__32128));
    InMux I__4051 (
            .O(N__32138),
            .I(N__32125));
    LocalMux I__4050 (
            .O(N__32131),
            .I(N__32122));
    LocalMux I__4049 (
            .O(N__32128),
            .I(N__32119));
    LocalMux I__4048 (
            .O(N__32125),
            .I(\c0.n20367 ));
    Odrv4 I__4047 (
            .O(N__32122),
            .I(\c0.n20367 ));
    Odrv4 I__4046 (
            .O(N__32119),
            .I(\c0.n20367 ));
    InMux I__4045 (
            .O(N__32112),
            .I(N__32109));
    LocalMux I__4044 (
            .O(N__32109),
            .I(N__32106));
    Odrv12 I__4043 (
            .O(N__32106),
            .I(\c0.n6_adj_4336 ));
    InMux I__4042 (
            .O(N__32103),
            .I(N__32100));
    LocalMux I__4041 (
            .O(N__32100),
            .I(N__32096));
    InMux I__4040 (
            .O(N__32099),
            .I(N__32093));
    Odrv4 I__4039 (
            .O(N__32096),
            .I(\c0.n22531 ));
    LocalMux I__4038 (
            .O(N__32093),
            .I(\c0.n22531 ));
    InMux I__4037 (
            .O(N__32088),
            .I(N__32085));
    LocalMux I__4036 (
            .O(N__32085),
            .I(N__32082));
    Span4Mux_v I__4035 (
            .O(N__32082),
            .I(N__32079));
    Sp12to4 I__4034 (
            .O(N__32079),
            .I(N__32076));
    Odrv12 I__4033 (
            .O(N__32076),
            .I(n25065));
    InMux I__4032 (
            .O(N__32073),
            .I(N__32070));
    LocalMux I__4031 (
            .O(N__32070),
            .I(\c0.n13741 ));
    CascadeMux I__4030 (
            .O(N__32067),
            .I(\c0.n14_adj_4317_cascade_ ));
    InMux I__4029 (
            .O(N__32064),
            .I(N__32061));
    LocalMux I__4028 (
            .O(N__32061),
            .I(\c0.n15_adj_4318 ));
    InMux I__4027 (
            .O(N__32058),
            .I(N__32055));
    LocalMux I__4026 (
            .O(N__32055),
            .I(\c0.n6_adj_4330 ));
    CascadeMux I__4025 (
            .O(N__32052),
            .I(\c0.n21323_cascade_ ));
    InMux I__4024 (
            .O(N__32049),
            .I(N__32046));
    LocalMux I__4023 (
            .O(N__32046),
            .I(\c0.n14_adj_4368 ));
    CascadeMux I__4022 (
            .O(N__32043),
            .I(\c0.n12488_cascade_ ));
    InMux I__4021 (
            .O(N__32040),
            .I(N__32037));
    LocalMux I__4020 (
            .O(N__32037),
            .I(N__32034));
    Odrv4 I__4019 (
            .O(N__32034),
            .I(\c0.n20379 ));
    CascadeMux I__4018 (
            .O(N__32031),
            .I(\c0.n13531_cascade_ ));
    InMux I__4017 (
            .O(N__32028),
            .I(N__32025));
    LocalMux I__4016 (
            .O(N__32025),
            .I(N__32022));
    Span4Mux_v I__4015 (
            .O(N__32022),
            .I(N__32018));
    InMux I__4014 (
            .O(N__32021),
            .I(N__32015));
    Odrv4 I__4013 (
            .O(N__32018),
            .I(\c0.n22294 ));
    LocalMux I__4012 (
            .O(N__32015),
            .I(\c0.n22294 ));
    InMux I__4011 (
            .O(N__32010),
            .I(\c0.rx.n19718 ));
    CascadeMux I__4010 (
            .O(N__32007),
            .I(N__32004));
    InMux I__4009 (
            .O(N__32004),
            .I(N__31996));
    InMux I__4008 (
            .O(N__32003),
            .I(N__31996));
    InMux I__4007 (
            .O(N__32002),
            .I(N__31993));
    InMux I__4006 (
            .O(N__32001),
            .I(N__31990));
    LocalMux I__4005 (
            .O(N__31996),
            .I(N__31987));
    LocalMux I__4004 (
            .O(N__31993),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__4003 (
            .O(N__31990),
            .I(\c0.rx.r_Clock_Count_4 ));
    Odrv4 I__4002 (
            .O(N__31987),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__4001 (
            .O(N__31980),
            .I(\c0.rx.n19719 ));
    InMux I__4000 (
            .O(N__31977),
            .I(N__31967));
    InMux I__3999 (
            .O(N__31976),
            .I(N__31967));
    InMux I__3998 (
            .O(N__31975),
            .I(N__31967));
    InMux I__3997 (
            .O(N__31974),
            .I(N__31964));
    LocalMux I__3996 (
            .O(N__31967),
            .I(N__31961));
    LocalMux I__3995 (
            .O(N__31964),
            .I(\c0.rx.r_Clock_Count_5 ));
    Odrv4 I__3994 (
            .O(N__31961),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__3993 (
            .O(N__31956),
            .I(\c0.rx.n19720 ));
    InMux I__3992 (
            .O(N__31953),
            .I(N__31950));
    LocalMux I__3991 (
            .O(N__31950),
            .I(N__31944));
    InMux I__3990 (
            .O(N__31949),
            .I(N__31939));
    InMux I__3989 (
            .O(N__31948),
            .I(N__31939));
    InMux I__3988 (
            .O(N__31947),
            .I(N__31936));
    Span4Mux_v I__3987 (
            .O(N__31944),
            .I(N__31933));
    LocalMux I__3986 (
            .O(N__31939),
            .I(N__31930));
    LocalMux I__3985 (
            .O(N__31936),
            .I(\c0.rx.r_Clock_Count_6 ));
    Odrv4 I__3984 (
            .O(N__31933),
            .I(\c0.rx.r_Clock_Count_6 ));
    Odrv4 I__3983 (
            .O(N__31930),
            .I(\c0.rx.r_Clock_Count_6 ));
    InMux I__3982 (
            .O(N__31923),
            .I(\c0.rx.n19721 ));
    InMux I__3981 (
            .O(N__31920),
            .I(\c0.rx.n19722 ));
    InMux I__3980 (
            .O(N__31917),
            .I(N__31914));
    LocalMux I__3979 (
            .O(N__31914),
            .I(N__31911));
    Span4Mux_h I__3978 (
            .O(N__31911),
            .I(N__31908));
    Span4Mux_v I__3977 (
            .O(N__31908),
            .I(N__31904));
    InMux I__3976 (
            .O(N__31907),
            .I(N__31901));
    Sp12to4 I__3975 (
            .O(N__31904),
            .I(N__31895));
    LocalMux I__3974 (
            .O(N__31901),
            .I(N__31891));
    InMux I__3973 (
            .O(N__31900),
            .I(N__31888));
    InMux I__3972 (
            .O(N__31899),
            .I(N__31885));
    InMux I__3971 (
            .O(N__31898),
            .I(N__31882));
    Span12Mux_v I__3970 (
            .O(N__31895),
            .I(N__31879));
    InMux I__3969 (
            .O(N__31894),
            .I(N__31876));
    Span4Mux_v I__3968 (
            .O(N__31891),
            .I(N__31871));
    LocalMux I__3967 (
            .O(N__31888),
            .I(N__31871));
    LocalMux I__3966 (
            .O(N__31885),
            .I(N__31868));
    LocalMux I__3965 (
            .O(N__31882),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv12 I__3964 (
            .O(N__31879),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__3963 (
            .O(N__31876),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__3962 (
            .O(N__31871),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__3961 (
            .O(N__31868),
            .I(\c0.rx.r_Clock_Count_7 ));
    SRMux I__3960 (
            .O(N__31857),
            .I(N__31854));
    LocalMux I__3959 (
            .O(N__31854),
            .I(N__31851));
    Span4Mux_h I__3958 (
            .O(N__31851),
            .I(N__31848));
    Odrv4 I__3957 (
            .O(N__31848),
            .I(n14895));
    SRMux I__3956 (
            .O(N__31845),
            .I(N__31842));
    LocalMux I__3955 (
            .O(N__31842),
            .I(N__31839));
    Odrv4 I__3954 (
            .O(N__31839),
            .I(\c0.n21645 ));
    CascadeMux I__3953 (
            .O(N__31836),
            .I(\c0.n22638_cascade_ ));
    CascadeMux I__3952 (
            .O(N__31833),
            .I(n14895_cascade_));
    CascadeMux I__3951 (
            .O(N__31830),
            .I(n24921_cascade_));
    InMux I__3950 (
            .O(N__31827),
            .I(N__31824));
    LocalMux I__3949 (
            .O(N__31824),
            .I(N__31821));
    Odrv12 I__3948 (
            .O(N__31821),
            .I(n24922));
    InMux I__3947 (
            .O(N__31818),
            .I(N__31815));
    LocalMux I__3946 (
            .O(N__31815),
            .I(\c0.rx.n24916 ));
    InMux I__3945 (
            .O(N__31812),
            .I(N__31809));
    LocalMux I__3944 (
            .O(N__31809),
            .I(\c0.rx.n8 ));
    InMux I__3943 (
            .O(N__31806),
            .I(N__31800));
    InMux I__3942 (
            .O(N__31805),
            .I(N__31797));
    InMux I__3941 (
            .O(N__31804),
            .I(N__31792));
    InMux I__3940 (
            .O(N__31803),
            .I(N__31792));
    LocalMux I__3939 (
            .O(N__31800),
            .I(r_Clock_Count_0));
    LocalMux I__3938 (
            .O(N__31797),
            .I(r_Clock_Count_0));
    LocalMux I__3937 (
            .O(N__31792),
            .I(r_Clock_Count_0));
    InMux I__3936 (
            .O(N__31785),
            .I(N__31782));
    LocalMux I__3935 (
            .O(N__31782),
            .I(n226));
    InMux I__3934 (
            .O(N__31779),
            .I(bfn_11_26_0_));
    InMux I__3933 (
            .O(N__31776),
            .I(N__31768));
    InMux I__3932 (
            .O(N__31775),
            .I(N__31768));
    InMux I__3931 (
            .O(N__31774),
            .I(N__31765));
    InMux I__3930 (
            .O(N__31773),
            .I(N__31762));
    LocalMux I__3929 (
            .O(N__31768),
            .I(N__31759));
    LocalMux I__3928 (
            .O(N__31765),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__3927 (
            .O(N__31762),
            .I(\c0.rx.r_Clock_Count_1 ));
    Odrv4 I__3926 (
            .O(N__31759),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__3925 (
            .O(N__31752),
            .I(\c0.rx.n19716 ));
    InMux I__3924 (
            .O(N__31749),
            .I(N__31743));
    InMux I__3923 (
            .O(N__31748),
            .I(N__31740));
    InMux I__3922 (
            .O(N__31747),
            .I(N__31735));
    InMux I__3921 (
            .O(N__31746),
            .I(N__31735));
    LocalMux I__3920 (
            .O(N__31743),
            .I(N__31732));
    LocalMux I__3919 (
            .O(N__31740),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__3918 (
            .O(N__31735),
            .I(\c0.rx.r_Clock_Count_2 ));
    Odrv4 I__3917 (
            .O(N__31732),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__3916 (
            .O(N__31725),
            .I(\c0.rx.n19717 ));
    InMux I__3915 (
            .O(N__31722),
            .I(N__31717));
    CascadeMux I__3914 (
            .O(N__31721),
            .I(N__31714));
    InMux I__3913 (
            .O(N__31720),
            .I(N__31710));
    LocalMux I__3912 (
            .O(N__31717),
            .I(N__31707));
    InMux I__3911 (
            .O(N__31714),
            .I(N__31702));
    InMux I__3910 (
            .O(N__31713),
            .I(N__31702));
    LocalMux I__3909 (
            .O(N__31710),
            .I(\c0.rx.r_Clock_Count_3 ));
    Odrv4 I__3908 (
            .O(N__31707),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__3907 (
            .O(N__31702),
            .I(\c0.rx.r_Clock_Count_3 ));
    CascadeMux I__3906 (
            .O(N__31695),
            .I(\c0.rx.n9_cascade_ ));
    InMux I__3905 (
            .O(N__31692),
            .I(N__31688));
    InMux I__3904 (
            .O(N__31691),
            .I(N__31684));
    LocalMux I__3903 (
            .O(N__31688),
            .I(N__31681));
    InMux I__3902 (
            .O(N__31687),
            .I(N__31678));
    LocalMux I__3901 (
            .O(N__31684),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__3900 (
            .O(N__31681),
            .I(\c0.FRAME_MATCHER_state_30 ));
    LocalMux I__3899 (
            .O(N__31678),
            .I(\c0.FRAME_MATCHER_state_30 ));
    CascadeMux I__3898 (
            .O(N__31671),
            .I(\c0.rx.n17531_cascade_ ));
    InMux I__3897 (
            .O(N__31668),
            .I(N__31665));
    LocalMux I__3896 (
            .O(N__31665),
            .I(\c0.rx.n17590 ));
    InMux I__3895 (
            .O(N__31662),
            .I(N__31659));
    LocalMux I__3894 (
            .O(N__31659),
            .I(N__31655));
    InMux I__3893 (
            .O(N__31658),
            .I(N__31651));
    Sp12to4 I__3892 (
            .O(N__31655),
            .I(N__31648));
    InMux I__3891 (
            .O(N__31654),
            .I(N__31645));
    LocalMux I__3890 (
            .O(N__31651),
            .I(N__31642));
    Span12Mux_v I__3889 (
            .O(N__31648),
            .I(N__31639));
    LocalMux I__3888 (
            .O(N__31645),
            .I(N__31636));
    Span4Mux_h I__3887 (
            .O(N__31642),
            .I(N__31633));
    Odrv12 I__3886 (
            .O(N__31639),
            .I(\c0.rx.n17848 ));
    Odrv4 I__3885 (
            .O(N__31636),
            .I(\c0.rx.n17848 ));
    Odrv4 I__3884 (
            .O(N__31633),
            .I(\c0.rx.n17848 ));
    InMux I__3883 (
            .O(N__31626),
            .I(N__31623));
    LocalMux I__3882 (
            .O(N__31623),
            .I(\c0.rx.n14 ));
    CascadeMux I__3881 (
            .O(N__31620),
            .I(\c0.rx.n24697_cascade_ ));
    CascadeMux I__3880 (
            .O(N__31617),
            .I(\c0.rx.n24914_cascade_ ));
    CascadeMux I__3879 (
            .O(N__31614),
            .I(N__31611));
    InMux I__3878 (
            .O(N__31611),
            .I(N__31608));
    LocalMux I__3877 (
            .O(N__31608),
            .I(\c0.n24255 ));
    SRMux I__3876 (
            .O(N__31605),
            .I(N__31602));
    LocalMux I__3875 (
            .O(N__31602),
            .I(N__31599));
    Sp12to4 I__3874 (
            .O(N__31599),
            .I(N__31596));
    Odrv12 I__3873 (
            .O(N__31596),
            .I(\c0.n21583 ));
    InMux I__3872 (
            .O(N__31593),
            .I(N__31589));
    InMux I__3871 (
            .O(N__31592),
            .I(N__31586));
    LocalMux I__3870 (
            .O(N__31589),
            .I(N__31582));
    LocalMux I__3869 (
            .O(N__31586),
            .I(N__31579));
    InMux I__3868 (
            .O(N__31585),
            .I(N__31576));
    Span4Mux_h I__3867 (
            .O(N__31582),
            .I(N__31573));
    Span4Mux_h I__3866 (
            .O(N__31579),
            .I(N__31570));
    LocalMux I__3865 (
            .O(N__31576),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv4 I__3864 (
            .O(N__31573),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv4 I__3863 (
            .O(N__31570),
            .I(\c0.FRAME_MATCHER_state_26 ));
    InMux I__3862 (
            .O(N__31563),
            .I(N__31560));
    LocalMux I__3861 (
            .O(N__31560),
            .I(N__31555));
    InMux I__3860 (
            .O(N__31559),
            .I(N__31552));
    InMux I__3859 (
            .O(N__31558),
            .I(N__31549));
    Span4Mux_h I__3858 (
            .O(N__31555),
            .I(N__31546));
    LocalMux I__3857 (
            .O(N__31552),
            .I(\c0.FRAME_MATCHER_state_17 ));
    LocalMux I__3856 (
            .O(N__31549),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__3855 (
            .O(N__31546),
            .I(\c0.FRAME_MATCHER_state_17 ));
    CascadeMux I__3854 (
            .O(N__31539),
            .I(\c0.n14530_cascade_ ));
    CascadeMux I__3853 (
            .O(N__31536),
            .I(N__31533));
    InMux I__3852 (
            .O(N__31533),
            .I(N__31529));
    InMux I__3851 (
            .O(N__31532),
            .I(N__31526));
    LocalMux I__3850 (
            .O(N__31529),
            .I(N__31523));
    LocalMux I__3849 (
            .O(N__31526),
            .I(data_out_frame_11_6));
    Odrv12 I__3848 (
            .O(N__31523),
            .I(data_out_frame_11_6));
    CascadeMux I__3847 (
            .O(N__31518),
            .I(\c0.n25098_cascade_ ));
    InMux I__3846 (
            .O(N__31515),
            .I(N__31512));
    LocalMux I__3845 (
            .O(N__31512),
            .I(\c0.n25101 ));
    CascadeMux I__3844 (
            .O(N__31509),
            .I(N__31506));
    InMux I__3843 (
            .O(N__31506),
            .I(N__31500));
    InMux I__3842 (
            .O(N__31505),
            .I(N__31500));
    LocalMux I__3841 (
            .O(N__31500),
            .I(data_out_frame_6_5));
    CascadeMux I__3840 (
            .O(N__31497),
            .I(N__31494));
    InMux I__3839 (
            .O(N__31494),
            .I(N__31490));
    InMux I__3838 (
            .O(N__31493),
            .I(N__31487));
    LocalMux I__3837 (
            .O(N__31490),
            .I(data_out_frame_5_5));
    LocalMux I__3836 (
            .O(N__31487),
            .I(data_out_frame_5_5));
    InMux I__3835 (
            .O(N__31482),
            .I(N__31479));
    LocalMux I__3834 (
            .O(N__31479),
            .I(\c0.n5_adj_4679 ));
    CascadeMux I__3833 (
            .O(N__31476),
            .I(\c0.n25016_cascade_ ));
    InMux I__3832 (
            .O(N__31473),
            .I(N__31470));
    LocalMux I__3831 (
            .O(N__31470),
            .I(N__31467));
    Odrv4 I__3830 (
            .O(N__31467),
            .I(\c0.n24794 ));
    InMux I__3829 (
            .O(N__31464),
            .I(N__31461));
    LocalMux I__3828 (
            .O(N__31461),
            .I(\c0.n5_adj_4700 ));
    InMux I__3827 (
            .O(N__31458),
            .I(N__31454));
    InMux I__3826 (
            .O(N__31457),
            .I(N__31451));
    LocalMux I__3825 (
            .O(N__31454),
            .I(data_out_frame_10_2));
    LocalMux I__3824 (
            .O(N__31451),
            .I(data_out_frame_10_2));
    CascadeMux I__3823 (
            .O(N__31446),
            .I(N__31442));
    InMux I__3822 (
            .O(N__31445),
            .I(N__31437));
    InMux I__3821 (
            .O(N__31442),
            .I(N__31437));
    LocalMux I__3820 (
            .O(N__31437),
            .I(data_out_frame_11_0));
    CascadeMux I__3819 (
            .O(N__31434),
            .I(N__31431));
    InMux I__3818 (
            .O(N__31431),
            .I(N__31428));
    LocalMux I__3817 (
            .O(N__31428),
            .I(N__31425));
    Odrv4 I__3816 (
            .O(N__31425),
            .I(\c0.n11_adj_4703 ));
    CascadeMux I__3815 (
            .O(N__31422),
            .I(\c0.n24945_cascade_ ));
    CascadeMux I__3814 (
            .O(N__31419),
            .I(N__31412));
    InMux I__3813 (
            .O(N__31418),
            .I(N__31409));
    CascadeMux I__3812 (
            .O(N__31417),
            .I(N__31406));
    CascadeMux I__3811 (
            .O(N__31416),
            .I(N__31402));
    InMux I__3810 (
            .O(N__31415),
            .I(N__31396));
    InMux I__3809 (
            .O(N__31412),
            .I(N__31396));
    LocalMux I__3808 (
            .O(N__31409),
            .I(N__31392));
    InMux I__3807 (
            .O(N__31406),
            .I(N__31389));
    InMux I__3806 (
            .O(N__31405),
            .I(N__31386));
    InMux I__3805 (
            .O(N__31402),
            .I(N__31381));
    InMux I__3804 (
            .O(N__31401),
            .I(N__31381));
    LocalMux I__3803 (
            .O(N__31396),
            .I(N__31378));
    CascadeMux I__3802 (
            .O(N__31395),
            .I(N__31375));
    Span4Mux_v I__3801 (
            .O(N__31392),
            .I(N__31372));
    LocalMux I__3800 (
            .O(N__31389),
            .I(N__31369));
    LocalMux I__3799 (
            .O(N__31386),
            .I(N__31366));
    LocalMux I__3798 (
            .O(N__31381),
            .I(N__31363));
    Span4Mux_v I__3797 (
            .O(N__31378),
            .I(N__31360));
    InMux I__3796 (
            .O(N__31375),
            .I(N__31357));
    Span4Mux_h I__3795 (
            .O(N__31372),
            .I(N__31352));
    Span4Mux_v I__3794 (
            .O(N__31369),
            .I(N__31352));
    Span4Mux_v I__3793 (
            .O(N__31366),
            .I(N__31347));
    Span4Mux_v I__3792 (
            .O(N__31363),
            .I(N__31347));
    Span4Mux_v I__3791 (
            .O(N__31360),
            .I(N__31344));
    LocalMux I__3790 (
            .O(N__31357),
            .I(N__31341));
    Odrv4 I__3789 (
            .O(N__31352),
            .I(n24682));
    Odrv4 I__3788 (
            .O(N__31347),
            .I(n24682));
    Odrv4 I__3787 (
            .O(N__31344),
            .I(n24682));
    Odrv12 I__3786 (
            .O(N__31341),
            .I(n24682));
    CascadeMux I__3785 (
            .O(N__31332),
            .I(\c0.n24797_cascade_ ));
    CascadeMux I__3784 (
            .O(N__31329),
            .I(N__31325));
    InMux I__3783 (
            .O(N__31328),
            .I(N__31320));
    InMux I__3782 (
            .O(N__31325),
            .I(N__31305));
    InMux I__3781 (
            .O(N__31324),
            .I(N__31305));
    InMux I__3780 (
            .O(N__31323),
            .I(N__31305));
    LocalMux I__3779 (
            .O(N__31320),
            .I(N__31300));
    InMux I__3778 (
            .O(N__31319),
            .I(N__31297));
    CascadeMux I__3777 (
            .O(N__31318),
            .I(N__31294));
    InMux I__3776 (
            .O(N__31317),
            .I(N__31291));
    InMux I__3775 (
            .O(N__31316),
            .I(N__31286));
    InMux I__3774 (
            .O(N__31315),
            .I(N__31286));
    InMux I__3773 (
            .O(N__31314),
            .I(N__31281));
    InMux I__3772 (
            .O(N__31313),
            .I(N__31281));
    InMux I__3771 (
            .O(N__31312),
            .I(N__31278));
    LocalMux I__3770 (
            .O(N__31305),
            .I(N__31275));
    CascadeMux I__3769 (
            .O(N__31304),
            .I(N__31272));
    CascadeMux I__3768 (
            .O(N__31303),
            .I(N__31267));
    Span4Mux_h I__3767 (
            .O(N__31300),
            .I(N__31261));
    LocalMux I__3766 (
            .O(N__31297),
            .I(N__31261));
    InMux I__3765 (
            .O(N__31294),
            .I(N__31258));
    LocalMux I__3764 (
            .O(N__31291),
            .I(N__31255));
    LocalMux I__3763 (
            .O(N__31286),
            .I(N__31248));
    LocalMux I__3762 (
            .O(N__31281),
            .I(N__31248));
    LocalMux I__3761 (
            .O(N__31278),
            .I(N__31248));
    Span4Mux_v I__3760 (
            .O(N__31275),
            .I(N__31245));
    InMux I__3759 (
            .O(N__31272),
            .I(N__31242));
    InMux I__3758 (
            .O(N__31271),
            .I(N__31237));
    InMux I__3757 (
            .O(N__31270),
            .I(N__31237));
    InMux I__3756 (
            .O(N__31267),
            .I(N__31234));
    InMux I__3755 (
            .O(N__31266),
            .I(N__31231));
    Span4Mux_v I__3754 (
            .O(N__31261),
            .I(N__31226));
    LocalMux I__3753 (
            .O(N__31258),
            .I(N__31226));
    Span4Mux_v I__3752 (
            .O(N__31255),
            .I(N__31219));
    Span4Mux_v I__3751 (
            .O(N__31248),
            .I(N__31219));
    Span4Mux_v I__3750 (
            .O(N__31245),
            .I(N__31219));
    LocalMux I__3749 (
            .O(N__31242),
            .I(N__31214));
    LocalMux I__3748 (
            .O(N__31237),
            .I(N__31214));
    LocalMux I__3747 (
            .O(N__31234),
            .I(N__31211));
    LocalMux I__3746 (
            .O(N__31231),
            .I(byte_transmit_counter_4));
    Odrv4 I__3745 (
            .O(N__31226),
            .I(byte_transmit_counter_4));
    Odrv4 I__3744 (
            .O(N__31219),
            .I(byte_transmit_counter_4));
    Odrv12 I__3743 (
            .O(N__31214),
            .I(byte_transmit_counter_4));
    Odrv4 I__3742 (
            .O(N__31211),
            .I(byte_transmit_counter_4));
    InMux I__3741 (
            .O(N__31200),
            .I(N__31194));
    InMux I__3740 (
            .O(N__31199),
            .I(N__31191));
    InMux I__3739 (
            .O(N__31198),
            .I(N__31186));
    InMux I__3738 (
            .O(N__31197),
            .I(N__31183));
    LocalMux I__3737 (
            .O(N__31194),
            .I(N__31178));
    LocalMux I__3736 (
            .O(N__31191),
            .I(N__31178));
    InMux I__3735 (
            .O(N__31190),
            .I(N__31173));
    InMux I__3734 (
            .O(N__31189),
            .I(N__31170));
    LocalMux I__3733 (
            .O(N__31186),
            .I(N__31167));
    LocalMux I__3732 (
            .O(N__31183),
            .I(N__31162));
    Span4Mux_h I__3731 (
            .O(N__31178),
            .I(N__31162));
    InMux I__3730 (
            .O(N__31177),
            .I(N__31159));
    InMux I__3729 (
            .O(N__31176),
            .I(N__31153));
    LocalMux I__3728 (
            .O(N__31173),
            .I(N__31150));
    LocalMux I__3727 (
            .O(N__31170),
            .I(N__31147));
    Span4Mux_v I__3726 (
            .O(N__31167),
            .I(N__31140));
    Span4Mux_v I__3725 (
            .O(N__31162),
            .I(N__31140));
    LocalMux I__3724 (
            .O(N__31159),
            .I(N__31140));
    InMux I__3723 (
            .O(N__31158),
            .I(N__31137));
    InMux I__3722 (
            .O(N__31157),
            .I(N__31134));
    InMux I__3721 (
            .O(N__31156),
            .I(N__31131));
    LocalMux I__3720 (
            .O(N__31153),
            .I(N__31128));
    Span4Mux_h I__3719 (
            .O(N__31150),
            .I(N__31125));
    Span4Mux_v I__3718 (
            .O(N__31147),
            .I(N__31120));
    Span4Mux_v I__3717 (
            .O(N__31140),
            .I(N__31120));
    LocalMux I__3716 (
            .O(N__31137),
            .I(N__31115));
    LocalMux I__3715 (
            .O(N__31134),
            .I(N__31115));
    LocalMux I__3714 (
            .O(N__31131),
            .I(byte_transmit_counter_3));
    Odrv12 I__3713 (
            .O(N__31128),
            .I(byte_transmit_counter_3));
    Odrv4 I__3712 (
            .O(N__31125),
            .I(byte_transmit_counter_3));
    Odrv4 I__3711 (
            .O(N__31120),
            .I(byte_transmit_counter_3));
    Odrv4 I__3710 (
            .O(N__31115),
            .I(byte_transmit_counter_3));
    CascadeMux I__3709 (
            .O(N__31104),
            .I(n24799_cascade_));
    InMux I__3708 (
            .O(N__31101),
            .I(N__31098));
    LocalMux I__3707 (
            .O(N__31098),
            .I(n25012));
    InMux I__3706 (
            .O(N__31095),
            .I(N__31092));
    LocalMux I__3705 (
            .O(N__31092),
            .I(N__31089));
    Span4Mux_h I__3704 (
            .O(N__31089),
            .I(N__31086));
    Odrv4 I__3703 (
            .O(N__31086),
            .I(n10_adj_4775));
    CascadeMux I__3702 (
            .O(N__31083),
            .I(N__31080));
    InMux I__3701 (
            .O(N__31080),
            .I(N__31077));
    LocalMux I__3700 (
            .O(N__31077),
            .I(N__31074));
    Odrv4 I__3699 (
            .O(N__31074),
            .I(\c0.n24953 ));
    InMux I__3698 (
            .O(N__31071),
            .I(N__31068));
    LocalMux I__3697 (
            .O(N__31068),
            .I(N__31065));
    Span4Mux_h I__3696 (
            .O(N__31065),
            .I(N__31062));
    Odrv4 I__3695 (
            .O(N__31062),
            .I(\c0.n24803 ));
    CascadeMux I__3694 (
            .O(N__31059),
            .I(N__31055));
    InMux I__3693 (
            .O(N__31058),
            .I(N__31052));
    InMux I__3692 (
            .O(N__31055),
            .I(N__31049));
    LocalMux I__3691 (
            .O(N__31052),
            .I(data_out_frame_8_2));
    LocalMux I__3690 (
            .O(N__31049),
            .I(data_out_frame_8_2));
    CascadeMux I__3689 (
            .O(N__31044),
            .I(\c0.n25059_cascade_ ));
    CascadeMux I__3688 (
            .O(N__31041),
            .I(n25004_cascade_));
    InMux I__3687 (
            .O(N__31038),
            .I(N__31035));
    LocalMux I__3686 (
            .O(N__31035),
            .I(N__31032));
    Odrv4 I__3685 (
            .O(N__31032),
            .I(n10_adj_4778));
    InMux I__3684 (
            .O(N__31029),
            .I(N__31026));
    LocalMux I__3683 (
            .O(N__31026),
            .I(\c0.n24809 ));
    InMux I__3682 (
            .O(N__31023),
            .I(N__31020));
    LocalMux I__3681 (
            .O(N__31020),
            .I(n24811));
    InMux I__3680 (
            .O(N__31017),
            .I(N__31014));
    LocalMux I__3679 (
            .O(N__31014),
            .I(N__31011));
    Span4Mux_v I__3678 (
            .O(N__31011),
            .I(N__31008));
    Odrv4 I__3677 (
            .O(N__31008),
            .I(n24904));
    CascadeMux I__3676 (
            .O(N__31005),
            .I(N__31001));
    InMux I__3675 (
            .O(N__31004),
            .I(N__30998));
    InMux I__3674 (
            .O(N__31001),
            .I(N__30995));
    LocalMux I__3673 (
            .O(N__30998),
            .I(N__30992));
    LocalMux I__3672 (
            .O(N__30995),
            .I(N__30989));
    Span4Mux_h I__3671 (
            .O(N__30992),
            .I(N__30986));
    Odrv12 I__3670 (
            .O(N__30989),
            .I(data_out_frame_28_3));
    Odrv4 I__3669 (
            .O(N__30986),
            .I(data_out_frame_28_3));
    CascadeMux I__3668 (
            .O(N__30981),
            .I(\c0.n25110_cascade_ ));
    InMux I__3667 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__3666 (
            .O(N__30975),
            .I(\c0.n25113 ));
    InMux I__3665 (
            .O(N__30972),
            .I(N__30969));
    LocalMux I__3664 (
            .O(N__30969),
            .I(\c0.n25056 ));
    InMux I__3663 (
            .O(N__30966),
            .I(N__30963));
    LocalMux I__3662 (
            .O(N__30963),
            .I(N__30959));
    InMux I__3661 (
            .O(N__30962),
            .I(N__30956));
    Span12Mux_s10_h I__3660 (
            .O(N__30959),
            .I(N__30953));
    LocalMux I__3659 (
            .O(N__30956),
            .I(data_out_frame_10_3));
    Odrv12 I__3658 (
            .O(N__30953),
            .I(data_out_frame_10_3));
    CascadeMux I__3657 (
            .O(N__30948),
            .I(N__30945));
    InMux I__3656 (
            .O(N__30945),
            .I(N__30942));
    LocalMux I__3655 (
            .O(N__30942),
            .I(N__30938));
    InMux I__3654 (
            .O(N__30941),
            .I(N__30935));
    Span4Mux_v I__3653 (
            .O(N__30938),
            .I(N__30932));
    LocalMux I__3652 (
            .O(N__30935),
            .I(\c0.n21362 ));
    Odrv4 I__3651 (
            .O(N__30932),
            .I(\c0.n21362 ));
    CascadeMux I__3650 (
            .O(N__30927),
            .I(N__30924));
    InMux I__3649 (
            .O(N__30924),
            .I(N__30921));
    LocalMux I__3648 (
            .O(N__30921),
            .I(N__30918));
    Odrv4 I__3647 (
            .O(N__30918),
            .I(\c0.n11_adj_4572 ));
    CascadeMux I__3646 (
            .O(N__30915),
            .I(N__30912));
    InMux I__3645 (
            .O(N__30912),
            .I(N__30906));
    InMux I__3644 (
            .O(N__30911),
            .I(N__30906));
    LocalMux I__3643 (
            .O(N__30906),
            .I(data_out_frame_13_0));
    InMux I__3642 (
            .O(N__30903),
            .I(N__30899));
    InMux I__3641 (
            .O(N__30902),
            .I(N__30896));
    LocalMux I__3640 (
            .O(N__30899),
            .I(N__30893));
    LocalMux I__3639 (
            .O(N__30896),
            .I(data_out_frame_6_2));
    Odrv4 I__3638 (
            .O(N__30893),
            .I(data_out_frame_6_2));
    CascadeMux I__3637 (
            .O(N__30888),
            .I(\c0.n5_adj_4650_cascade_ ));
    InMux I__3636 (
            .O(N__30885),
            .I(N__30882));
    LocalMux I__3635 (
            .O(N__30882),
            .I(N__30879));
    Odrv12 I__3634 (
            .O(N__30879),
            .I(\c0.n6_adj_4649 ));
    CascadeMux I__3633 (
            .O(N__30876),
            .I(n22735_cascade_));
    CascadeMux I__3632 (
            .O(N__30873),
            .I(N__30870));
    InMux I__3631 (
            .O(N__30870),
            .I(N__30867));
    LocalMux I__3630 (
            .O(N__30867),
            .I(\c0.n22757 ));
    CascadeMux I__3629 (
            .O(N__30864),
            .I(\c0.n20_adj_4699_cascade_ ));
    InMux I__3628 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__3627 (
            .O(N__30858),
            .I(n22285));
    InMux I__3626 (
            .O(N__30855),
            .I(N__30852));
    LocalMux I__3625 (
            .O(N__30852),
            .I(N__30849));
    Odrv4 I__3624 (
            .O(N__30849),
            .I(\c0.n6_adj_4210 ));
    InMux I__3623 (
            .O(N__30846),
            .I(N__30839));
    InMux I__3622 (
            .O(N__30845),
            .I(N__30839));
    InMux I__3621 (
            .O(N__30844),
            .I(N__30836));
    LocalMux I__3620 (
            .O(N__30839),
            .I(\c0.n13683 ));
    LocalMux I__3619 (
            .O(N__30836),
            .I(\c0.n13683 ));
    CascadeMux I__3618 (
            .O(N__30831),
            .I(\c0.n22534_cascade_ ));
    CascadeMux I__3617 (
            .O(N__30828),
            .I(\c0.n20415_cascade_ ));
    InMux I__3616 (
            .O(N__30825),
            .I(N__30820));
    InMux I__3615 (
            .O(N__30824),
            .I(N__30815));
    InMux I__3614 (
            .O(N__30823),
            .I(N__30815));
    LocalMux I__3613 (
            .O(N__30820),
            .I(\c0.n20384 ));
    LocalMux I__3612 (
            .O(N__30815),
            .I(\c0.n20384 ));
    CascadeMux I__3611 (
            .O(N__30810),
            .I(N__30806));
    InMux I__3610 (
            .O(N__30809),
            .I(N__30803));
    InMux I__3609 (
            .O(N__30806),
            .I(N__30800));
    LocalMux I__3608 (
            .O(N__30803),
            .I(\c0.n22544 ));
    LocalMux I__3607 (
            .O(N__30800),
            .I(\c0.n22544 ));
    CascadeMux I__3606 (
            .O(N__30795),
            .I(N__30792));
    InMux I__3605 (
            .O(N__30792),
            .I(N__30789));
    LocalMux I__3604 (
            .O(N__30789),
            .I(\c0.data_out_frame_28_5 ));
    InMux I__3603 (
            .O(N__30786),
            .I(N__30783));
    LocalMux I__3602 (
            .O(N__30783),
            .I(N__30780));
    Span4Mux_v I__3601 (
            .O(N__30780),
            .I(N__30777));
    Odrv4 I__3600 (
            .O(N__30777),
            .I(\c0.n26_adj_4680 ));
    InMux I__3599 (
            .O(N__30774),
            .I(N__30767));
    InMux I__3598 (
            .O(N__30773),
            .I(N__30767));
    InMux I__3597 (
            .O(N__30772),
            .I(N__30764));
    LocalMux I__3596 (
            .O(N__30767),
            .I(\c0.n22478 ));
    LocalMux I__3595 (
            .O(N__30764),
            .I(\c0.n22478 ));
    InMux I__3594 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__3593 (
            .O(N__30756),
            .I(n22735));
    InMux I__3592 (
            .O(N__30753),
            .I(N__30750));
    LocalMux I__3591 (
            .O(N__30750),
            .I(\c0.n6_adj_4456 ));
    CascadeMux I__3590 (
            .O(N__30747),
            .I(n21484_cascade_));
    InMux I__3589 (
            .O(N__30744),
            .I(N__30740));
    InMux I__3588 (
            .O(N__30743),
            .I(N__30737));
    LocalMux I__3587 (
            .O(N__30740),
            .I(\c0.n22246 ));
    LocalMux I__3586 (
            .O(N__30737),
            .I(\c0.n22246 ));
    InMux I__3585 (
            .O(N__30732),
            .I(N__30728));
    InMux I__3584 (
            .O(N__30731),
            .I(N__30725));
    LocalMux I__3583 (
            .O(N__30728),
            .I(N__30722));
    LocalMux I__3582 (
            .O(N__30725),
            .I(data_out_frame_7_3));
    Odrv4 I__3581 (
            .O(N__30722),
            .I(data_out_frame_7_3));
    InMux I__3580 (
            .O(N__30717),
            .I(N__30714));
    LocalMux I__3579 (
            .O(N__30714),
            .I(\c0.n10_adj_4313 ));
    CascadeMux I__3578 (
            .O(N__30711),
            .I(N__30708));
    InMux I__3577 (
            .O(N__30708),
            .I(N__30705));
    LocalMux I__3576 (
            .O(N__30705),
            .I(N__30701));
    InMux I__3575 (
            .O(N__30704),
            .I(N__30698));
    Span4Mux_v I__3574 (
            .O(N__30701),
            .I(N__30695));
    LocalMux I__3573 (
            .O(N__30698),
            .I(data_out_frame_11_3));
    Odrv4 I__3572 (
            .O(N__30695),
            .I(data_out_frame_11_3));
    InMux I__3571 (
            .O(N__30690),
            .I(N__30687));
    LocalMux I__3570 (
            .O(N__30687),
            .I(\c0.n22534 ));
    CascadeMux I__3569 (
            .O(N__30684),
            .I(\c0.n22246_cascade_ ));
    InMux I__3568 (
            .O(N__30681),
            .I(N__30677));
    InMux I__3567 (
            .O(N__30680),
            .I(N__30674));
    LocalMux I__3566 (
            .O(N__30677),
            .I(N__30671));
    LocalMux I__3565 (
            .O(N__30674),
            .I(\c0.n22846 ));
    Odrv4 I__3564 (
            .O(N__30671),
            .I(\c0.n22846 ));
    CascadeMux I__3563 (
            .O(N__30666),
            .I(\c0.n20379_cascade_ ));
    InMux I__3562 (
            .O(N__30663),
            .I(N__30660));
    LocalMux I__3561 (
            .O(N__30660),
            .I(N__30653));
    InMux I__3560 (
            .O(N__30659),
            .I(N__30646));
    InMux I__3559 (
            .O(N__30658),
            .I(N__30646));
    InMux I__3558 (
            .O(N__30657),
            .I(N__30646));
    InMux I__3557 (
            .O(N__30656),
            .I(N__30643));
    Span4Mux_v I__3556 (
            .O(N__30653),
            .I(N__30640));
    LocalMux I__3555 (
            .O(N__30646),
            .I(N__30637));
    LocalMux I__3554 (
            .O(N__30643),
            .I(A_filtered_adj_4763));
    Odrv4 I__3553 (
            .O(N__30640),
            .I(A_filtered_adj_4763));
    Odrv12 I__3552 (
            .O(N__30637),
            .I(A_filtered_adj_4763));
    InMux I__3551 (
            .O(N__30630),
            .I(N__30627));
    LocalMux I__3550 (
            .O(N__30627),
            .I(N__30624));
    Span4Mux_v I__3549 (
            .O(N__30624),
            .I(N__30619));
    InMux I__3548 (
            .O(N__30623),
            .I(N__30614));
    InMux I__3547 (
            .O(N__30622),
            .I(N__30614));
    Odrv4 I__3546 (
            .O(N__30619),
            .I(\quad_counter1.B_delayed ));
    LocalMux I__3545 (
            .O(N__30614),
            .I(\quad_counter1.B_delayed ));
    InMux I__3544 (
            .O(N__30609),
            .I(N__30603));
    InMux I__3543 (
            .O(N__30608),
            .I(N__30603));
    LocalMux I__3542 (
            .O(N__30603),
            .I(\c0.data_out_frame_29__7__N_849 ));
    SRMux I__3541 (
            .O(N__30600),
            .I(N__30597));
    LocalMux I__3540 (
            .O(N__30597),
            .I(\c0.n21597 ));
    SRMux I__3539 (
            .O(N__30594),
            .I(N__30591));
    LocalMux I__3538 (
            .O(N__30591),
            .I(N__30588));
    Odrv4 I__3537 (
            .O(N__30588),
            .I(\c0.n21587 ));
    CascadeMux I__3536 (
            .O(N__30585),
            .I(\c0.n10_adj_4303_cascade_ ));
    CascadeMux I__3535 (
            .O(N__30582),
            .I(N__30578));
    InMux I__3534 (
            .O(N__30581),
            .I(N__30574));
    InMux I__3533 (
            .O(N__30578),
            .I(N__30569));
    InMux I__3532 (
            .O(N__30577),
            .I(N__30569));
    LocalMux I__3531 (
            .O(N__30574),
            .I(N__30566));
    LocalMux I__3530 (
            .O(N__30569),
            .I(N__30562));
    Span4Mux_h I__3529 (
            .O(N__30566),
            .I(N__30559));
    InMux I__3528 (
            .O(N__30565),
            .I(N__30556));
    Span12Mux_v I__3527 (
            .O(N__30562),
            .I(N__30551));
    Span4Mux_v I__3526 (
            .O(N__30559),
            .I(N__30548));
    LocalMux I__3525 (
            .O(N__30556),
            .I(N__30545));
    InMux I__3524 (
            .O(N__30555),
            .I(N__30542));
    InMux I__3523 (
            .O(N__30554),
            .I(N__30539));
    Odrv12 I__3522 (
            .O(N__30551),
            .I(\c0.r_SM_Main_2_N_3754_0 ));
    Odrv4 I__3521 (
            .O(N__30548),
            .I(\c0.r_SM_Main_2_N_3754_0 ));
    Odrv4 I__3520 (
            .O(N__30545),
            .I(\c0.r_SM_Main_2_N_3754_0 ));
    LocalMux I__3519 (
            .O(N__30542),
            .I(\c0.r_SM_Main_2_N_3754_0 ));
    LocalMux I__3518 (
            .O(N__30539),
            .I(\c0.r_SM_Main_2_N_3754_0 ));
    InMux I__3517 (
            .O(N__30528),
            .I(N__30521));
    InMux I__3516 (
            .O(N__30527),
            .I(N__30521));
    InMux I__3515 (
            .O(N__30526),
            .I(N__30517));
    LocalMux I__3514 (
            .O(N__30521),
            .I(N__30514));
    InMux I__3513 (
            .O(N__30520),
            .I(N__30511));
    LocalMux I__3512 (
            .O(N__30517),
            .I(N__30508));
    Span4Mux_v I__3511 (
            .O(N__30514),
            .I(N__30505));
    LocalMux I__3510 (
            .O(N__30511),
            .I(\c0.tx_active ));
    Odrv4 I__3509 (
            .O(N__30508),
            .I(\c0.tx_active ));
    Odrv4 I__3508 (
            .O(N__30505),
            .I(\c0.tx_active ));
    CascadeMux I__3507 (
            .O(N__30498),
            .I(\c0.n5_cascade_ ));
    SRMux I__3506 (
            .O(N__30495),
            .I(N__30492));
    LocalMux I__3505 (
            .O(N__30492),
            .I(N__30489));
    Span4Mux_h I__3504 (
            .O(N__30489),
            .I(N__30486));
    Odrv4 I__3503 (
            .O(N__30486),
            .I(\c0.n21585 ));
    InMux I__3502 (
            .O(N__30483),
            .I(N__30480));
    LocalMux I__3501 (
            .O(N__30480),
            .I(\c0.n3 ));
    CascadeMux I__3500 (
            .O(N__30477),
            .I(\c0.n8_adj_4740_cascade_ ));
    CascadeMux I__3499 (
            .O(N__30474),
            .I(\c0.n22952_cascade_ ));
    CEMux I__3498 (
            .O(N__30471),
            .I(N__30468));
    LocalMux I__3497 (
            .O(N__30468),
            .I(\c0.n14380 ));
    CascadeMux I__3496 (
            .O(N__30465),
            .I(\c0.n14380_cascade_ ));
    SRMux I__3495 (
            .O(N__30462),
            .I(N__30459));
    LocalMux I__3494 (
            .O(N__30459),
            .I(\c0.n14942 ));
    InMux I__3493 (
            .O(N__30456),
            .I(N__30453));
    LocalMux I__3492 (
            .O(N__30453),
            .I(\c0.n4728 ));
    CascadeMux I__3491 (
            .O(N__30450),
            .I(\c0.n4728_cascade_ ));
    InMux I__3490 (
            .O(N__30447),
            .I(N__30444));
    LocalMux I__3489 (
            .O(N__30444),
            .I(\c0.n58_adj_4742 ));
    SRMux I__3488 (
            .O(N__30441),
            .I(N__30438));
    LocalMux I__3487 (
            .O(N__30438),
            .I(N__30434));
    InMux I__3486 (
            .O(N__30437),
            .I(N__30431));
    Odrv4 I__3485 (
            .O(N__30434),
            .I(\c0.n22952 ));
    LocalMux I__3484 (
            .O(N__30431),
            .I(\c0.n22952 ));
    InMux I__3483 (
            .O(N__30426),
            .I(N__30423));
    LocalMux I__3482 (
            .O(N__30423),
            .I(n25008));
    InMux I__3481 (
            .O(N__30420),
            .I(N__30417));
    LocalMux I__3480 (
            .O(N__30417),
            .I(\c0.n11_adj_4681 ));
    InMux I__3479 (
            .O(N__30414),
            .I(N__30411));
    LocalMux I__3478 (
            .O(N__30411),
            .I(N__30408));
    Odrv4 I__3477 (
            .O(N__30408),
            .I(\c0.n24897 ));
    InMux I__3476 (
            .O(N__30405),
            .I(N__30399));
    InMux I__3475 (
            .O(N__30404),
            .I(N__30399));
    LocalMux I__3474 (
            .O(N__30399),
            .I(data_out_frame_5_0));
    InMux I__3473 (
            .O(N__30396),
            .I(N__30390));
    InMux I__3472 (
            .O(N__30395),
            .I(N__30390));
    LocalMux I__3471 (
            .O(N__30390),
            .I(data_out_frame_0_2));
    InMux I__3470 (
            .O(N__30387),
            .I(N__30383));
    InMux I__3469 (
            .O(N__30386),
            .I(N__30380));
    LocalMux I__3468 (
            .O(N__30383),
            .I(N__30377));
    LocalMux I__3467 (
            .O(N__30380),
            .I(data_out_frame_12_5));
    Odrv4 I__3466 (
            .O(N__30377),
            .I(data_out_frame_12_5));
    InMux I__3465 (
            .O(N__30372),
            .I(N__30369));
    LocalMux I__3464 (
            .O(N__30369),
            .I(N__30366));
    Odrv12 I__3463 (
            .O(N__30366),
            .I(\c0.n24900 ));
    CascadeMux I__3462 (
            .O(N__30363),
            .I(n14247_cascade_));
    InMux I__3461 (
            .O(N__30360),
            .I(N__30354));
    InMux I__3460 (
            .O(N__30359),
            .I(N__30354));
    LocalMux I__3459 (
            .O(N__30354),
            .I(data_out_frame_0_3));
    InMux I__3458 (
            .O(N__30351),
            .I(N__30348));
    LocalMux I__3457 (
            .O(N__30348),
            .I(N__30345));
    Span4Mux_v I__3456 (
            .O(N__30345),
            .I(N__30342));
    Odrv4 I__3455 (
            .O(N__30342),
            .I(n24796));
    InMux I__3454 (
            .O(N__30339),
            .I(N__30336));
    LocalMux I__3453 (
            .O(N__30336),
            .I(N__30332));
    InMux I__3452 (
            .O(N__30335),
            .I(N__30329));
    Span4Mux_h I__3451 (
            .O(N__30332),
            .I(N__30326));
    LocalMux I__3450 (
            .O(N__30329),
            .I(data_out_frame_7_7));
    Odrv4 I__3449 (
            .O(N__30326),
            .I(data_out_frame_7_7));
    CascadeMux I__3448 (
            .O(N__30321),
            .I(n24805_cascade_));
    InMux I__3447 (
            .O(N__30318),
            .I(N__30315));
    LocalMux I__3446 (
            .O(N__30315),
            .I(n10_adj_4780));
    CascadeMux I__3445 (
            .O(N__30312),
            .I(N__30309));
    InMux I__3444 (
            .O(N__30309),
            .I(N__30305));
    InMux I__3443 (
            .O(N__30308),
            .I(N__30302));
    LocalMux I__3442 (
            .O(N__30305),
            .I(N__30299));
    LocalMux I__3441 (
            .O(N__30302),
            .I(data_out_frame_11_5));
    Odrv4 I__3440 (
            .O(N__30299),
            .I(data_out_frame_11_5));
    CascadeMux I__3439 (
            .O(N__30294),
            .I(\c0.n25092_cascade_ ));
    CascadeMux I__3438 (
            .O(N__30291),
            .I(\c0.n25095_cascade_ ));
    CascadeMux I__3437 (
            .O(N__30288),
            .I(N__30285));
    InMux I__3436 (
            .O(N__30285),
            .I(N__30282));
    LocalMux I__3435 (
            .O(N__30282),
            .I(N__30279));
    Span4Mux_v I__3434 (
            .O(N__30279),
            .I(N__30276));
    Odrv4 I__3433 (
            .O(N__30276),
            .I(n25014));
    CascadeMux I__3432 (
            .O(N__30273),
            .I(N__30270));
    InMux I__3431 (
            .O(N__30270),
            .I(N__30264));
    InMux I__3430 (
            .O(N__30269),
            .I(N__30264));
    LocalMux I__3429 (
            .O(N__30264),
            .I(data_out_frame_9_5));
    CascadeMux I__3428 (
            .O(N__30261),
            .I(\c0.n20341_cascade_ ));
    InMux I__3427 (
            .O(N__30258),
            .I(N__30255));
    LocalMux I__3426 (
            .O(N__30255),
            .I(N__30251));
    InMux I__3425 (
            .O(N__30254),
            .I(N__30248));
    Span4Mux_v I__3424 (
            .O(N__30251),
            .I(N__30245));
    LocalMux I__3423 (
            .O(N__30248),
            .I(data_out_frame_13_7));
    Odrv4 I__3422 (
            .O(N__30245),
            .I(data_out_frame_13_7));
    InMux I__3421 (
            .O(N__30240),
            .I(N__30237));
    LocalMux I__3420 (
            .O(N__30237),
            .I(N__30233));
    InMux I__3419 (
            .O(N__30236),
            .I(N__30230));
    Span4Mux_v I__3418 (
            .O(N__30233),
            .I(N__30227));
    LocalMux I__3417 (
            .O(N__30230),
            .I(data_out_frame_10_7));
    Odrv4 I__3416 (
            .O(N__30227),
            .I(data_out_frame_10_7));
    CascadeMux I__3415 (
            .O(N__30222),
            .I(N__30218));
    CascadeMux I__3414 (
            .O(N__30221),
            .I(N__30214));
    InMux I__3413 (
            .O(N__30218),
            .I(N__30210));
    InMux I__3412 (
            .O(N__30217),
            .I(N__30207));
    InMux I__3411 (
            .O(N__30214),
            .I(N__30204));
    InMux I__3410 (
            .O(N__30213),
            .I(N__30198));
    LocalMux I__3409 (
            .O(N__30210),
            .I(N__30195));
    LocalMux I__3408 (
            .O(N__30207),
            .I(N__30192));
    LocalMux I__3407 (
            .O(N__30204),
            .I(N__30189));
    InMux I__3406 (
            .O(N__30203),
            .I(N__30184));
    InMux I__3405 (
            .O(N__30202),
            .I(N__30184));
    InMux I__3404 (
            .O(N__30201),
            .I(N__30181));
    LocalMux I__3403 (
            .O(N__30198),
            .I(N__30178));
    Span4Mux_h I__3402 (
            .O(N__30195),
            .I(N__30175));
    Span4Mux_v I__3401 (
            .O(N__30192),
            .I(N__30168));
    Span4Mux_h I__3400 (
            .O(N__30189),
            .I(N__30168));
    LocalMux I__3399 (
            .O(N__30184),
            .I(N__30168));
    LocalMux I__3398 (
            .O(N__30181),
            .I(N__30165));
    Span4Mux_h I__3397 (
            .O(N__30178),
            .I(N__30162));
    Span4Mux_v I__3396 (
            .O(N__30175),
            .I(N__30159));
    Span4Mux_v I__3395 (
            .O(N__30168),
            .I(N__30156));
    Odrv12 I__3394 (
            .O(N__30165),
            .I(n9603));
    Odrv4 I__3393 (
            .O(N__30162),
            .I(n9603));
    Odrv4 I__3392 (
            .O(N__30159),
            .I(n9603));
    Odrv4 I__3391 (
            .O(N__30156),
            .I(n9603));
    CascadeMux I__3390 (
            .O(N__30147),
            .I(N__30143));
    CascadeMux I__3389 (
            .O(N__30146),
            .I(N__30140));
    InMux I__3388 (
            .O(N__30143),
            .I(N__30135));
    InMux I__3387 (
            .O(N__30140),
            .I(N__30132));
    InMux I__3386 (
            .O(N__30139),
            .I(N__30126));
    CascadeMux I__3385 (
            .O(N__30138),
            .I(N__30122));
    LocalMux I__3384 (
            .O(N__30135),
            .I(N__30119));
    LocalMux I__3383 (
            .O(N__30132),
            .I(N__30116));
    InMux I__3382 (
            .O(N__30131),
            .I(N__30113));
    CascadeMux I__3381 (
            .O(N__30130),
            .I(N__30110));
    InMux I__3380 (
            .O(N__30129),
            .I(N__30107));
    LocalMux I__3379 (
            .O(N__30126),
            .I(N__30104));
    InMux I__3378 (
            .O(N__30125),
            .I(N__30099));
    InMux I__3377 (
            .O(N__30122),
            .I(N__30099));
    Span4Mux_h I__3376 (
            .O(N__30119),
            .I(N__30096));
    Span4Mux_v I__3375 (
            .O(N__30116),
            .I(N__30091));
    LocalMux I__3374 (
            .O(N__30113),
            .I(N__30091));
    InMux I__3373 (
            .O(N__30110),
            .I(N__30087));
    LocalMux I__3372 (
            .O(N__30107),
            .I(N__30084));
    Span4Mux_h I__3371 (
            .O(N__30104),
            .I(N__30081));
    LocalMux I__3370 (
            .O(N__30099),
            .I(N__30078));
    Sp12to4 I__3369 (
            .O(N__30096),
            .I(N__30073));
    Sp12to4 I__3368 (
            .O(N__30091),
            .I(N__30073));
    InMux I__3367 (
            .O(N__30090),
            .I(N__30069));
    LocalMux I__3366 (
            .O(N__30087),
            .I(N__30064));
    Span4Mux_h I__3365 (
            .O(N__30084),
            .I(N__30064));
    Span4Mux_v I__3364 (
            .O(N__30081),
            .I(N__30061));
    Span12Mux_v I__3363 (
            .O(N__30078),
            .I(N__30058));
    Span12Mux_v I__3362 (
            .O(N__30073),
            .I(N__30055));
    InMux I__3361 (
            .O(N__30072),
            .I(N__30052));
    LocalMux I__3360 (
            .O(N__30069),
            .I(byte_transmit_counter_5));
    Odrv4 I__3359 (
            .O(N__30064),
            .I(byte_transmit_counter_5));
    Odrv4 I__3358 (
            .O(N__30061),
            .I(byte_transmit_counter_5));
    Odrv12 I__3357 (
            .O(N__30058),
            .I(byte_transmit_counter_5));
    Odrv12 I__3356 (
            .O(N__30055),
            .I(byte_transmit_counter_5));
    LocalMux I__3355 (
            .O(N__30052),
            .I(byte_transmit_counter_5));
    CascadeMux I__3354 (
            .O(N__30039),
            .I(N__30036));
    InMux I__3353 (
            .O(N__30036),
            .I(N__30033));
    LocalMux I__3352 (
            .O(N__30033),
            .I(N__30029));
    InMux I__3351 (
            .O(N__30032),
            .I(N__30026));
    Span4Mux_h I__3350 (
            .O(N__30029),
            .I(N__30023));
    LocalMux I__3349 (
            .O(N__30026),
            .I(r_Tx_Data_0));
    Odrv4 I__3348 (
            .O(N__30023),
            .I(r_Tx_Data_0));
    InMux I__3347 (
            .O(N__30018),
            .I(N__30014));
    InMux I__3346 (
            .O(N__30017),
            .I(N__30011));
    LocalMux I__3345 (
            .O(N__30014),
            .I(N__30008));
    LocalMux I__3344 (
            .O(N__30011),
            .I(data_out_frame_13_6));
    Odrv4 I__3343 (
            .O(N__30008),
            .I(data_out_frame_13_6));
    InMux I__3342 (
            .O(N__30003),
            .I(N__30000));
    LocalMux I__3341 (
            .O(N__30000),
            .I(N__29996));
    InMux I__3340 (
            .O(N__29999),
            .I(N__29993));
    Span4Mux_h I__3339 (
            .O(N__29996),
            .I(N__29990));
    LocalMux I__3338 (
            .O(N__29993),
            .I(data_out_frame_8_3));
    Odrv4 I__3337 (
            .O(N__29990),
            .I(data_out_frame_8_3));
    CascadeMux I__3336 (
            .O(N__29985),
            .I(\c0.n24033_cascade_ ));
    CascadeMux I__3335 (
            .O(N__29982),
            .I(n21307_cascade_));
    CascadeMux I__3334 (
            .O(N__29979),
            .I(\c0.n7_cascade_ ));
    InMux I__3333 (
            .O(N__29976),
            .I(N__29973));
    LocalMux I__3332 (
            .O(N__29973),
            .I(\c0.n23918 ));
    InMux I__3331 (
            .O(N__29970),
            .I(N__29967));
    LocalMux I__3330 (
            .O(N__29967),
            .I(N__29963));
    InMux I__3329 (
            .O(N__29966),
            .I(N__29960));
    Span4Mux_v I__3328 (
            .O(N__29963),
            .I(N__29957));
    LocalMux I__3327 (
            .O(N__29960),
            .I(r_Tx_Data_2));
    Odrv4 I__3326 (
            .O(N__29957),
            .I(r_Tx_Data_2));
    InMux I__3325 (
            .O(N__29952),
            .I(N__29949));
    LocalMux I__3324 (
            .O(N__29949),
            .I(\c0.n22163 ));
    CascadeMux I__3323 (
            .O(N__29946),
            .I(\c0.n6_adj_4297_cascade_ ));
    InMux I__3322 (
            .O(N__29943),
            .I(N__29940));
    LocalMux I__3321 (
            .O(N__29940),
            .I(\c0.data_out_frame_28_4 ));
    CascadeMux I__3320 (
            .O(N__29937),
            .I(n26_cascade_));
    InMux I__3319 (
            .O(N__29934),
            .I(N__29931));
    LocalMux I__3318 (
            .O(N__29931),
            .I(N__29928));
    Odrv4 I__3317 (
            .O(N__29928),
            .I(n25021));
    InMux I__3316 (
            .O(N__29925),
            .I(N__29922));
    LocalMux I__3315 (
            .O(N__29922),
            .I(N__29919));
    Odrv4 I__3314 (
            .O(N__29919),
            .I(n25022));
    CascadeMux I__3313 (
            .O(N__29916),
            .I(\c0.n21391_cascade_ ));
    CascadeMux I__3312 (
            .O(N__29913),
            .I(\c0.n21362_cascade_ ));
    CascadeMux I__3311 (
            .O(N__29910),
            .I(\c0.n21244_cascade_ ));
    CascadeMux I__3310 (
            .O(N__29907),
            .I(N__29903));
    InMux I__3309 (
            .O(N__29906),
            .I(N__29900));
    InMux I__3308 (
            .O(N__29903),
            .I(N__29897));
    LocalMux I__3307 (
            .O(N__29900),
            .I(N__29892));
    LocalMux I__3306 (
            .O(N__29897),
            .I(N__29892));
    Span4Mux_h I__3305 (
            .O(N__29892),
            .I(N__29888));
    InMux I__3304 (
            .O(N__29891),
            .I(N__29885));
    Span4Mux_h I__3303 (
            .O(N__29888),
            .I(N__29882));
    LocalMux I__3302 (
            .O(N__29885),
            .I(B_filtered_adj_4764));
    Odrv4 I__3301 (
            .O(N__29882),
            .I(B_filtered_adj_4764));
    InMux I__3300 (
            .O(N__29877),
            .I(N__29874));
    LocalMux I__3299 (
            .O(N__29874),
            .I(\quad_counter1.A_delayed ));
    CascadeMux I__3298 (
            .O(N__29871),
            .I(N__29867));
    InMux I__3297 (
            .O(N__29870),
            .I(N__29864));
    InMux I__3296 (
            .O(N__29867),
            .I(N__29861));
    LocalMux I__3295 (
            .O(N__29864),
            .I(r_Tx_Data_4));
    LocalMux I__3294 (
            .O(N__29861),
            .I(r_Tx_Data_4));
    CascadeMux I__3293 (
            .O(N__29856),
            .I(n9806_cascade_));
    InMux I__3292 (
            .O(N__29853),
            .I(N__29847));
    InMux I__3291 (
            .O(N__29852),
            .I(N__29847));
    LocalMux I__3290 (
            .O(N__29847),
            .I(N__29842));
    InMux I__3289 (
            .O(N__29846),
            .I(N__29837));
    InMux I__3288 (
            .O(N__29845),
            .I(N__29837));
    Span4Mux_h I__3287 (
            .O(N__29842),
            .I(N__29834));
    LocalMux I__3286 (
            .O(N__29837),
            .I(N__29831));
    Span4Mux_h I__3285 (
            .O(N__29834),
            .I(N__29828));
    Span12Mux_h I__3284 (
            .O(N__29831),
            .I(N__29825));
    Span4Mux_v I__3283 (
            .O(N__29828),
            .I(N__29822));
    Odrv12 I__3282 (
            .O(N__29825),
            .I(PIN_12_c));
    Odrv4 I__3281 (
            .O(N__29822),
            .I(PIN_12_c));
    InMux I__3280 (
            .O(N__29817),
            .I(N__29810));
    InMux I__3279 (
            .O(N__29816),
            .I(N__29810));
    InMux I__3278 (
            .O(N__29815),
            .I(N__29807));
    LocalMux I__3277 (
            .O(N__29810),
            .I(quadA_delayed_adj_4767));
    LocalMux I__3276 (
            .O(N__29807),
            .I(quadA_delayed_adj_4767));
    InMux I__3275 (
            .O(N__29802),
            .I(N__29799));
    LocalMux I__3274 (
            .O(N__29799),
            .I(n9806));
    CEMux I__3273 (
            .O(N__29796),
            .I(N__29793));
    LocalMux I__3272 (
            .O(N__29793),
            .I(N__29790));
    Span4Mux_h I__3271 (
            .O(N__29790),
            .I(N__29786));
    CEMux I__3270 (
            .O(N__29789),
            .I(N__29783));
    Odrv4 I__3269 (
            .O(N__29786),
            .I(n14345));
    LocalMux I__3268 (
            .O(N__29783),
            .I(n14345));
    SRMux I__3267 (
            .O(N__29778),
            .I(N__29774));
    SRMux I__3266 (
            .O(N__29777),
            .I(N__29771));
    LocalMux I__3265 (
            .O(N__29774),
            .I(N__29767));
    LocalMux I__3264 (
            .O(N__29771),
            .I(N__29764));
    InMux I__3263 (
            .O(N__29770),
            .I(N__29761));
    Span4Mux_h I__3262 (
            .O(N__29767),
            .I(N__29758));
    Span4Mux_h I__3261 (
            .O(N__29764),
            .I(N__29755));
    LocalMux I__3260 (
            .O(N__29761),
            .I(a_delay_counter_15__N_4123_adj_4772));
    Odrv4 I__3259 (
            .O(N__29758),
            .I(a_delay_counter_15__N_4123_adj_4772));
    Odrv4 I__3258 (
            .O(N__29755),
            .I(a_delay_counter_15__N_4123_adj_4772));
    CascadeMux I__3257 (
            .O(N__29748),
            .I(n14345_cascade_));
    InMux I__3256 (
            .O(N__29745),
            .I(N__29742));
    LocalMux I__3255 (
            .O(N__29742),
            .I(n39_adj_4770));
    InMux I__3254 (
            .O(N__29739),
            .I(N__29735));
    InMux I__3253 (
            .O(N__29738),
            .I(N__29732));
    LocalMux I__3252 (
            .O(N__29735),
            .I(\quad_counter1.a_delay_counter_5 ));
    LocalMux I__3251 (
            .O(N__29732),
            .I(\quad_counter1.a_delay_counter_5 ));
    InMux I__3250 (
            .O(N__29727),
            .I(N__29723));
    InMux I__3249 (
            .O(N__29726),
            .I(N__29720));
    LocalMux I__3248 (
            .O(N__29723),
            .I(\quad_counter1.a_delay_counter_11 ));
    LocalMux I__3247 (
            .O(N__29720),
            .I(\quad_counter1.a_delay_counter_11 ));
    CascadeMux I__3246 (
            .O(N__29715),
            .I(N__29711));
    InMux I__3245 (
            .O(N__29714),
            .I(N__29708));
    InMux I__3244 (
            .O(N__29711),
            .I(N__29705));
    LocalMux I__3243 (
            .O(N__29708),
            .I(\quad_counter1.a_delay_counter_4 ));
    LocalMux I__3242 (
            .O(N__29705),
            .I(\quad_counter1.a_delay_counter_4 ));
    InMux I__3241 (
            .O(N__29700),
            .I(N__29695));
    InMux I__3240 (
            .O(N__29699),
            .I(N__29690));
    InMux I__3239 (
            .O(N__29698),
            .I(N__29690));
    LocalMux I__3238 (
            .O(N__29695),
            .I(a_delay_counter_0_adj_4765));
    LocalMux I__3237 (
            .O(N__29690),
            .I(a_delay_counter_0_adj_4765));
    CascadeMux I__3236 (
            .O(N__29685),
            .I(N__29682));
    InMux I__3235 (
            .O(N__29682),
            .I(N__29679));
    LocalMux I__3234 (
            .O(N__29679),
            .I(\quad_counter1.n25 ));
    InMux I__3233 (
            .O(N__29676),
            .I(N__29672));
    InMux I__3232 (
            .O(N__29675),
            .I(N__29669));
    LocalMux I__3231 (
            .O(N__29672),
            .I(\quad_counter1.a_delay_counter_9 ));
    LocalMux I__3230 (
            .O(N__29669),
            .I(\quad_counter1.a_delay_counter_9 ));
    InMux I__3229 (
            .O(N__29664),
            .I(N__29660));
    InMux I__3228 (
            .O(N__29663),
            .I(N__29657));
    LocalMux I__3227 (
            .O(N__29660),
            .I(\quad_counter1.a_delay_counter_6 ));
    LocalMux I__3226 (
            .O(N__29657),
            .I(\quad_counter1.a_delay_counter_6 ));
    CascadeMux I__3225 (
            .O(N__29652),
            .I(N__29648));
    InMux I__3224 (
            .O(N__29651),
            .I(N__29645));
    InMux I__3223 (
            .O(N__29648),
            .I(N__29642));
    LocalMux I__3222 (
            .O(N__29645),
            .I(\quad_counter1.a_delay_counter_12 ));
    LocalMux I__3221 (
            .O(N__29642),
            .I(\quad_counter1.a_delay_counter_12 ));
    InMux I__3220 (
            .O(N__29637),
            .I(N__29633));
    InMux I__3219 (
            .O(N__29636),
            .I(N__29630));
    LocalMux I__3218 (
            .O(N__29633),
            .I(\quad_counter1.a_delay_counter_13 ));
    LocalMux I__3217 (
            .O(N__29630),
            .I(\quad_counter1.a_delay_counter_13 ));
    InMux I__3216 (
            .O(N__29625),
            .I(N__29622));
    LocalMux I__3215 (
            .O(N__29622),
            .I(\quad_counter1.n26 ));
    InMux I__3214 (
            .O(N__29619),
            .I(N__29615));
    InMux I__3213 (
            .O(N__29618),
            .I(N__29612));
    LocalMux I__3212 (
            .O(N__29615),
            .I(\quad_counter1.a_delay_counter_8 ));
    LocalMux I__3211 (
            .O(N__29612),
            .I(\quad_counter1.a_delay_counter_8 ));
    InMux I__3210 (
            .O(N__29607),
            .I(N__29603));
    InMux I__3209 (
            .O(N__29606),
            .I(N__29600));
    LocalMux I__3208 (
            .O(N__29603),
            .I(\quad_counter1.a_delay_counter_1 ));
    LocalMux I__3207 (
            .O(N__29600),
            .I(\quad_counter1.a_delay_counter_1 ));
    CascadeMux I__3206 (
            .O(N__29595),
            .I(N__29591));
    InMux I__3205 (
            .O(N__29594),
            .I(N__29588));
    InMux I__3204 (
            .O(N__29591),
            .I(N__29585));
    LocalMux I__3203 (
            .O(N__29588),
            .I(\quad_counter1.a_delay_counter_2 ));
    LocalMux I__3202 (
            .O(N__29585),
            .I(\quad_counter1.a_delay_counter_2 ));
    InMux I__3201 (
            .O(N__29580),
            .I(N__29576));
    InMux I__3200 (
            .O(N__29579),
            .I(N__29573));
    LocalMux I__3199 (
            .O(N__29576),
            .I(\quad_counter1.a_delay_counter_3 ));
    LocalMux I__3198 (
            .O(N__29573),
            .I(\quad_counter1.a_delay_counter_3 ));
    InMux I__3197 (
            .O(N__29568),
            .I(N__29565));
    LocalMux I__3196 (
            .O(N__29565),
            .I(\quad_counter1.n28 ));
    InMux I__3195 (
            .O(N__29562),
            .I(N__29558));
    InMux I__3194 (
            .O(N__29561),
            .I(N__29555));
    LocalMux I__3193 (
            .O(N__29558),
            .I(\quad_counter1.a_delay_counter_14 ));
    LocalMux I__3192 (
            .O(N__29555),
            .I(\quad_counter1.a_delay_counter_14 ));
    InMux I__3191 (
            .O(N__29550),
            .I(N__29546));
    InMux I__3190 (
            .O(N__29549),
            .I(N__29543));
    LocalMux I__3189 (
            .O(N__29546),
            .I(\quad_counter1.a_delay_counter_7 ));
    LocalMux I__3188 (
            .O(N__29543),
            .I(\quad_counter1.a_delay_counter_7 ));
    CascadeMux I__3187 (
            .O(N__29538),
            .I(N__29534));
    InMux I__3186 (
            .O(N__29537),
            .I(N__29531));
    InMux I__3185 (
            .O(N__29534),
            .I(N__29528));
    LocalMux I__3184 (
            .O(N__29531),
            .I(\quad_counter1.a_delay_counter_10 ));
    LocalMux I__3183 (
            .O(N__29528),
            .I(\quad_counter1.a_delay_counter_10 ));
    InMux I__3182 (
            .O(N__29523),
            .I(N__29519));
    InMux I__3181 (
            .O(N__29522),
            .I(N__29516));
    LocalMux I__3180 (
            .O(N__29519),
            .I(\quad_counter1.a_delay_counter_15 ));
    LocalMux I__3179 (
            .O(N__29516),
            .I(\quad_counter1.a_delay_counter_15 ));
    InMux I__3178 (
            .O(N__29511),
            .I(N__29508));
    LocalMux I__3177 (
            .O(N__29508),
            .I(\quad_counter1.n27 ));
    CascadeMux I__3176 (
            .O(N__29505),
            .I(N__29502));
    InMux I__3175 (
            .O(N__29502),
            .I(N__29498));
    InMux I__3174 (
            .O(N__29501),
            .I(N__29495));
    LocalMux I__3173 (
            .O(N__29498),
            .I(N__29491));
    LocalMux I__3172 (
            .O(N__29495),
            .I(N__29488));
    InMux I__3171 (
            .O(N__29494),
            .I(N__29485));
    Span12Mux_v I__3170 (
            .O(N__29491),
            .I(N__29482));
    Span4Mux_h I__3169 (
            .O(N__29488),
            .I(N__29479));
    LocalMux I__3168 (
            .O(N__29485),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv12 I__3167 (
            .O(N__29482),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv4 I__3166 (
            .O(N__29479),
            .I(\c0.FRAME_MATCHER_state_13 ));
    SRMux I__3165 (
            .O(N__29472),
            .I(N__29469));
    LocalMux I__3164 (
            .O(N__29469),
            .I(N__29466));
    Span4Mux_h I__3163 (
            .O(N__29466),
            .I(N__29463));
    Span4Mux_v I__3162 (
            .O(N__29463),
            .I(N__29460));
    Odrv4 I__3161 (
            .O(N__29460),
            .I(\c0.n21573 ));
    SRMux I__3160 (
            .O(N__29457),
            .I(N__29454));
    LocalMux I__3159 (
            .O(N__29454),
            .I(N__29451));
    Span4Mux_h I__3158 (
            .O(N__29451),
            .I(N__29448));
    Odrv4 I__3157 (
            .O(N__29448),
            .I(\c0.n21581 ));
    SRMux I__3156 (
            .O(N__29445),
            .I(N__29442));
    LocalMux I__3155 (
            .O(N__29442),
            .I(N__29439));
    Span4Mux_h I__3154 (
            .O(N__29439),
            .I(N__29436));
    Odrv4 I__3153 (
            .O(N__29436),
            .I(\c0.n21575 ));
    CascadeMux I__3152 (
            .O(N__29433),
            .I(N__29430));
    InMux I__3151 (
            .O(N__29430),
            .I(N__29426));
    CascadeMux I__3150 (
            .O(N__29429),
            .I(N__29423));
    LocalMux I__3149 (
            .O(N__29426),
            .I(N__29420));
    InMux I__3148 (
            .O(N__29423),
            .I(N__29416));
    Span4Mux_v I__3147 (
            .O(N__29420),
            .I(N__29413));
    InMux I__3146 (
            .O(N__29419),
            .I(N__29410));
    LocalMux I__3145 (
            .O(N__29416),
            .I(N__29405));
    Span4Mux_v I__3144 (
            .O(N__29413),
            .I(N__29405));
    LocalMux I__3143 (
            .O(N__29410),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__3142 (
            .O(N__29405),
            .I(\c0.FRAME_MATCHER_state_14 ));
    SRMux I__3141 (
            .O(N__29400),
            .I(N__29397));
    LocalMux I__3140 (
            .O(N__29397),
            .I(N__29394));
    Span4Mux_h I__3139 (
            .O(N__29394),
            .I(N__29391));
    Odrv4 I__3138 (
            .O(N__29391),
            .I(\c0.n21577 ));
    InMux I__3137 (
            .O(N__29388),
            .I(\c0.n19796 ));
    InMux I__3136 (
            .O(N__29385),
            .I(\c0.n19797 ));
    InMux I__3135 (
            .O(N__29382),
            .I(\c0.n19798 ));
    InMux I__3134 (
            .O(N__29379),
            .I(\c0.n19799 ));
    InMux I__3133 (
            .O(N__29376),
            .I(N__29372));
    InMux I__3132 (
            .O(N__29375),
            .I(N__29369));
    LocalMux I__3131 (
            .O(N__29372),
            .I(\c0.byte_transmit_counter_6 ));
    LocalMux I__3130 (
            .O(N__29369),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__3129 (
            .O(N__29364),
            .I(\c0.n19800 ));
    InMux I__3128 (
            .O(N__29361),
            .I(\c0.n19801 ));
    InMux I__3127 (
            .O(N__29358),
            .I(N__29354));
    InMux I__3126 (
            .O(N__29357),
            .I(N__29351));
    LocalMux I__3125 (
            .O(N__29354),
            .I(\c0.byte_transmit_counter_7 ));
    LocalMux I__3124 (
            .O(N__29351),
            .I(\c0.byte_transmit_counter_7 ));
    SRMux I__3123 (
            .O(N__29346),
            .I(N__29343));
    LocalMux I__3122 (
            .O(N__29343),
            .I(N__29340));
    Span4Mux_h I__3121 (
            .O(N__29340),
            .I(N__29337));
    Odrv4 I__3120 (
            .O(N__29337),
            .I(\c0.n21611 ));
    CascadeMux I__3119 (
            .O(N__29334),
            .I(N__29331));
    InMux I__3118 (
            .O(N__29331),
            .I(N__29327));
    InMux I__3117 (
            .O(N__29330),
            .I(N__29324));
    LocalMux I__3116 (
            .O(N__29327),
            .I(data_out_frame_12_6));
    LocalMux I__3115 (
            .O(N__29324),
            .I(data_out_frame_12_6));
    InMux I__3114 (
            .O(N__29319),
            .I(N__29316));
    LocalMux I__3113 (
            .O(N__29316),
            .I(\c0.n5_adj_4334 ));
    InMux I__3112 (
            .O(N__29313),
            .I(N__29310));
    LocalMux I__3111 (
            .O(N__29310),
            .I(\c0.n4_adj_4332 ));
    InMux I__3110 (
            .O(N__29307),
            .I(N__29304));
    LocalMux I__3109 (
            .O(N__29304),
            .I(N__29301));
    Span4Mux_v I__3108 (
            .O(N__29301),
            .I(N__29298));
    Odrv4 I__3107 (
            .O(N__29298),
            .I(\c0.n26_adj_4662 ));
    InMux I__3106 (
            .O(N__29295),
            .I(\c0.n19795 ));
    InMux I__3105 (
            .O(N__29292),
            .I(N__29288));
    InMux I__3104 (
            .O(N__29291),
            .I(N__29285));
    LocalMux I__3103 (
            .O(N__29288),
            .I(N__29282));
    LocalMux I__3102 (
            .O(N__29285),
            .I(r_Tx_Data_6));
    Odrv12 I__3101 (
            .O(N__29282),
            .I(r_Tx_Data_6));
    CascadeMux I__3100 (
            .O(N__29277),
            .I(N__29274));
    InMux I__3099 (
            .O(N__29274),
            .I(N__29270));
    InMux I__3098 (
            .O(N__29273),
            .I(N__29267));
    LocalMux I__3097 (
            .O(N__29270),
            .I(N__29264));
    LocalMux I__3096 (
            .O(N__29267),
            .I(data_out_frame_5_2));
    Odrv12 I__3095 (
            .O(N__29264),
            .I(data_out_frame_5_2));
    InMux I__3094 (
            .O(N__29259),
            .I(N__29253));
    InMux I__3093 (
            .O(N__29258),
            .I(N__29253));
    LocalMux I__3092 (
            .O(N__29253),
            .I(N__29250));
    Odrv4 I__3091 (
            .O(N__29250),
            .I(n17951));
    InMux I__3090 (
            .O(N__29247),
            .I(N__29232));
    InMux I__3089 (
            .O(N__29246),
            .I(N__29232));
    InMux I__3088 (
            .O(N__29245),
            .I(N__29232));
    InMux I__3087 (
            .O(N__29244),
            .I(N__29227));
    InMux I__3086 (
            .O(N__29243),
            .I(N__29227));
    InMux I__3085 (
            .O(N__29242),
            .I(N__29224));
    InMux I__3084 (
            .O(N__29241),
            .I(N__29221));
    InMux I__3083 (
            .O(N__29240),
            .I(N__29215));
    InMux I__3082 (
            .O(N__29239),
            .I(N__29215));
    LocalMux I__3081 (
            .O(N__29232),
            .I(N__29209));
    LocalMux I__3080 (
            .O(N__29227),
            .I(N__29206));
    LocalMux I__3079 (
            .O(N__29224),
            .I(N__29203));
    LocalMux I__3078 (
            .O(N__29221),
            .I(N__29200));
    InMux I__3077 (
            .O(N__29220),
            .I(N__29197));
    LocalMux I__3076 (
            .O(N__29215),
            .I(N__29194));
    InMux I__3075 (
            .O(N__29214),
            .I(N__29187));
    InMux I__3074 (
            .O(N__29213),
            .I(N__29187));
    InMux I__3073 (
            .O(N__29212),
            .I(N__29187));
    Span12Mux_s8_h I__3072 (
            .O(N__29209),
            .I(N__29180));
    Sp12to4 I__3071 (
            .O(N__29206),
            .I(N__29180));
    Span12Mux_s11_v I__3070 (
            .O(N__29203),
            .I(N__29180));
    Span4Mux_v I__3069 (
            .O(N__29200),
            .I(N__29175));
    LocalMux I__3068 (
            .O(N__29197),
            .I(N__29175));
    Span4Mux_h I__3067 (
            .O(N__29194),
            .I(N__29172));
    LocalMux I__3066 (
            .O(N__29187),
            .I(r_SM_Main_1_adj_4774));
    Odrv12 I__3065 (
            .O(N__29180),
            .I(r_SM_Main_1_adj_4774));
    Odrv4 I__3064 (
            .O(N__29175),
            .I(r_SM_Main_1_adj_4774));
    Odrv4 I__3063 (
            .O(N__29172),
            .I(r_SM_Main_1_adj_4774));
    InMux I__3062 (
            .O(N__29163),
            .I(N__29160));
    LocalMux I__3061 (
            .O(N__29160),
            .I(N__29157));
    Odrv12 I__3060 (
            .O(N__29157),
            .I(n25006));
    CascadeMux I__3059 (
            .O(N__29154),
            .I(N__29151));
    InMux I__3058 (
            .O(N__29151),
            .I(N__29148));
    LocalMux I__3057 (
            .O(N__29148),
            .I(N__29145));
    Span4Mux_h I__3056 (
            .O(N__29145),
            .I(N__29142));
    Odrv4 I__3055 (
            .O(N__29142),
            .I(\c0.n11_adj_4663 ));
    InMux I__3054 (
            .O(N__29139),
            .I(N__29136));
    LocalMux I__3053 (
            .O(N__29136),
            .I(N__29132));
    InMux I__3052 (
            .O(N__29135),
            .I(N__29129));
    Span4Mux_v I__3051 (
            .O(N__29132),
            .I(N__29126));
    LocalMux I__3050 (
            .O(N__29129),
            .I(data_out_frame_5_1));
    Odrv4 I__3049 (
            .O(N__29126),
            .I(data_out_frame_5_1));
    CascadeMux I__3048 (
            .O(N__29121),
            .I(N__29118));
    InMux I__3047 (
            .O(N__29118),
            .I(N__29112));
    InMux I__3046 (
            .O(N__29117),
            .I(N__29112));
    LocalMux I__3045 (
            .O(N__29112),
            .I(data_out_frame_13_3));
    InMux I__3044 (
            .O(N__29109),
            .I(N__29105));
    CascadeMux I__3043 (
            .O(N__29108),
            .I(N__29102));
    LocalMux I__3042 (
            .O(N__29105),
            .I(N__29099));
    InMux I__3041 (
            .O(N__29102),
            .I(N__29096));
    Span4Mux_h I__3040 (
            .O(N__29099),
            .I(N__29093));
    LocalMux I__3039 (
            .O(N__29096),
            .I(data_out_frame_8_7));
    Odrv4 I__3038 (
            .O(N__29093),
            .I(data_out_frame_8_7));
    CascadeMux I__3037 (
            .O(N__29088),
            .I(N__29085));
    InMux I__3036 (
            .O(N__29085),
            .I(N__29081));
    InMux I__3035 (
            .O(N__29084),
            .I(N__29078));
    LocalMux I__3034 (
            .O(N__29081),
            .I(N__29075));
    LocalMux I__3033 (
            .O(N__29078),
            .I(\c0.tx.r_Clock_Count_3 ));
    Odrv12 I__3032 (
            .O(N__29075),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__3031 (
            .O(N__29070),
            .I(\c0.tx.n19725 ));
    InMux I__3030 (
            .O(N__29067),
            .I(N__29063));
    InMux I__3029 (
            .O(N__29066),
            .I(N__29060));
    LocalMux I__3028 (
            .O(N__29063),
            .I(\c0.tx.r_Clock_Count_4 ));
    LocalMux I__3027 (
            .O(N__29060),
            .I(\c0.tx.r_Clock_Count_4 ));
    InMux I__3026 (
            .O(N__29055),
            .I(\c0.tx.n19726 ));
    InMux I__3025 (
            .O(N__29052),
            .I(N__29048));
    InMux I__3024 (
            .O(N__29051),
            .I(N__29045));
    LocalMux I__3023 (
            .O(N__29048),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__3022 (
            .O(N__29045),
            .I(\c0.tx.r_Clock_Count_5 ));
    InMux I__3021 (
            .O(N__29040),
            .I(\c0.tx.n19727 ));
    InMux I__3020 (
            .O(N__29037),
            .I(N__29033));
    InMux I__3019 (
            .O(N__29036),
            .I(N__29030));
    LocalMux I__3018 (
            .O(N__29033),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__3017 (
            .O(N__29030),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__3016 (
            .O(N__29025),
            .I(\c0.tx.n19728 ));
    InMux I__3015 (
            .O(N__29022),
            .I(N__29018));
    InMux I__3014 (
            .O(N__29021),
            .I(N__29015));
    LocalMux I__3013 (
            .O(N__29018),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__3012 (
            .O(N__29015),
            .I(\c0.tx.r_Clock_Count_7 ));
    InMux I__3011 (
            .O(N__29010),
            .I(\c0.tx.n19729 ));
    InMux I__3010 (
            .O(N__29007),
            .I(bfn_9_17_0_));
    CascadeMux I__3009 (
            .O(N__29004),
            .I(N__29000));
    InMux I__3008 (
            .O(N__29003),
            .I(N__28993));
    InMux I__3007 (
            .O(N__29000),
            .I(N__28993));
    InMux I__3006 (
            .O(N__28999),
            .I(N__28988));
    InMux I__3005 (
            .O(N__28998),
            .I(N__28988));
    LocalMux I__3004 (
            .O(N__28993),
            .I(N__28984));
    LocalMux I__3003 (
            .O(N__28988),
            .I(N__28981));
    InMux I__3002 (
            .O(N__28987),
            .I(N__28978));
    Span4Mux_v I__3001 (
            .O(N__28984),
            .I(N__28975));
    Span4Mux_h I__3000 (
            .O(N__28981),
            .I(N__28972));
    LocalMux I__2999 (
            .O(N__28978),
            .I(\c0.tx.r_Clock_Count_8 ));
    Odrv4 I__2998 (
            .O(N__28975),
            .I(\c0.tx.r_Clock_Count_8 ));
    Odrv4 I__2997 (
            .O(N__28972),
            .I(\c0.tx.r_Clock_Count_8 ));
    SRMux I__2996 (
            .O(N__28965),
            .I(N__28961));
    SRMux I__2995 (
            .O(N__28964),
            .I(N__28958));
    LocalMux I__2994 (
            .O(N__28961),
            .I(N__28955));
    LocalMux I__2993 (
            .O(N__28958),
            .I(N__28952));
    Span4Mux_h I__2992 (
            .O(N__28955),
            .I(N__28948));
    Span4Mux_h I__2991 (
            .O(N__28952),
            .I(N__28945));
    InMux I__2990 (
            .O(N__28951),
            .I(N__28942));
    Odrv4 I__2989 (
            .O(N__28948),
            .I(\c0.tx.n17199 ));
    Odrv4 I__2988 (
            .O(N__28945),
            .I(\c0.tx.n17199 ));
    LocalMux I__2987 (
            .O(N__28942),
            .I(\c0.tx.n17199 ));
    InMux I__2986 (
            .O(N__28935),
            .I(N__28932));
    LocalMux I__2985 (
            .O(N__28932),
            .I(N__28929));
    Span4Mux_v I__2984 (
            .O(N__28929),
            .I(N__28926));
    Odrv4 I__2983 (
            .O(N__28926),
            .I(\c0.tx.n4 ));
    CascadeMux I__2982 (
            .O(N__28923),
            .I(\c0.tx.n14290_cascade_ ));
    InMux I__2981 (
            .O(N__28920),
            .I(N__28917));
    LocalMux I__2980 (
            .O(N__28917),
            .I(N__28913));
    InMux I__2979 (
            .O(N__28916),
            .I(N__28910));
    Span4Mux_h I__2978 (
            .O(N__28913),
            .I(N__28907));
    LocalMux I__2977 (
            .O(N__28910),
            .I(data_out_frame_6_7));
    Odrv4 I__2976 (
            .O(N__28907),
            .I(data_out_frame_6_7));
    InMux I__2975 (
            .O(N__28902),
            .I(N__28899));
    LocalMux I__2974 (
            .O(N__28899),
            .I(\c0.n26_adj_4645 ));
    InMux I__2973 (
            .O(N__28896),
            .I(N__28893));
    LocalMux I__2972 (
            .O(N__28893),
            .I(n24808));
    InMux I__2971 (
            .O(N__28890),
            .I(N__28887));
    LocalMux I__2970 (
            .O(N__28887),
            .I(N__28884));
    Odrv4 I__2969 (
            .O(N__28884),
            .I(n10_adj_4779));
    CascadeMux I__2968 (
            .O(N__28881),
            .I(\c0.tx.n5_cascade_ ));
    InMux I__2967 (
            .O(N__28878),
            .I(N__28872));
    InMux I__2966 (
            .O(N__28877),
            .I(N__28865));
    InMux I__2965 (
            .O(N__28876),
            .I(N__28865));
    InMux I__2964 (
            .O(N__28875),
            .I(N__28865));
    LocalMux I__2963 (
            .O(N__28872),
            .I(N__28862));
    LocalMux I__2962 (
            .O(N__28865),
            .I(N__28859));
    Span4Mux_h I__2961 (
            .O(N__28862),
            .I(N__28856));
    Span4Mux_h I__2960 (
            .O(N__28859),
            .I(N__28853));
    Odrv4 I__2959 (
            .O(N__28856),
            .I(\c0.tx.n17904 ));
    Odrv4 I__2958 (
            .O(N__28853),
            .I(\c0.tx.n17904 ));
    InMux I__2957 (
            .O(N__28848),
            .I(N__28845));
    LocalMux I__2956 (
            .O(N__28845),
            .I(N__28842));
    Odrv12 I__2955 (
            .O(N__28842),
            .I(\c0.tx.n25051 ));
    InMux I__2954 (
            .O(N__28839),
            .I(bfn_9_16_0_));
    InMux I__2953 (
            .O(N__28836),
            .I(N__28832));
    InMux I__2952 (
            .O(N__28835),
            .I(N__28829));
    LocalMux I__2951 (
            .O(N__28832),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__2950 (
            .O(N__28829),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__2949 (
            .O(N__28824),
            .I(\c0.tx.n19723 ));
    InMux I__2948 (
            .O(N__28821),
            .I(N__28817));
    InMux I__2947 (
            .O(N__28820),
            .I(N__28814));
    LocalMux I__2946 (
            .O(N__28817),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__2945 (
            .O(N__28814),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__2944 (
            .O(N__28809),
            .I(\c0.tx.n19724 ));
    CascadeMux I__2943 (
            .O(N__28806),
            .I(n10_adj_4776_cascade_));
    InMux I__2942 (
            .O(N__28803),
            .I(N__28797));
    InMux I__2941 (
            .O(N__28802),
            .I(N__28797));
    LocalMux I__2940 (
            .O(N__28797),
            .I(r_Tx_Data_5));
    InMux I__2939 (
            .O(N__28794),
            .I(N__28791));
    LocalMux I__2938 (
            .O(N__28791),
            .I(\c0.tx.n25077 ));
    InMux I__2937 (
            .O(N__28788),
            .I(N__28782));
    InMux I__2936 (
            .O(N__28787),
            .I(N__28782));
    LocalMux I__2935 (
            .O(N__28782),
            .I(r_Tx_Data_7));
    CascadeMux I__2934 (
            .O(N__28779),
            .I(N__28775));
    InMux I__2933 (
            .O(N__28778),
            .I(N__28771));
    InMux I__2932 (
            .O(N__28775),
            .I(N__28768));
    InMux I__2931 (
            .O(N__28774),
            .I(N__28763));
    LocalMux I__2930 (
            .O(N__28771),
            .I(N__28758));
    LocalMux I__2929 (
            .O(N__28768),
            .I(N__28758));
    InMux I__2928 (
            .O(N__28767),
            .I(N__28752));
    InMux I__2927 (
            .O(N__28766),
            .I(N__28752));
    LocalMux I__2926 (
            .O(N__28763),
            .I(N__28749));
    Span4Mux_v I__2925 (
            .O(N__28758),
            .I(N__28746));
    InMux I__2924 (
            .O(N__28757),
            .I(N__28743));
    LocalMux I__2923 (
            .O(N__28752),
            .I(N__28740));
    Span4Mux_v I__2922 (
            .O(N__28749),
            .I(N__28735));
    Span4Mux_h I__2921 (
            .O(N__28746),
            .I(N__28735));
    LocalMux I__2920 (
            .O(N__28743),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv4 I__2919 (
            .O(N__28740),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv4 I__2918 (
            .O(N__28735),
            .I(\c0.tx.r_Bit_Index_0 ));
    CascadeMux I__2917 (
            .O(N__28728),
            .I(N__28723));
    InMux I__2916 (
            .O(N__28727),
            .I(N__28716));
    InMux I__2915 (
            .O(N__28726),
            .I(N__28713));
    InMux I__2914 (
            .O(N__28723),
            .I(N__28710));
    InMux I__2913 (
            .O(N__28722),
            .I(N__28701));
    InMux I__2912 (
            .O(N__28721),
            .I(N__28701));
    InMux I__2911 (
            .O(N__28720),
            .I(N__28701));
    InMux I__2910 (
            .O(N__28719),
            .I(N__28701));
    LocalMux I__2909 (
            .O(N__28716),
            .I(\c0.tx.r_Bit_Index_1 ));
    LocalMux I__2908 (
            .O(N__28713),
            .I(\c0.tx.r_Bit_Index_1 ));
    LocalMux I__2907 (
            .O(N__28710),
            .I(\c0.tx.r_Bit_Index_1 ));
    LocalMux I__2906 (
            .O(N__28701),
            .I(\c0.tx.r_Bit_Index_1 ));
    InMux I__2905 (
            .O(N__28692),
            .I(N__28689));
    LocalMux I__2904 (
            .O(N__28689),
            .I(\c0.tx.n25074 ));
    CascadeMux I__2903 (
            .O(N__28686),
            .I(N__28680));
    InMux I__2902 (
            .O(N__28685),
            .I(N__28676));
    InMux I__2901 (
            .O(N__28684),
            .I(N__28673));
    CascadeMux I__2900 (
            .O(N__28683),
            .I(N__28670));
    InMux I__2899 (
            .O(N__28680),
            .I(N__28663));
    InMux I__2898 (
            .O(N__28679),
            .I(N__28660));
    LocalMux I__2897 (
            .O(N__28676),
            .I(N__28655));
    LocalMux I__2896 (
            .O(N__28673),
            .I(N__28655));
    InMux I__2895 (
            .O(N__28670),
            .I(N__28652));
    InMux I__2894 (
            .O(N__28669),
            .I(N__28649));
    InMux I__2893 (
            .O(N__28668),
            .I(N__28644));
    InMux I__2892 (
            .O(N__28667),
            .I(N__28644));
    InMux I__2891 (
            .O(N__28666),
            .I(N__28641));
    LocalMux I__2890 (
            .O(N__28663),
            .I(N__28636));
    LocalMux I__2889 (
            .O(N__28660),
            .I(N__28636));
    Span4Mux_v I__2888 (
            .O(N__28655),
            .I(N__28633));
    LocalMux I__2887 (
            .O(N__28652),
            .I(N__28626));
    LocalMux I__2886 (
            .O(N__28649),
            .I(N__28626));
    LocalMux I__2885 (
            .O(N__28644),
            .I(N__28626));
    LocalMux I__2884 (
            .O(N__28641),
            .I(r_SM_Main_0));
    Odrv4 I__2883 (
            .O(N__28636),
            .I(r_SM_Main_0));
    Odrv4 I__2882 (
            .O(N__28633),
            .I(r_SM_Main_0));
    Odrv12 I__2881 (
            .O(N__28626),
            .I(r_SM_Main_0));
    CascadeMux I__2880 (
            .O(N__28617),
            .I(\c0.n24960_cascade_ ));
    CascadeMux I__2879 (
            .O(N__28614),
            .I(\c0.n24806_cascade_ ));
    InMux I__2878 (
            .O(N__28611),
            .I(N__28608));
    LocalMux I__2877 (
            .O(N__28608),
            .I(N__28605));
    Odrv4 I__2876 (
            .O(N__28605),
            .I(n24757));
    CascadeMux I__2875 (
            .O(N__28602),
            .I(n3_cascade_));
    IoInMux I__2874 (
            .O(N__28599),
            .I(N__28596));
    LocalMux I__2873 (
            .O(N__28596),
            .I(N__28593));
    IoSpan4Mux I__2872 (
            .O(N__28593),
            .I(N__28589));
    InMux I__2871 (
            .O(N__28592),
            .I(N__28586));
    Span4Mux_s0_h I__2870 (
            .O(N__28589),
            .I(N__28581));
    LocalMux I__2869 (
            .O(N__28586),
            .I(N__28581));
    Span4Mux_h I__2868 (
            .O(N__28581),
            .I(N__28578));
    Span4Mux_v I__2867 (
            .O(N__28578),
            .I(N__28575));
    Span4Mux_h I__2866 (
            .O(N__28575),
            .I(N__28571));
    InMux I__2865 (
            .O(N__28574),
            .I(N__28568));
    Odrv4 I__2864 (
            .O(N__28571),
            .I(tx_o));
    LocalMux I__2863 (
            .O(N__28568),
            .I(tx_o));
    InMux I__2862 (
            .O(N__28563),
            .I(N__28560));
    LocalMux I__2861 (
            .O(N__28560),
            .I(N__28556));
    InMux I__2860 (
            .O(N__28559),
            .I(N__28553));
    Span4Mux_h I__2859 (
            .O(N__28556),
            .I(N__28550));
    LocalMux I__2858 (
            .O(N__28553),
            .I(r_Tx_Data_3));
    Odrv4 I__2857 (
            .O(N__28550),
            .I(r_Tx_Data_3));
    InMux I__2856 (
            .O(N__28545),
            .I(N__28542));
    LocalMux I__2855 (
            .O(N__28542),
            .I(\c0.tx.n19492 ));
    InMux I__2854 (
            .O(N__28539),
            .I(N__28536));
    LocalMux I__2853 (
            .O(N__28536),
            .I(N__28533));
    Span4Mux_v I__2852 (
            .O(N__28533),
            .I(N__28527));
    InMux I__2851 (
            .O(N__28532),
            .I(N__28520));
    InMux I__2850 (
            .O(N__28531),
            .I(N__28520));
    InMux I__2849 (
            .O(N__28530),
            .I(N__28520));
    Odrv4 I__2848 (
            .O(N__28527),
            .I(\c0.tx.n22949 ));
    LocalMux I__2847 (
            .O(N__28520),
            .I(\c0.tx.n22949 ));
    CascadeMux I__2846 (
            .O(N__28515),
            .I(\c0.tx.n19492_cascade_ ));
    InMux I__2845 (
            .O(N__28512),
            .I(N__28509));
    LocalMux I__2844 (
            .O(N__28509),
            .I(N__28505));
    InMux I__2843 (
            .O(N__28508),
            .I(N__28502));
    Span4Mux_v I__2842 (
            .O(N__28505),
            .I(N__28499));
    LocalMux I__2841 (
            .O(N__28502),
            .I(r_Tx_Data_1));
    Odrv4 I__2840 (
            .O(N__28499),
            .I(r_Tx_Data_1));
    InMux I__2839 (
            .O(N__28494),
            .I(N__28491));
    LocalMux I__2838 (
            .O(N__28491),
            .I(\c0.tx.n25080 ));
    CascadeMux I__2837 (
            .O(N__28488),
            .I(\c0.tx.n25083_cascade_ ));
    InMux I__2836 (
            .O(N__28485),
            .I(N__28482));
    LocalMux I__2835 (
            .O(N__28482),
            .I(\c0.tx.o_Tx_Serial_N_3782 ));
    InMux I__2834 (
            .O(N__28479),
            .I(N__28476));
    LocalMux I__2833 (
            .O(N__28476),
            .I(N__28473));
    Span4Mux_h I__2832 (
            .O(N__28473),
            .I(N__28470));
    Odrv4 I__2831 (
            .O(N__28470),
            .I(n10));
    CascadeMux I__2830 (
            .O(N__28467),
            .I(N__28464));
    InMux I__2829 (
            .O(N__28464),
            .I(N__28459));
    InMux I__2828 (
            .O(N__28463),
            .I(N__28454));
    InMux I__2827 (
            .O(N__28462),
            .I(N__28454));
    LocalMux I__2826 (
            .O(N__28459),
            .I(\c0.tx.r_Bit_Index_2 ));
    LocalMux I__2825 (
            .O(N__28454),
            .I(\c0.tx.r_Bit_Index_2 ));
    CascadeMux I__2824 (
            .O(N__28449),
            .I(N__28446));
    InMux I__2823 (
            .O(N__28446),
            .I(N__28443));
    LocalMux I__2822 (
            .O(N__28443),
            .I(N__28440));
    Span4Mux_v I__2821 (
            .O(N__28440),
            .I(N__28436));
    InMux I__2820 (
            .O(N__28439),
            .I(N__28433));
    Odrv4 I__2819 (
            .O(N__28436),
            .I(\c0.tx.n17832 ));
    LocalMux I__2818 (
            .O(N__28433),
            .I(\c0.tx.n17832 ));
    InMux I__2817 (
            .O(N__28428),
            .I(\quad_counter1.n19714 ));
    InMux I__2816 (
            .O(N__28425),
            .I(\quad_counter1.n19715 ));
    CascadeMux I__2815 (
            .O(N__28422),
            .I(N__28419));
    InMux I__2814 (
            .O(N__28419),
            .I(N__28415));
    InMux I__2813 (
            .O(N__28418),
            .I(N__28411));
    LocalMux I__2812 (
            .O(N__28415),
            .I(N__28407));
    InMux I__2811 (
            .O(N__28414),
            .I(N__28402));
    LocalMux I__2810 (
            .O(N__28411),
            .I(N__28399));
    InMux I__2809 (
            .O(N__28410),
            .I(N__28396));
    Span4Mux_h I__2808 (
            .O(N__28407),
            .I(N__28393));
    InMux I__2807 (
            .O(N__28406),
            .I(N__28390));
    InMux I__2806 (
            .O(N__28405),
            .I(N__28387));
    LocalMux I__2805 (
            .O(N__28402),
            .I(\c0.tx.r_SM_Main_2 ));
    Odrv4 I__2804 (
            .O(N__28399),
            .I(\c0.tx.r_SM_Main_2 ));
    LocalMux I__2803 (
            .O(N__28396),
            .I(\c0.tx.r_SM_Main_2 ));
    Odrv4 I__2802 (
            .O(N__28393),
            .I(\c0.tx.r_SM_Main_2 ));
    LocalMux I__2801 (
            .O(N__28390),
            .I(\c0.tx.r_SM_Main_2 ));
    LocalMux I__2800 (
            .O(N__28387),
            .I(\c0.tx.r_SM_Main_2 ));
    InMux I__2799 (
            .O(N__28374),
            .I(N__28369));
    InMux I__2798 (
            .O(N__28373),
            .I(N__28366));
    InMux I__2797 (
            .O(N__28372),
            .I(N__28363));
    LocalMux I__2796 (
            .O(N__28369),
            .I(N__28358));
    LocalMux I__2795 (
            .O(N__28366),
            .I(N__28358));
    LocalMux I__2794 (
            .O(N__28363),
            .I(N__28352));
    Span4Mux_h I__2793 (
            .O(N__28358),
            .I(N__28352));
    InMux I__2792 (
            .O(N__28357),
            .I(N__28349));
    Span4Mux_v I__2791 (
            .O(N__28352),
            .I(N__28346));
    LocalMux I__2790 (
            .O(N__28349),
            .I(r_SM_Main_2_N_3751_1));
    Odrv4 I__2789 (
            .O(N__28346),
            .I(r_SM_Main_2_N_3751_1));
    InMux I__2788 (
            .O(N__28341),
            .I(N__28338));
    LocalMux I__2787 (
            .O(N__28338),
            .I(\c0.tx.n3843 ));
    InMux I__2786 (
            .O(N__28335),
            .I(\quad_counter1.n19705 ));
    InMux I__2785 (
            .O(N__28332),
            .I(\quad_counter1.n19706 ));
    InMux I__2784 (
            .O(N__28329),
            .I(\quad_counter1.n19707 ));
    InMux I__2783 (
            .O(N__28326),
            .I(bfn_9_8_0_));
    InMux I__2782 (
            .O(N__28323),
            .I(\quad_counter1.n19709 ));
    InMux I__2781 (
            .O(N__28320),
            .I(\quad_counter1.n19710 ));
    InMux I__2780 (
            .O(N__28317),
            .I(\quad_counter1.n19711 ));
    InMux I__2779 (
            .O(N__28314),
            .I(\quad_counter1.n19712 ));
    InMux I__2778 (
            .O(N__28311),
            .I(\quad_counter1.n19713 ));
    InMux I__2777 (
            .O(N__28308),
            .I(N__28304));
    InMux I__2776 (
            .O(N__28307),
            .I(N__28301));
    LocalMux I__2775 (
            .O(N__28304),
            .I(N__28298));
    LocalMux I__2774 (
            .O(N__28301),
            .I(data_out_frame_9_7));
    Odrv4 I__2773 (
            .O(N__28298),
            .I(data_out_frame_9_7));
    InMux I__2772 (
            .O(N__28293),
            .I(N__28290));
    LocalMux I__2771 (
            .O(N__28290),
            .I(N__28287));
    Odrv12 I__2770 (
            .O(N__28287),
            .I(\c0.rx.n24875 ));
    InMux I__2769 (
            .O(N__28284),
            .I(N__28281));
    LocalMux I__2768 (
            .O(N__28281),
            .I(\c0.rx.n25068 ));
    InMux I__2767 (
            .O(N__28278),
            .I(bfn_9_7_0_));
    InMux I__2766 (
            .O(N__28275),
            .I(\quad_counter1.n19701 ));
    InMux I__2765 (
            .O(N__28272),
            .I(\quad_counter1.n19702 ));
    InMux I__2764 (
            .O(N__28269),
            .I(\quad_counter1.n19703 ));
    InMux I__2763 (
            .O(N__28266),
            .I(\quad_counter1.n19704 ));
    CascadeMux I__2762 (
            .O(N__28263),
            .I(\c0.n25104_cascade_ ));
    InMux I__2761 (
            .O(N__28260),
            .I(N__28257));
    LocalMux I__2760 (
            .O(N__28257),
            .I(N__28254));
    Odrv12 I__2759 (
            .O(N__28254),
            .I(\c0.n25107 ));
    InMux I__2758 (
            .O(N__28251),
            .I(N__28247));
    InMux I__2757 (
            .O(N__28250),
            .I(N__28244));
    LocalMux I__2756 (
            .O(N__28247),
            .I(N__28241));
    LocalMux I__2755 (
            .O(N__28244),
            .I(data_out_frame_5_7));
    Odrv4 I__2754 (
            .O(N__28241),
            .I(data_out_frame_5_7));
    InMux I__2753 (
            .O(N__28236),
            .I(N__28233));
    LocalMux I__2752 (
            .O(N__28233),
            .I(n25071));
    CascadeMux I__2751 (
            .O(N__28230),
            .I(n3821_cascade_));
    CascadeMux I__2750 (
            .O(N__28227),
            .I(\c0.tx.n6_cascade_ ));
    InMux I__2749 (
            .O(N__28224),
            .I(N__28221));
    LocalMux I__2748 (
            .O(N__28221),
            .I(N__28218));
    Odrv4 I__2747 (
            .O(N__28218),
            .I(\c0.n25089 ));
    InMux I__2746 (
            .O(N__28215),
            .I(N__28212));
    LocalMux I__2745 (
            .O(N__28212),
            .I(N__28209));
    Odrv4 I__2744 (
            .O(N__28209),
            .I(n25018));
    InMux I__2743 (
            .O(N__28206),
            .I(N__28203));
    LocalMux I__2742 (
            .O(N__28203),
            .I(\c0.tx.n23980 ));
    CascadeMux I__2741 (
            .O(N__28200),
            .I(\c0.n5_adj_4712_cascade_ ));
    InMux I__2740 (
            .O(N__28197),
            .I(N__28194));
    LocalMux I__2739 (
            .O(N__28194),
            .I(N__28191));
    Odrv4 I__2738 (
            .O(N__28191),
            .I(\c0.n24800 ));
    InMux I__2737 (
            .O(N__28188),
            .I(N__28185));
    LocalMux I__2736 (
            .O(N__28185),
            .I(N__28182));
    Odrv4 I__2735 (
            .O(N__28182),
            .I(\c0.tx.n5_adj_4207 ));
    InMux I__2734 (
            .O(N__28179),
            .I(N__28176));
    LocalMux I__2733 (
            .O(N__28176),
            .I(\c0.n24949 ));
    InMux I__2732 (
            .O(N__28173),
            .I(N__28170));
    LocalMux I__2731 (
            .O(N__28170),
            .I(N__28167));
    Odrv4 I__2730 (
            .O(N__28167),
            .I(n10_adj_4777));
    CascadeMux I__2729 (
            .O(N__28164),
            .I(\c0.n25086_cascade_ ));
    InMux I__2728 (
            .O(N__28161),
            .I(N__28157));
    InMux I__2727 (
            .O(N__28160),
            .I(N__28154));
    LocalMux I__2726 (
            .O(N__28157),
            .I(data_out_frame_9_3));
    LocalMux I__2725 (
            .O(N__28154),
            .I(data_out_frame_9_3));
    CascadeMux I__2724 (
            .O(N__28149),
            .I(n24802_cascade_));
    CascadeMux I__2723 (
            .O(N__28146),
            .I(\c0.n11_adj_4715_cascade_ ));
    InMux I__2722 (
            .O(N__28143),
            .I(N__28140));
    LocalMux I__2721 (
            .O(N__28140),
            .I(n25010));
    InMux I__2720 (
            .O(N__28137),
            .I(N__28130));
    InMux I__2719 (
            .O(N__28136),
            .I(N__28125));
    InMux I__2718 (
            .O(N__28135),
            .I(N__28125));
    InMux I__2717 (
            .O(N__28134),
            .I(N__28122));
    InMux I__2716 (
            .O(N__28133),
            .I(N__28119));
    LocalMux I__2715 (
            .O(N__28130),
            .I(N__28114));
    LocalMux I__2714 (
            .O(N__28125),
            .I(N__28114));
    LocalMux I__2713 (
            .O(N__28122),
            .I(N__28111));
    LocalMux I__2712 (
            .O(N__28119),
            .I(N__28106));
    Span4Mux_h I__2711 (
            .O(N__28114),
            .I(N__28106));
    Odrv4 I__2710 (
            .O(N__28111),
            .I(A_filtered));
    Odrv4 I__2709 (
            .O(N__28106),
            .I(A_filtered));
    InMux I__2708 (
            .O(N__28101),
            .I(N__28098));
    LocalMux I__2707 (
            .O(N__28098),
            .I(n8628));
    CascadeMux I__2706 (
            .O(N__28095),
            .I(n9603_cascade_));
    CascadeMux I__2705 (
            .O(N__28092),
            .I(N__28087));
    InMux I__2704 (
            .O(N__28091),
            .I(N__28084));
    CascadeMux I__2703 (
            .O(N__28090),
            .I(N__28081));
    InMux I__2702 (
            .O(N__28087),
            .I(N__28078));
    LocalMux I__2701 (
            .O(N__28084),
            .I(N__28075));
    InMux I__2700 (
            .O(N__28081),
            .I(N__28072));
    LocalMux I__2699 (
            .O(N__28078),
            .I(B_filtered));
    Odrv4 I__2698 (
            .O(N__28075),
            .I(B_filtered));
    LocalMux I__2697 (
            .O(N__28072),
            .I(B_filtered));
    CascadeMux I__2696 (
            .O(N__28065),
            .I(N__28061));
    InMux I__2695 (
            .O(N__28064),
            .I(N__28057));
    InMux I__2694 (
            .O(N__28061),
            .I(N__28052));
    InMux I__2693 (
            .O(N__28060),
            .I(N__28052));
    LocalMux I__2692 (
            .O(N__28057),
            .I(N__28047));
    LocalMux I__2691 (
            .O(N__28052),
            .I(N__28047));
    Odrv4 I__2690 (
            .O(N__28047),
            .I(\quad_counter0.B_delayed ));
    InMux I__2689 (
            .O(N__28044),
            .I(\quad_counter0.n19685 ));
    InMux I__2688 (
            .O(N__28041),
            .I(N__28037));
    InMux I__2687 (
            .O(N__28040),
            .I(N__28034));
    LocalMux I__2686 (
            .O(N__28037),
            .I(\quad_counter0.a_delay_counter_15 ));
    LocalMux I__2685 (
            .O(N__28034),
            .I(\quad_counter0.a_delay_counter_15 ));
    CascadeMux I__2684 (
            .O(N__28029),
            .I(N__28026));
    InMux I__2683 (
            .O(N__28026),
            .I(N__28021));
    CEMux I__2682 (
            .O(N__28025),
            .I(N__28018));
    CEMux I__2681 (
            .O(N__28024),
            .I(N__28015));
    LocalMux I__2680 (
            .O(N__28021),
            .I(n14469));
    LocalMux I__2679 (
            .O(N__28018),
            .I(n14469));
    LocalMux I__2678 (
            .O(N__28015),
            .I(n14469));
    SRMux I__2677 (
            .O(N__28008),
            .I(N__28004));
    InMux I__2676 (
            .O(N__28007),
            .I(N__28000));
    LocalMux I__2675 (
            .O(N__28004),
            .I(N__27997));
    SRMux I__2674 (
            .O(N__28003),
            .I(N__27994));
    LocalMux I__2673 (
            .O(N__28000),
            .I(N__27991));
    Odrv12 I__2672 (
            .O(N__27997),
            .I(a_delay_counter_15__N_4123));
    LocalMux I__2671 (
            .O(N__27994),
            .I(a_delay_counter_15__N_4123));
    Odrv4 I__2670 (
            .O(N__27991),
            .I(a_delay_counter_15__N_4123));
    InMux I__2669 (
            .O(N__27984),
            .I(N__27980));
    InMux I__2668 (
            .O(N__27983),
            .I(N__27977));
    LocalMux I__2667 (
            .O(N__27980),
            .I(N__27974));
    LocalMux I__2666 (
            .O(N__27977),
            .I(\quad_counter1.b_delay_counter_13 ));
    Odrv4 I__2665 (
            .O(N__27974),
            .I(\quad_counter1.b_delay_counter_13 ));
    InMux I__2664 (
            .O(N__27969),
            .I(N__27965));
    InMux I__2663 (
            .O(N__27968),
            .I(N__27962));
    LocalMux I__2662 (
            .O(N__27965),
            .I(\quad_counter1.b_delay_counter_1 ));
    LocalMux I__2661 (
            .O(N__27962),
            .I(\quad_counter1.b_delay_counter_1 ));
    CascadeMux I__2660 (
            .O(N__27957),
            .I(N__27953));
    InMux I__2659 (
            .O(N__27956),
            .I(N__27950));
    InMux I__2658 (
            .O(N__27953),
            .I(N__27947));
    LocalMux I__2657 (
            .O(N__27950),
            .I(\quad_counter1.b_delay_counter_2 ));
    LocalMux I__2656 (
            .O(N__27947),
            .I(\quad_counter1.b_delay_counter_2 ));
    InMux I__2655 (
            .O(N__27942),
            .I(N__27938));
    InMux I__2654 (
            .O(N__27941),
            .I(N__27935));
    LocalMux I__2653 (
            .O(N__27938),
            .I(\quad_counter1.b_delay_counter_5 ));
    LocalMux I__2652 (
            .O(N__27935),
            .I(\quad_counter1.b_delay_counter_5 ));
    InMux I__2651 (
            .O(N__27930),
            .I(N__27927));
    LocalMux I__2650 (
            .O(N__27927),
            .I(N__27924));
    Odrv4 I__2649 (
            .O(N__27924),
            .I(\quad_counter1.n28_adj_4199 ));
    InMux I__2648 (
            .O(N__27921),
            .I(N__27916));
    InMux I__2647 (
            .O(N__27920),
            .I(N__27913));
    InMux I__2646 (
            .O(N__27919),
            .I(N__27910));
    LocalMux I__2645 (
            .O(N__27916),
            .I(N__27904));
    LocalMux I__2644 (
            .O(N__27913),
            .I(N__27904));
    LocalMux I__2643 (
            .O(N__27910),
            .I(N__27901));
    InMux I__2642 (
            .O(N__27909),
            .I(N__27898));
    Span4Mux_v I__2641 (
            .O(N__27904),
            .I(N__27891));
    Span4Mux_h I__2640 (
            .O(N__27901),
            .I(N__27891));
    LocalMux I__2639 (
            .O(N__27898),
            .I(N__27891));
    Span4Mux_h I__2638 (
            .O(N__27891),
            .I(N__27888));
    Span4Mux_v I__2637 (
            .O(N__27888),
            .I(N__27885));
    Odrv4 I__2636 (
            .O(N__27885),
            .I(PIN_7_c));
    InMux I__2635 (
            .O(N__27882),
            .I(N__27878));
    CascadeMux I__2634 (
            .O(N__27881),
            .I(N__27875));
    LocalMux I__2633 (
            .O(N__27878),
            .I(N__27872));
    InMux I__2632 (
            .O(N__27875),
            .I(N__27868));
    Span4Mux_h I__2631 (
            .O(N__27872),
            .I(N__27865));
    InMux I__2630 (
            .O(N__27871),
            .I(N__27862));
    LocalMux I__2629 (
            .O(N__27868),
            .I(quadA_delayed));
    Odrv4 I__2628 (
            .O(N__27865),
            .I(quadA_delayed));
    LocalMux I__2627 (
            .O(N__27862),
            .I(quadA_delayed));
    InMux I__2626 (
            .O(N__27855),
            .I(N__27851));
    InMux I__2625 (
            .O(N__27854),
            .I(N__27848));
    LocalMux I__2624 (
            .O(N__27851),
            .I(\quad_counter1.b_delay_counter_14 ));
    LocalMux I__2623 (
            .O(N__27848),
            .I(\quad_counter1.b_delay_counter_14 ));
    InMux I__2622 (
            .O(N__27843),
            .I(N__27839));
    InMux I__2621 (
            .O(N__27842),
            .I(N__27836));
    LocalMux I__2620 (
            .O(N__27839),
            .I(\quad_counter1.b_delay_counter_7 ));
    LocalMux I__2619 (
            .O(N__27836),
            .I(\quad_counter1.b_delay_counter_7 ));
    CascadeMux I__2618 (
            .O(N__27831),
            .I(N__27827));
    InMux I__2617 (
            .O(N__27830),
            .I(N__27824));
    InMux I__2616 (
            .O(N__27827),
            .I(N__27821));
    LocalMux I__2615 (
            .O(N__27824),
            .I(\quad_counter1.b_delay_counter_12 ));
    LocalMux I__2614 (
            .O(N__27821),
            .I(\quad_counter1.b_delay_counter_12 ));
    InMux I__2613 (
            .O(N__27816),
            .I(N__27812));
    InMux I__2612 (
            .O(N__27815),
            .I(N__27809));
    LocalMux I__2611 (
            .O(N__27812),
            .I(\quad_counter1.b_delay_counter_15 ));
    LocalMux I__2610 (
            .O(N__27809),
            .I(\quad_counter1.b_delay_counter_15 ));
    InMux I__2609 (
            .O(N__27804),
            .I(N__27801));
    LocalMux I__2608 (
            .O(N__27801),
            .I(\quad_counter1.n27_adj_4201 ));
    InMux I__2607 (
            .O(N__27798),
            .I(N__27794));
    InMux I__2606 (
            .O(N__27797),
            .I(N__27791));
    LocalMux I__2605 (
            .O(N__27794),
            .I(\quad_counter0.a_delay_counter_7 ));
    LocalMux I__2604 (
            .O(N__27791),
            .I(\quad_counter0.a_delay_counter_7 ));
    InMux I__2603 (
            .O(N__27786),
            .I(\quad_counter0.n19677 ));
    InMux I__2602 (
            .O(N__27783),
            .I(N__27779));
    InMux I__2601 (
            .O(N__27782),
            .I(N__27776));
    LocalMux I__2600 (
            .O(N__27779),
            .I(\quad_counter0.a_delay_counter_8 ));
    LocalMux I__2599 (
            .O(N__27776),
            .I(\quad_counter0.a_delay_counter_8 ));
    InMux I__2598 (
            .O(N__27771),
            .I(bfn_6_14_0_));
    InMux I__2597 (
            .O(N__27768),
            .I(N__27764));
    InMux I__2596 (
            .O(N__27767),
            .I(N__27761));
    LocalMux I__2595 (
            .O(N__27764),
            .I(\quad_counter0.a_delay_counter_9 ));
    LocalMux I__2594 (
            .O(N__27761),
            .I(\quad_counter0.a_delay_counter_9 ));
    InMux I__2593 (
            .O(N__27756),
            .I(\quad_counter0.n19679 ));
    CascadeMux I__2592 (
            .O(N__27753),
            .I(N__27749));
    InMux I__2591 (
            .O(N__27752),
            .I(N__27746));
    InMux I__2590 (
            .O(N__27749),
            .I(N__27743));
    LocalMux I__2589 (
            .O(N__27746),
            .I(\quad_counter0.a_delay_counter_10 ));
    LocalMux I__2588 (
            .O(N__27743),
            .I(\quad_counter0.a_delay_counter_10 ));
    InMux I__2587 (
            .O(N__27738),
            .I(\quad_counter0.n19680 ));
    InMux I__2586 (
            .O(N__27735),
            .I(N__27731));
    InMux I__2585 (
            .O(N__27734),
            .I(N__27728));
    LocalMux I__2584 (
            .O(N__27731),
            .I(\quad_counter0.a_delay_counter_11 ));
    LocalMux I__2583 (
            .O(N__27728),
            .I(\quad_counter0.a_delay_counter_11 ));
    InMux I__2582 (
            .O(N__27723),
            .I(\quad_counter0.n19681 ));
    InMux I__2581 (
            .O(N__27720),
            .I(N__27716));
    InMux I__2580 (
            .O(N__27719),
            .I(N__27713));
    LocalMux I__2579 (
            .O(N__27716),
            .I(\quad_counter0.a_delay_counter_12 ));
    LocalMux I__2578 (
            .O(N__27713),
            .I(\quad_counter0.a_delay_counter_12 ));
    InMux I__2577 (
            .O(N__27708),
            .I(\quad_counter0.n19682 ));
    InMux I__2576 (
            .O(N__27705),
            .I(N__27701));
    InMux I__2575 (
            .O(N__27704),
            .I(N__27698));
    LocalMux I__2574 (
            .O(N__27701),
            .I(\quad_counter0.a_delay_counter_13 ));
    LocalMux I__2573 (
            .O(N__27698),
            .I(\quad_counter0.a_delay_counter_13 ));
    InMux I__2572 (
            .O(N__27693),
            .I(\quad_counter0.n19683 ));
    InMux I__2571 (
            .O(N__27690),
            .I(N__27686));
    InMux I__2570 (
            .O(N__27689),
            .I(N__27683));
    LocalMux I__2569 (
            .O(N__27686),
            .I(\quad_counter0.a_delay_counter_14 ));
    LocalMux I__2568 (
            .O(N__27683),
            .I(\quad_counter0.a_delay_counter_14 ));
    InMux I__2567 (
            .O(N__27678),
            .I(\quad_counter0.n19684 ));
    InMux I__2566 (
            .O(N__27675),
            .I(N__27671));
    InMux I__2565 (
            .O(N__27674),
            .I(N__27668));
    LocalMux I__2564 (
            .O(N__27671),
            .I(\quad_counter0.b_delay_counter_10 ));
    LocalMux I__2563 (
            .O(N__27668),
            .I(\quad_counter0.b_delay_counter_10 ));
    InMux I__2562 (
            .O(N__27663),
            .I(N__27659));
    InMux I__2561 (
            .O(N__27662),
            .I(N__27656));
    LocalMux I__2560 (
            .O(N__27659),
            .I(\quad_counter0.b_delay_counter_11 ));
    LocalMux I__2559 (
            .O(N__27656),
            .I(\quad_counter0.b_delay_counter_11 ));
    CascadeMux I__2558 (
            .O(N__27651),
            .I(\quad_counter0.n24_adj_4758_cascade_ ));
    InMux I__2557 (
            .O(N__27648),
            .I(N__27645));
    LocalMux I__2556 (
            .O(N__27645),
            .I(\quad_counter0.n18 ));
    InMux I__2555 (
            .O(N__27642),
            .I(N__27639));
    LocalMux I__2554 (
            .O(N__27639),
            .I(\quad_counter0.n26_adj_4759 ));
    InMux I__2553 (
            .O(N__27636),
            .I(N__27631));
    InMux I__2552 (
            .O(N__27635),
            .I(N__27626));
    InMux I__2551 (
            .O(N__27634),
            .I(N__27626));
    LocalMux I__2550 (
            .O(N__27631),
            .I(a_delay_counter_0));
    LocalMux I__2549 (
            .O(N__27626),
            .I(a_delay_counter_0));
    InMux I__2548 (
            .O(N__27621),
            .I(N__27618));
    LocalMux I__2547 (
            .O(N__27618),
            .I(N__27615));
    Odrv4 I__2546 (
            .O(N__27615),
            .I(n39));
    InMux I__2545 (
            .O(N__27612),
            .I(bfn_6_13_0_));
    InMux I__2544 (
            .O(N__27609),
            .I(N__27605));
    InMux I__2543 (
            .O(N__27608),
            .I(N__27602));
    LocalMux I__2542 (
            .O(N__27605),
            .I(\quad_counter0.a_delay_counter_1 ));
    LocalMux I__2541 (
            .O(N__27602),
            .I(\quad_counter0.a_delay_counter_1 ));
    InMux I__2540 (
            .O(N__27597),
            .I(\quad_counter0.n19671 ));
    CascadeMux I__2539 (
            .O(N__27594),
            .I(N__27590));
    InMux I__2538 (
            .O(N__27593),
            .I(N__27587));
    InMux I__2537 (
            .O(N__27590),
            .I(N__27584));
    LocalMux I__2536 (
            .O(N__27587),
            .I(\quad_counter0.a_delay_counter_2 ));
    LocalMux I__2535 (
            .O(N__27584),
            .I(\quad_counter0.a_delay_counter_2 ));
    InMux I__2534 (
            .O(N__27579),
            .I(\quad_counter0.n19672 ));
    InMux I__2533 (
            .O(N__27576),
            .I(N__27572));
    InMux I__2532 (
            .O(N__27575),
            .I(N__27569));
    LocalMux I__2531 (
            .O(N__27572),
            .I(\quad_counter0.a_delay_counter_3 ));
    LocalMux I__2530 (
            .O(N__27569),
            .I(\quad_counter0.a_delay_counter_3 ));
    InMux I__2529 (
            .O(N__27564),
            .I(\quad_counter0.n19673 ));
    CascadeMux I__2528 (
            .O(N__27561),
            .I(N__27557));
    InMux I__2527 (
            .O(N__27560),
            .I(N__27554));
    InMux I__2526 (
            .O(N__27557),
            .I(N__27551));
    LocalMux I__2525 (
            .O(N__27554),
            .I(\quad_counter0.a_delay_counter_4 ));
    LocalMux I__2524 (
            .O(N__27551),
            .I(\quad_counter0.a_delay_counter_4 ));
    InMux I__2523 (
            .O(N__27546),
            .I(\quad_counter0.n19674 ));
    InMux I__2522 (
            .O(N__27543),
            .I(N__27539));
    InMux I__2521 (
            .O(N__27542),
            .I(N__27536));
    LocalMux I__2520 (
            .O(N__27539),
            .I(\quad_counter0.a_delay_counter_5 ));
    LocalMux I__2519 (
            .O(N__27536),
            .I(\quad_counter0.a_delay_counter_5 ));
    InMux I__2518 (
            .O(N__27531),
            .I(\quad_counter0.n19675 ));
    CascadeMux I__2517 (
            .O(N__27528),
            .I(N__27524));
    InMux I__2516 (
            .O(N__27527),
            .I(N__27521));
    InMux I__2515 (
            .O(N__27524),
            .I(N__27518));
    LocalMux I__2514 (
            .O(N__27521),
            .I(\quad_counter0.a_delay_counter_6 ));
    LocalMux I__2513 (
            .O(N__27518),
            .I(\quad_counter0.a_delay_counter_6 ));
    InMux I__2512 (
            .O(N__27513),
            .I(\quad_counter0.n19676 ));
    InMux I__2511 (
            .O(N__27510),
            .I(\quad_counter0.n19666 ));
    InMux I__2510 (
            .O(N__27507),
            .I(\quad_counter0.n19667 ));
    InMux I__2509 (
            .O(N__27504),
            .I(N__27500));
    InMux I__2508 (
            .O(N__27503),
            .I(N__27497));
    LocalMux I__2507 (
            .O(N__27500),
            .I(\quad_counter0.b_delay_counter_13 ));
    LocalMux I__2506 (
            .O(N__27497),
            .I(\quad_counter0.b_delay_counter_13 ));
    InMux I__2505 (
            .O(N__27492),
            .I(\quad_counter0.n19668 ));
    InMux I__2504 (
            .O(N__27489),
            .I(\quad_counter0.n19669 ));
    InMux I__2503 (
            .O(N__27486),
            .I(\quad_counter0.n19670 ));
    CEMux I__2502 (
            .O(N__27483),
            .I(N__27479));
    CEMux I__2501 (
            .O(N__27482),
            .I(N__27476));
    LocalMux I__2500 (
            .O(N__27479),
            .I(N__27473));
    LocalMux I__2499 (
            .O(N__27476),
            .I(N__27470));
    Span4Mux_v I__2498 (
            .O(N__27473),
            .I(N__27466));
    Span4Mux_v I__2497 (
            .O(N__27470),
            .I(N__27463));
    InMux I__2496 (
            .O(N__27469),
            .I(N__27460));
    Odrv4 I__2495 (
            .O(N__27466),
            .I(n14315));
    Odrv4 I__2494 (
            .O(N__27463),
            .I(n14315));
    LocalMux I__2493 (
            .O(N__27460),
            .I(n14315));
    SRMux I__2492 (
            .O(N__27453),
            .I(N__27449));
    SRMux I__2491 (
            .O(N__27452),
            .I(N__27445));
    LocalMux I__2490 (
            .O(N__27449),
            .I(N__27442));
    InMux I__2489 (
            .O(N__27448),
            .I(N__27439));
    LocalMux I__2488 (
            .O(N__27445),
            .I(N__27435));
    Span4Mux_h I__2487 (
            .O(N__27442),
            .I(N__27432));
    LocalMux I__2486 (
            .O(N__27439),
            .I(N__27429));
    InMux I__2485 (
            .O(N__27438),
            .I(N__27426));
    Odrv4 I__2484 (
            .O(N__27435),
            .I(b_delay_counter_15__N_4140));
    Odrv4 I__2483 (
            .O(N__27432),
            .I(b_delay_counter_15__N_4140));
    Odrv4 I__2482 (
            .O(N__27429),
            .I(b_delay_counter_15__N_4140));
    LocalMux I__2481 (
            .O(N__27426),
            .I(b_delay_counter_15__N_4140));
    InMux I__2480 (
            .O(N__27417),
            .I(N__27413));
    InMux I__2479 (
            .O(N__27416),
            .I(N__27408));
    LocalMux I__2478 (
            .O(N__27413),
            .I(N__27405));
    InMux I__2477 (
            .O(N__27412),
            .I(N__27402));
    InMux I__2476 (
            .O(N__27411),
            .I(N__27399));
    LocalMux I__2475 (
            .O(N__27408),
            .I(N__27392));
    Span4Mux_h I__2474 (
            .O(N__27405),
            .I(N__27392));
    LocalMux I__2473 (
            .O(N__27402),
            .I(N__27392));
    LocalMux I__2472 (
            .O(N__27399),
            .I(N__27389));
    Sp12to4 I__2471 (
            .O(N__27392),
            .I(N__27386));
    Span4Mux_h I__2470 (
            .O(N__27389),
            .I(N__27383));
    Span12Mux_v I__2469 (
            .O(N__27386),
            .I(N__27380));
    Span4Mux_v I__2468 (
            .O(N__27383),
            .I(N__27377));
    Odrv12 I__2467 (
            .O(N__27380),
            .I(PIN_8_c));
    Odrv4 I__2466 (
            .O(N__27377),
            .I(PIN_8_c));
    InMux I__2465 (
            .O(N__27372),
            .I(N__27369));
    LocalMux I__2464 (
            .O(N__27369),
            .I(N__27365));
    InMux I__2463 (
            .O(N__27368),
            .I(N__27362));
    Span4Mux_v I__2462 (
            .O(N__27365),
            .I(N__27358));
    LocalMux I__2461 (
            .O(N__27362),
            .I(N__27355));
    InMux I__2460 (
            .O(N__27361),
            .I(N__27352));
    Odrv4 I__2459 (
            .O(N__27358),
            .I(quadB_delayed));
    Odrv4 I__2458 (
            .O(N__27355),
            .I(quadB_delayed));
    LocalMux I__2457 (
            .O(N__27352),
            .I(quadB_delayed));
    InMux I__2456 (
            .O(N__27345),
            .I(N__27342));
    LocalMux I__2455 (
            .O(N__27342),
            .I(n12942));
    InMux I__2454 (
            .O(N__27339),
            .I(N__27335));
    InMux I__2453 (
            .O(N__27338),
            .I(N__27332));
    LocalMux I__2452 (
            .O(N__27335),
            .I(\quad_counter0.b_delay_counter_15 ));
    LocalMux I__2451 (
            .O(N__27332),
            .I(\quad_counter0.b_delay_counter_15 ));
    InMux I__2450 (
            .O(N__27327),
            .I(N__27323));
    InMux I__2449 (
            .O(N__27326),
            .I(N__27320));
    LocalMux I__2448 (
            .O(N__27323),
            .I(\quad_counter0.b_delay_counter_8 ));
    LocalMux I__2447 (
            .O(N__27320),
            .I(\quad_counter0.b_delay_counter_8 ));
    InMux I__2446 (
            .O(N__27315),
            .I(N__27312));
    LocalMux I__2445 (
            .O(N__27312),
            .I(\quad_counter0.A_delayed ));
    InMux I__2444 (
            .O(N__27309),
            .I(N__27305));
    InMux I__2443 (
            .O(N__27308),
            .I(N__27302));
    LocalMux I__2442 (
            .O(N__27305),
            .I(N__27299));
    LocalMux I__2441 (
            .O(N__27302),
            .I(\quad_counter0.b_delay_counter_7 ));
    Odrv4 I__2440 (
            .O(N__27299),
            .I(\quad_counter0.b_delay_counter_7 ));
    InMux I__2439 (
            .O(N__27294),
            .I(N__27290));
    InMux I__2438 (
            .O(N__27293),
            .I(N__27287));
    LocalMux I__2437 (
            .O(N__27290),
            .I(\quad_counter0.b_delay_counter_12 ));
    LocalMux I__2436 (
            .O(N__27287),
            .I(\quad_counter0.b_delay_counter_12 ));
    CascadeMux I__2435 (
            .O(N__27282),
            .I(N__27279));
    InMux I__2434 (
            .O(N__27279),
            .I(N__27275));
    InMux I__2433 (
            .O(N__27278),
            .I(N__27272));
    LocalMux I__2432 (
            .O(N__27275),
            .I(N__27269));
    LocalMux I__2431 (
            .O(N__27272),
            .I(\quad_counter0.b_delay_counter_5 ));
    Odrv4 I__2430 (
            .O(N__27269),
            .I(\quad_counter0.b_delay_counter_5 ));
    InMux I__2429 (
            .O(N__27264),
            .I(N__27260));
    InMux I__2428 (
            .O(N__27263),
            .I(N__27257));
    LocalMux I__2427 (
            .O(N__27260),
            .I(\quad_counter0.b_delay_counter_14 ));
    LocalMux I__2426 (
            .O(N__27257),
            .I(\quad_counter0.b_delay_counter_14 ));
    InMux I__2425 (
            .O(N__27252),
            .I(N__27248));
    InMux I__2424 (
            .O(N__27251),
            .I(N__27245));
    LocalMux I__2423 (
            .O(N__27248),
            .I(\quad_counter0.b_delay_counter_2 ));
    LocalMux I__2422 (
            .O(N__27245),
            .I(\quad_counter0.b_delay_counter_2 ));
    InMux I__2421 (
            .O(N__27240),
            .I(\quad_counter0.n19657 ));
    InMux I__2420 (
            .O(N__27237),
            .I(N__27233));
    InMux I__2419 (
            .O(N__27236),
            .I(N__27230));
    LocalMux I__2418 (
            .O(N__27233),
            .I(\quad_counter0.b_delay_counter_3 ));
    LocalMux I__2417 (
            .O(N__27230),
            .I(\quad_counter0.b_delay_counter_3 ));
    InMux I__2416 (
            .O(N__27225),
            .I(\quad_counter0.n19658 ));
    InMux I__2415 (
            .O(N__27222),
            .I(N__27218));
    InMux I__2414 (
            .O(N__27221),
            .I(N__27215));
    LocalMux I__2413 (
            .O(N__27218),
            .I(\quad_counter0.b_delay_counter_4 ));
    LocalMux I__2412 (
            .O(N__27215),
            .I(\quad_counter0.b_delay_counter_4 ));
    InMux I__2411 (
            .O(N__27210),
            .I(\quad_counter0.n19659 ));
    InMux I__2410 (
            .O(N__27207),
            .I(\quad_counter0.n19660 ));
    CascadeMux I__2409 (
            .O(N__27204),
            .I(N__27200));
    InMux I__2408 (
            .O(N__27203),
            .I(N__27197));
    InMux I__2407 (
            .O(N__27200),
            .I(N__27194));
    LocalMux I__2406 (
            .O(N__27197),
            .I(\quad_counter0.b_delay_counter_6 ));
    LocalMux I__2405 (
            .O(N__27194),
            .I(\quad_counter0.b_delay_counter_6 ));
    InMux I__2404 (
            .O(N__27189),
            .I(\quad_counter0.n19661 ));
    InMux I__2403 (
            .O(N__27186),
            .I(\quad_counter0.n19662 ));
    InMux I__2402 (
            .O(N__27183),
            .I(bfn_6_11_0_));
    InMux I__2401 (
            .O(N__27180),
            .I(N__27176));
    InMux I__2400 (
            .O(N__27179),
            .I(N__27173));
    LocalMux I__2399 (
            .O(N__27176),
            .I(\quad_counter0.b_delay_counter_9 ));
    LocalMux I__2398 (
            .O(N__27173),
            .I(\quad_counter0.b_delay_counter_9 ));
    InMux I__2397 (
            .O(N__27168),
            .I(\quad_counter0.n19664 ));
    InMux I__2396 (
            .O(N__27165),
            .I(\quad_counter0.n19665 ));
    InMux I__2395 (
            .O(N__27162),
            .I(N__27158));
    InMux I__2394 (
            .O(N__27161),
            .I(N__27155));
    LocalMux I__2393 (
            .O(N__27158),
            .I(N__27152));
    LocalMux I__2392 (
            .O(N__27155),
            .I(\quad_counter1.b_delay_counter_10 ));
    Odrv4 I__2391 (
            .O(N__27152),
            .I(\quad_counter1.b_delay_counter_10 ));
    InMux I__2390 (
            .O(N__27147),
            .I(\quad_counter1.n19695 ));
    InMux I__2389 (
            .O(N__27144),
            .I(N__27140));
    InMux I__2388 (
            .O(N__27143),
            .I(N__27137));
    LocalMux I__2387 (
            .O(N__27140),
            .I(N__27134));
    LocalMux I__2386 (
            .O(N__27137),
            .I(\quad_counter1.b_delay_counter_11 ));
    Odrv4 I__2385 (
            .O(N__27134),
            .I(\quad_counter1.b_delay_counter_11 ));
    InMux I__2384 (
            .O(N__27129),
            .I(\quad_counter1.n19696 ));
    InMux I__2383 (
            .O(N__27126),
            .I(\quad_counter1.n19697 ));
    InMux I__2382 (
            .O(N__27123),
            .I(\quad_counter1.n19698 ));
    InMux I__2381 (
            .O(N__27120),
            .I(\quad_counter1.n19699 ));
    InMux I__2380 (
            .O(N__27117),
            .I(\quad_counter1.n19700 ));
    CEMux I__2379 (
            .O(N__27114),
            .I(N__27110));
    CEMux I__2378 (
            .O(N__27113),
            .I(N__27107));
    LocalMux I__2377 (
            .O(N__27110),
            .I(N__27104));
    LocalMux I__2376 (
            .O(N__27107),
            .I(N__27101));
    Odrv4 I__2375 (
            .O(N__27104),
            .I(n14425));
    Odrv12 I__2374 (
            .O(N__27101),
            .I(n14425));
    SRMux I__2373 (
            .O(N__27096),
            .I(N__27092));
    SRMux I__2372 (
            .O(N__27095),
            .I(N__27089));
    LocalMux I__2371 (
            .O(N__27092),
            .I(N__27086));
    LocalMux I__2370 (
            .O(N__27089),
            .I(N__27083));
    Span4Mux_v I__2369 (
            .O(N__27086),
            .I(N__27077));
    Span4Mux_h I__2368 (
            .O(N__27083),
            .I(N__27077));
    InMux I__2367 (
            .O(N__27082),
            .I(N__27074));
    Odrv4 I__2366 (
            .O(N__27077),
            .I(b_delay_counter_15__N_4140_adj_4773));
    LocalMux I__2365 (
            .O(N__27074),
            .I(b_delay_counter_15__N_4140_adj_4773));
    CascadeMux I__2364 (
            .O(N__27069),
            .I(N__27065));
    InMux I__2363 (
            .O(N__27068),
            .I(N__27062));
    InMux I__2362 (
            .O(N__27065),
            .I(N__27058));
    LocalMux I__2361 (
            .O(N__27062),
            .I(N__27055));
    InMux I__2360 (
            .O(N__27061),
            .I(N__27052));
    LocalMux I__2359 (
            .O(N__27058),
            .I(b_delay_counter_0));
    Odrv4 I__2358 (
            .O(N__27055),
            .I(b_delay_counter_0));
    LocalMux I__2357 (
            .O(N__27052),
            .I(b_delay_counter_0));
    InMux I__2356 (
            .O(N__27045),
            .I(N__27042));
    LocalMux I__2355 (
            .O(N__27042),
            .I(n187));
    InMux I__2354 (
            .O(N__27039),
            .I(bfn_6_10_0_));
    InMux I__2353 (
            .O(N__27036),
            .I(N__27032));
    InMux I__2352 (
            .O(N__27035),
            .I(N__27029));
    LocalMux I__2351 (
            .O(N__27032),
            .I(\quad_counter0.b_delay_counter_1 ));
    LocalMux I__2350 (
            .O(N__27029),
            .I(\quad_counter0.b_delay_counter_1 ));
    InMux I__2349 (
            .O(N__27024),
            .I(\quad_counter0.n19656 ));
    InMux I__2348 (
            .O(N__27021),
            .I(\quad_counter1.n19686 ));
    InMux I__2347 (
            .O(N__27018),
            .I(\quad_counter1.n19687 ));
    InMux I__2346 (
            .O(N__27015),
            .I(N__27011));
    InMux I__2345 (
            .O(N__27014),
            .I(N__27008));
    LocalMux I__2344 (
            .O(N__27011),
            .I(\quad_counter1.b_delay_counter_3 ));
    LocalMux I__2343 (
            .O(N__27008),
            .I(\quad_counter1.b_delay_counter_3 ));
    InMux I__2342 (
            .O(N__27003),
            .I(\quad_counter1.n19688 ));
    CascadeMux I__2341 (
            .O(N__27000),
            .I(N__26996));
    InMux I__2340 (
            .O(N__26999),
            .I(N__26993));
    InMux I__2339 (
            .O(N__26996),
            .I(N__26990));
    LocalMux I__2338 (
            .O(N__26993),
            .I(\quad_counter1.b_delay_counter_4 ));
    LocalMux I__2337 (
            .O(N__26990),
            .I(\quad_counter1.b_delay_counter_4 ));
    InMux I__2336 (
            .O(N__26985),
            .I(\quad_counter1.n19689 ));
    InMux I__2335 (
            .O(N__26982),
            .I(\quad_counter1.n19690 ));
    InMux I__2334 (
            .O(N__26979),
            .I(N__26975));
    InMux I__2333 (
            .O(N__26978),
            .I(N__26972));
    LocalMux I__2332 (
            .O(N__26975),
            .I(\quad_counter1.b_delay_counter_6 ));
    LocalMux I__2331 (
            .O(N__26972),
            .I(\quad_counter1.b_delay_counter_6 ));
    InMux I__2330 (
            .O(N__26967),
            .I(\quad_counter1.n19691 ));
    InMux I__2329 (
            .O(N__26964),
            .I(\quad_counter1.n19692 ));
    CascadeMux I__2328 (
            .O(N__26961),
            .I(N__26958));
    InMux I__2327 (
            .O(N__26958),
            .I(N__26954));
    InMux I__2326 (
            .O(N__26957),
            .I(N__26951));
    LocalMux I__2325 (
            .O(N__26954),
            .I(N__26948));
    LocalMux I__2324 (
            .O(N__26951),
            .I(\quad_counter1.b_delay_counter_8 ));
    Odrv4 I__2323 (
            .O(N__26948),
            .I(\quad_counter1.b_delay_counter_8 ));
    InMux I__2322 (
            .O(N__26943),
            .I(bfn_5_18_0_));
    InMux I__2321 (
            .O(N__26940),
            .I(N__26936));
    InMux I__2320 (
            .O(N__26939),
            .I(N__26933));
    LocalMux I__2319 (
            .O(N__26936),
            .I(N__26930));
    LocalMux I__2318 (
            .O(N__26933),
            .I(\quad_counter1.b_delay_counter_9 ));
    Odrv4 I__2317 (
            .O(N__26930),
            .I(\quad_counter1.b_delay_counter_9 ));
    InMux I__2316 (
            .O(N__26925),
            .I(\quad_counter1.n19694 ));
    CascadeMux I__2315 (
            .O(N__26922),
            .I(\quad_counter0.n27_adj_4756_cascade_ ));
    InMux I__2314 (
            .O(N__26919),
            .I(N__26916));
    LocalMux I__2313 (
            .O(N__26916),
            .I(\quad_counter0.n25_adj_4757 ));
    CascadeMux I__2312 (
            .O(N__26913),
            .I(n9809_cascade_));
    InMux I__2311 (
            .O(N__26910),
            .I(N__26907));
    LocalMux I__2310 (
            .O(N__26907),
            .I(N__26904));
    Odrv12 I__2309 (
            .O(N__26904),
            .I(n9809));
    CascadeMux I__2308 (
            .O(N__26901),
            .I(\quad_counter1.n25_adj_4202_cascade_ ));
    InMux I__2307 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__2306 (
            .O(N__26895),
            .I(N__26892));
    Odrv12 I__2305 (
            .O(N__26892),
            .I(n12940));
    InMux I__2304 (
            .O(N__26889),
            .I(N__26886));
    LocalMux I__2303 (
            .O(N__26886),
            .I(N__26883));
    Span4Mux_v I__2302 (
            .O(N__26883),
            .I(N__26878));
    InMux I__2301 (
            .O(N__26882),
            .I(N__26875));
    InMux I__2300 (
            .O(N__26881),
            .I(N__26872));
    Span4Mux_v I__2299 (
            .O(N__26878),
            .I(N__26866));
    LocalMux I__2298 (
            .O(N__26875),
            .I(N__26866));
    LocalMux I__2297 (
            .O(N__26872),
            .I(N__26863));
    InMux I__2296 (
            .O(N__26871),
            .I(N__26860));
    Span4Mux_v I__2295 (
            .O(N__26866),
            .I(N__26857));
    Span12Mux_v I__2294 (
            .O(N__26863),
            .I(N__26852));
    LocalMux I__2293 (
            .O(N__26860),
            .I(N__26852));
    Span4Mux_v I__2292 (
            .O(N__26857),
            .I(N__26849));
    Span12Mux_v I__2291 (
            .O(N__26852),
            .I(N__26844));
    Sp12to4 I__2290 (
            .O(N__26849),
            .I(N__26844));
    Odrv12 I__2289 (
            .O(N__26844),
            .I(PIN_13_c));
    CascadeMux I__2288 (
            .O(N__26841),
            .I(n12940_cascade_));
    InMux I__2287 (
            .O(N__26838),
            .I(N__26834));
    CascadeMux I__2286 (
            .O(N__26837),
            .I(N__26830));
    LocalMux I__2285 (
            .O(N__26834),
            .I(N__26827));
    InMux I__2284 (
            .O(N__26833),
            .I(N__26824));
    InMux I__2283 (
            .O(N__26830),
            .I(N__26821));
    Span4Mux_v I__2282 (
            .O(N__26827),
            .I(N__26818));
    LocalMux I__2281 (
            .O(N__26824),
            .I(N__26815));
    LocalMux I__2280 (
            .O(N__26821),
            .I(quadB_delayed_adj_4768));
    Odrv4 I__2279 (
            .O(N__26818),
            .I(quadB_delayed_adj_4768));
    Odrv12 I__2278 (
            .O(N__26815),
            .I(quadB_delayed_adj_4768));
    CascadeMux I__2277 (
            .O(N__26808),
            .I(n14425_cascade_));
    InMux I__2276 (
            .O(N__26805),
            .I(N__26802));
    LocalMux I__2275 (
            .O(N__26802),
            .I(\quad_counter1.n26_adj_4200 ));
    InMux I__2274 (
            .O(N__26799),
            .I(N__26794));
    InMux I__2273 (
            .O(N__26798),
            .I(N__26789));
    InMux I__2272 (
            .O(N__26797),
            .I(N__26789));
    LocalMux I__2271 (
            .O(N__26794),
            .I(b_delay_counter_0_adj_4766));
    LocalMux I__2270 (
            .O(N__26789),
            .I(b_delay_counter_0_adj_4766));
    InMux I__2269 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__2268 (
            .O(N__26781),
            .I(n187_adj_4771));
    InMux I__2267 (
            .O(N__26778),
            .I(bfn_5_17_0_));
    CascadeMux I__2266 (
            .O(N__26775),
            .I(\quad_counter0.n25_adj_4760_cascade_ ));
    CascadeMux I__2265 (
            .O(N__26772),
            .I(n12942_cascade_));
    InMux I__2264 (
            .O(N__26769),
            .I(N__26766));
    LocalMux I__2263 (
            .O(N__26766),
            .I(\quad_counter0.n28_adj_4754 ));
    InMux I__2262 (
            .O(N__26763),
            .I(N__26760));
    LocalMux I__2261 (
            .O(N__26760),
            .I(\quad_counter0.n26_adj_4755 ));
    IoInMux I__2260 (
            .O(N__26757),
            .I(N__26754));
    LocalMux I__2259 (
            .O(N__26754),
            .I(tx_enable));
    IoInMux I__2258 (
            .O(N__26751),
            .I(N__26748));
    LocalMux I__2257 (
            .O(N__26748),
            .I(N__26745));
    IoSpan4Mux I__2256 (
            .O(N__26745),
            .I(N__26742));
    Span4Mux_s3_v I__2255 (
            .O(N__26742),
            .I(N__26739));
    Span4Mux_v I__2254 (
            .O(N__26739),
            .I(N__26736));
    Sp12to4 I__2253 (
            .O(N__26736),
            .I(N__26732));
    InMux I__2252 (
            .O(N__26735),
            .I(N__26729));
    Span12Mux_v I__2251 (
            .O(N__26732),
            .I(N__26724));
    LocalMux I__2250 (
            .O(N__26729),
            .I(N__26724));
    Span12Mux_v I__2249 (
            .O(N__26724),
            .I(N__26721));
    Odrv12 I__2248 (
            .O(N__26721),
            .I(LED_c));
    InMux I__2247 (
            .O(N__26718),
            .I(N__26715));
    LocalMux I__2246 (
            .O(N__26715),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__2245 (
            .O(N__26712),
            .I(\quad_counter0.n22_cascade_ ));
    IoInMux I__2244 (
            .O(N__26709),
            .I(N__26706));
    LocalMux I__2243 (
            .O(N__26706),
            .I(N__26703));
    IoSpan4Mux I__2242 (
            .O(N__26703),
            .I(N__26700));
    IoSpan4Mux I__2241 (
            .O(N__26700),
            .I(N__26697));
    IoSpan4Mux I__2240 (
            .O(N__26697),
            .I(N__26694));
    Odrv4 I__2239 (
            .O(N__26694),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\quad_counter1.n19738 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\quad_counter1.n19746 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\quad_counter1.n19754 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\quad_counter1.n19762 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\quad_counter0.n19770 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\quad_counter0.n19778 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\quad_counter0.n19786 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\quad_counter0.n19794 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\quad_counter1.n19693 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\quad_counter1.n19708 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(\quad_counter0.n19663 ),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(\quad_counter0.n19678 ),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\c0.tx.n19730 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_11_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_26_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_19_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_1_0_));
    defparam IN_MUX_bfv_19_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_2_0_ (
            .carryinitin(\c0.n19625_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_2_0_));
    defparam IN_MUX_bfv_19_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_3_0_ (
            .carryinitin(\c0.n19626_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_3_0_));
    defparam IN_MUX_bfv_19_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_4_0_ (
            .carryinitin(\c0.n19627_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_4_0_));
    defparam IN_MUX_bfv_19_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_5_0_ (
            .carryinitin(\c0.n19628_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_5_0_));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(\c0.n19629_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(\c0.n19630_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\c0.n19631_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_19_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_9_0_ (
            .carryinitin(\c0.n19632_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_9_0_));
    defparam IN_MUX_bfv_19_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_10_0_ (
            .carryinitin(\c0.n19633_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_10_0_));
    defparam IN_MUX_bfv_19_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_11_0_ (
            .carryinitin(\c0.n19634_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_11_0_));
    defparam IN_MUX_bfv_19_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_12_0_ (
            .carryinitin(\c0.n19635_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_12_0_));
    defparam IN_MUX_bfv_19_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_13_0_ (
            .carryinitin(\c0.n19636_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_13_0_));
    defparam IN_MUX_bfv_19_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_14_0_ (
            .carryinitin(\c0.n19637_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_14_0_));
    defparam IN_MUX_bfv_19_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_15_0_ (
            .carryinitin(\c0.n19638_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_15_0_));
    defparam IN_MUX_bfv_19_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_16_0_ (
            .carryinitin(\c0.n19639_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_16_0_));
    defparam IN_MUX_bfv_19_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_17_0_ (
            .carryinitin(\c0.n19640_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_17_0_));
    defparam IN_MUX_bfv_19_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_18_0_ (
            .carryinitin(\c0.n19641_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_18_0_));
    defparam IN_MUX_bfv_19_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_19_0_ (
            .carryinitin(\c0.n19642_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_19_0_));
    defparam IN_MUX_bfv_19_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_20_0_ (
            .carryinitin(\c0.n19643_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_20_0_));
    defparam IN_MUX_bfv_19_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_21_0_ (
            .carryinitin(\c0.n19644_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_21_0_));
    defparam IN_MUX_bfv_19_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_22_0_ (
            .carryinitin(\c0.n19645_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_22_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(\c0.n19646_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_19_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_24_0_ (
            .carryinitin(\c0.n19647_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_24_0_));
    defparam IN_MUX_bfv_19_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_25_0_ (
            .carryinitin(\c0.n19648_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_25_0_));
    defparam IN_MUX_bfv_19_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_26_0_ (
            .carryinitin(\c0.n19649_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_26_0_));
    defparam IN_MUX_bfv_19_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_27_0_ (
            .carryinitin(\c0.n19650_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_27_0_));
    defparam IN_MUX_bfv_19_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_28_0_ (
            .carryinitin(\c0.n19651_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_28_0_));
    defparam IN_MUX_bfv_19_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_29_0_ (
            .carryinitin(\c0.n19652_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_29_0_));
    defparam IN_MUX_bfv_19_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_30_0_ (
            .carryinitin(\c0.n19653_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_30_0_));
    defparam IN_MUX_bfv_19_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_31_0_ (
            .carryinitin(\c0.n19654_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_31_0_));
    defparam IN_MUX_bfv_19_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_32_0_ (
            .carryinitin(\c0.n19655_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_19_32_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__26709),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_4_5 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28592),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_R_49_LC_3_16_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_49_LC_3_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_49_LC_3_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_R_49_LC_3_16_6  (
            .in0(N__26735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_Rx_Data_R ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78562),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_delayed_62_LC_4_12_3 .C_ON=1'b0;
    defparam \quad_counter1.quadB_delayed_62_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadB_delayed_62_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.quadB_delayed_62_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26871),
            .lcout(quadB_delayed_adj_4768),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78571),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadB_delayed_62_LC_4_13_0 .C_ON=1'b0;
    defparam \quad_counter0.quadB_delayed_62_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadB_delayed_62_LC_4_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.quadB_delayed_62_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27411),
            .lcout(quadB_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78569),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_4_16_3 .C_ON=1'b0;
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_4_16_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.quadB_I_0_79_2_lut_LC_4_16_3  (
            .in0(N__26881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26833),
            .lcout(b_delay_counter_15__N_4140_adj_4773),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_4_16_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_4_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26718),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78564),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i0_LC_5_10_1 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i0_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i0_LC_5_10_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \quad_counter0.b_delay_counter__i0_LC_5_10_1  (
            .in0(N__27448),
            .in1(N__27045),
            .in2(N__27069),
            .in3(N__27469),
            .lcout(b_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78592),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_65_LC_5_11_2 .C_ON=1'b0;
    defparam \quad_counter1.B_65_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_65_LC_5_11_2 .LUT_INIT=16'b1010101011101000;
    LogicCell40 \quad_counter1.B_65_LC_5_11_2  (
            .in0(N__29891),
            .in1(N__26882),
            .in2(N__26837),
            .in3(N__26898),
            .lcout(B_filtered_adj_4764),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78584),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_LC_5_11_3 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_LC_5_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_LC_5_11_3  (
            .in0(N__27236),
            .in1(N__27221),
            .in2(N__27204),
            .in3(N__27179),
            .lcout(),
            .ltout(\quad_counter0.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_3_lut_LC_5_11_4 .C_ON=1'b0;
    defparam \quad_counter0.i11_3_lut_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_3_lut_LC_5_11_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter0.i11_3_lut_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__27035),
            .in2(N__26712),
            .in3(N__27503),
            .lcout(),
            .ltout(\quad_counter0.n25_adj_4760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_4_lut_LC_5_11_5 .C_ON=1'b0;
    defparam \quad_counter0.i2_4_lut_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_4_lut_LC_5_11_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \quad_counter0.i2_4_lut_LC_5_11_5  (
            .in0(N__27068),
            .in1(N__27251),
            .in2(N__26775),
            .in3(N__27642),
            .lcout(n12942),
            .ltout(n12942_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_5_11_6.C_ON=1'b0;
    defparam i1_4_lut_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_5_11_6.LUT_INIT=16'b1110110011011100;
    LogicCell40 i1_4_lut_LC_5_11_6 (
            .in0(N__27417),
            .in1(N__27438),
            .in2(N__26772),
            .in3(N__27368),
            .lcout(n14315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadB_I_0_79_2_lut_LC_5_12_2 .C_ON=1'b0;
    defparam \quad_counter0.quadB_I_0_79_2_lut_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadB_I_0_79_2_lut_LC_5_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.quadB_I_0_79_2_lut_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__27412),
            .in2(_gnd_net_),
            .in3(N__27361),
            .lcout(b_delay_counter_15__N_4140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_LC_5_13_0 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_LC_5_13_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter0.i9_4_lut_LC_5_13_0  (
            .in0(N__27542),
            .in1(N__27734),
            .in2(N__27561),
            .in3(N__27634),
            .lcout(\quad_counter0.n25_adj_4757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_LC_5_13_2 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_LC_5_13_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter0.i12_4_lut_LC_5_13_2  (
            .in0(N__27575),
            .in1(N__27782),
            .in2(N__27594),
            .in3(N__27608),
            .lcout(\quad_counter0.n28_adj_4754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_delayed_67_LC_5_13_5 .C_ON=1'b0;
    defparam \quad_counter0.A_delayed_67_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_delayed_67_LC_5_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.A_delayed_67_LC_5_13_5  (
            .in0(N__28133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78572),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i0_LC_5_13_6 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i0_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i0_LC_5_13_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \quad_counter0.a_delay_counter__i0_LC_5_13_6  (
            .in0(N__28007),
            .in1(N__27621),
            .in2(N__28029),
            .in3(N__27635),
            .lcout(a_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78572),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_LC_5_14_0 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_LC_5_14_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_LC_5_14_0  (
            .in0(N__27719),
            .in1(N__27704),
            .in2(N__27528),
            .in3(N__27767),
            .lcout(\quad_counter0.n26_adj_4755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_LC_5_14_1 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_LC_5_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_LC_5_14_1  (
            .in0(N__27689),
            .in1(N__27797),
            .in2(N__27753),
            .in3(N__28040),
            .lcout(),
            .ltout(\quad_counter0.n27_adj_4756_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_LC_5_14_2 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_LC_5_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_LC_5_14_2  (
            .in0(N__26769),
            .in1(N__26763),
            .in2(N__26922),
            .in3(N__26919),
            .lcout(n9809),
            .ltout(n9809_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_2055_LC_5_14_3.C_ON=1'b0;
    defparam i1_3_lut_adj_2055_LC_5_14_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_2055_LC_5_14_3.LUT_INIT=16'b1111010111111010;
    LogicCell40 i1_3_lut_adj_2055_LC_5_14_3 (
            .in0(N__27920),
            .in1(_gnd_net_),
            .in2(N__26913),
            .in3(N__27882),
            .lcout(n14469),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_63_LC_5_16_0 .C_ON=1'b0;
    defparam \quad_counter0.A_63_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_63_LC_5_16_0 .LUT_INIT=16'b1111111001000000;
    LogicCell40 \quad_counter0.A_63_LC_5_16_0  (
            .in0(N__26910),
            .in1(N__27909),
            .in2(N__27881),
            .in3(N__28134),
            .lcout(A_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1164_LC_5_16_1 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1164_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1164_LC_5_16_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1164_LC_5_16_1  (
            .in0(N__26940),
            .in1(N__27014),
            .in2(N__27000),
            .in3(N__26797),
            .lcout(),
            .ltout(\quad_counter1.n25_adj_4202_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_adj_1165_LC_5_16_2 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_adj_1165_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_adj_1165_LC_5_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_adj_1165_LC_5_16_2  (
            .in0(N__27930),
            .in1(N__26805),
            .in2(N__26901),
            .in3(N__27804),
            .lcout(n12940),
            .ltout(n12940_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_2054_LC_5_16_3.C_ON=1'b0;
    defparam i1_3_lut_adj_2054_LC_5_16_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_2054_LC_5_16_3.LUT_INIT=16'b1111001111111100;
    LogicCell40 i1_3_lut_adj_2054_LC_5_16_3 (
            .in0(_gnd_net_),
            .in1(N__26889),
            .in2(N__26841),
            .in3(N__26838),
            .lcout(n14425),
            .ltout(n14425_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i0_LC_5_16_4 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i0_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i0_LC_5_16_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \quad_counter1.b_delay_counter__i0_LC_5_16_4  (
            .in0(N__26798),
            .in1(N__26784),
            .in2(N__26808),
            .in3(N__27082),
            .lcout(b_delay_counter_0_adj_4766),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1162_LC_5_16_5 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1162_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1162_LC_5_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1162_LC_5_16_5  (
            .in0(N__27144),
            .in1(N__27162),
            .in2(N__26961),
            .in3(N__26978),
            .lcout(\quad_counter1.n26_adj_4200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_86_2_lut_LC_5_17_0 .C_ON=1'b1;
    defparam \quad_counter1.add_86_2_lut_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_86_2_lut_LC_5_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_86_2_lut_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__26799),
            .in2(_gnd_net_),
            .in3(N__26778),
            .lcout(n187_adj_4771),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\quad_counter1.n19686 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i1_LC_5_17_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i1_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i1_LC_5_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i1_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__27969),
            .in2(_gnd_net_),
            .in3(N__27021),
            .lcout(\quad_counter1.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n19686 ),
            .carryout(\quad_counter1.n19687 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i2_LC_5_17_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i2_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i2_LC_5_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i2_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__27956),
            .in2(_gnd_net_),
            .in3(N__27018),
            .lcout(\quad_counter1.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n19687 ),
            .carryout(\quad_counter1.n19688 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i3_LC_5_17_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i3_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i3_LC_5_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i3_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__27015),
            .in2(_gnd_net_),
            .in3(N__27003),
            .lcout(\quad_counter1.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n19688 ),
            .carryout(\quad_counter1.n19689 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i4_LC_5_17_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i4_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i4_LC_5_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i4_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__26999),
            .in2(_gnd_net_),
            .in3(N__26985),
            .lcout(\quad_counter1.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n19689 ),
            .carryout(\quad_counter1.n19690 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i5_LC_5_17_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i5_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i5_LC_5_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i5_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__27942),
            .in2(_gnd_net_),
            .in3(N__26982),
            .lcout(\quad_counter1.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n19690 ),
            .carryout(\quad_counter1.n19691 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i6_LC_5_17_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i6_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i6_LC_5_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i6_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__26979),
            .in2(_gnd_net_),
            .in3(N__26967),
            .lcout(\quad_counter1.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n19691 ),
            .carryout(\quad_counter1.n19692 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i7_LC_5_17_7 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i7_LC_5_17_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i7_LC_5_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i7_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__27843),
            .in2(_gnd_net_),
            .in3(N__26964),
            .lcout(\quad_counter1.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n19692 ),
            .carryout(\quad_counter1.n19693 ),
            .clk(N__78563),
            .ce(N__27114),
            .sr(N__27095));
    defparam \quad_counter1.b_delay_counter__i8_LC_5_18_0 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i8_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i8_LC_5_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i8_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__26957),
            .in2(_gnd_net_),
            .in3(N__26943),
            .lcout(\quad_counter1.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\quad_counter1.n19694 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i9_LC_5_18_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i9_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i9_LC_5_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i9_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__26939),
            .in2(_gnd_net_),
            .in3(N__26925),
            .lcout(\quad_counter1.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n19694 ),
            .carryout(\quad_counter1.n19695 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i10_LC_5_18_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i10_LC_5_18_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i10_LC_5_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i10_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__27161),
            .in2(_gnd_net_),
            .in3(N__27147),
            .lcout(\quad_counter1.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n19695 ),
            .carryout(\quad_counter1.n19696 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i11_LC_5_18_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i11_LC_5_18_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i11_LC_5_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i11_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__27143),
            .in2(_gnd_net_),
            .in3(N__27129),
            .lcout(\quad_counter1.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n19696 ),
            .carryout(\quad_counter1.n19697 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i12_LC_5_18_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i12_LC_5_18_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i12_LC_5_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i12_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(N__27830),
            .in2(_gnd_net_),
            .in3(N__27126),
            .lcout(\quad_counter1.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n19697 ),
            .carryout(\quad_counter1.n19698 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i13_LC_5_18_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i13_LC_5_18_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i13_LC_5_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i13_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(N__27983),
            .in2(_gnd_net_),
            .in3(N__27123),
            .lcout(\quad_counter1.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n19698 ),
            .carryout(\quad_counter1.n19699 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i14_LC_5_18_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i14_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i14_LC_5_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i14_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(N__27855),
            .in2(_gnd_net_),
            .in3(N__27120),
            .lcout(\quad_counter1.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n19699 ),
            .carryout(\quad_counter1.n19700 ),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter1.b_delay_counter__i15_LC_5_18_7 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i15_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i15_LC_5_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i15_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(N__27816),
            .in2(_gnd_net_),
            .in3(N__27117),
            .lcout(\quad_counter1.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78566),
            .ce(N__27113),
            .sr(N__27096));
    defparam \quad_counter0.add_86_2_lut_LC_6_10_0 .C_ON=1'b1;
    defparam \quad_counter0.add_86_2_lut_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_2_lut_LC_6_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_86_2_lut_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__27061),
            .in2(_gnd_net_),
            .in3(N__27039),
            .lcout(n187),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\quad_counter0.n19656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i1_LC_6_10_1 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i1_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i1_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__27036),
            .in2(_gnd_net_),
            .in3(N__27024),
            .lcout(\quad_counter0.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n19656 ),
            .carryout(\quad_counter0.n19657 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i2_LC_6_10_2 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i2_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i2_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i2_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__27252),
            .in2(_gnd_net_),
            .in3(N__27240),
            .lcout(\quad_counter0.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n19657 ),
            .carryout(\quad_counter0.n19658 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i3_LC_6_10_3 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i3_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i3_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i3_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__27237),
            .in2(_gnd_net_),
            .in3(N__27225),
            .lcout(\quad_counter0.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n19658 ),
            .carryout(\quad_counter0.n19659 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i4_LC_6_10_4 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i4_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i4_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i4_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__27222),
            .in2(_gnd_net_),
            .in3(N__27210),
            .lcout(\quad_counter0.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n19659 ),
            .carryout(\quad_counter0.n19660 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i5_LC_6_10_5 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i5_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i5_LC_6_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i5_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__27278),
            .in2(_gnd_net_),
            .in3(N__27207),
            .lcout(\quad_counter0.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n19660 ),
            .carryout(\quad_counter0.n19661 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i6_LC_6_10_6 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i6_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i6_LC_6_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i6_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__27203),
            .in2(_gnd_net_),
            .in3(N__27189),
            .lcout(\quad_counter0.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n19661 ),
            .carryout(\quad_counter0.n19662 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i7_LC_6_10_7 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i7_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i7_LC_6_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i7_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(N__27308),
            .in2(_gnd_net_),
            .in3(N__27186),
            .lcout(\quad_counter0.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n19662 ),
            .carryout(\quad_counter0.n19663 ),
            .clk(N__78602),
            .ce(N__27483),
            .sr(N__27452));
    defparam \quad_counter0.b_delay_counter__i8_LC_6_11_0 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i8_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i8_LC_6_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i8_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__27327),
            .in2(_gnd_net_),
            .in3(N__27183),
            .lcout(\quad_counter0.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\quad_counter0.n19664 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i9_LC_6_11_1 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i9_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i9_LC_6_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i9_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__27180),
            .in2(_gnd_net_),
            .in3(N__27168),
            .lcout(\quad_counter0.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n19664 ),
            .carryout(\quad_counter0.n19665 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i10_LC_6_11_2 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i10_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i10_LC_6_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i10_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__27675),
            .in2(_gnd_net_),
            .in3(N__27165),
            .lcout(\quad_counter0.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n19665 ),
            .carryout(\quad_counter0.n19666 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i11_LC_6_11_3 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i11_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i11_LC_6_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i11_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__27663),
            .in2(_gnd_net_),
            .in3(N__27510),
            .lcout(\quad_counter0.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n19666 ),
            .carryout(\quad_counter0.n19667 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i12_LC_6_11_4 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i12_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i12_LC_6_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i12_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__27294),
            .in2(_gnd_net_),
            .in3(N__27507),
            .lcout(\quad_counter0.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n19667 ),
            .carryout(\quad_counter0.n19668 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i13_LC_6_11_5 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i13_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i13_LC_6_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i13_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__27504),
            .in2(_gnd_net_),
            .in3(N__27492),
            .lcout(\quad_counter0.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n19668 ),
            .carryout(\quad_counter0.n19669 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i14_LC_6_11_6 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i14_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i14_LC_6_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i14_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__27264),
            .in2(_gnd_net_),
            .in3(N__27489),
            .lcout(\quad_counter0.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n19669 ),
            .carryout(\quad_counter0.n19670 ),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.b_delay_counter__i15_LC_6_11_7 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i15_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i15_LC_6_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i15_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__27339),
            .in2(_gnd_net_),
            .in3(N__27486),
            .lcout(\quad_counter0.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78593),
            .ce(N__27482),
            .sr(N__27453));
    defparam \quad_counter0.B_65_LC_6_12_0 .C_ON=1'b0;
    defparam \quad_counter0.B_65_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_65_LC_6_12_0 .LUT_INIT=16'b1111000011101000;
    LogicCell40 \quad_counter0.B_65_LC_6_12_0  (
            .in0(N__27416),
            .in1(N__27372),
            .in2(N__28092),
            .in3(N__27345),
            .lcout(B_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78585),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_2_lut_LC_6_12_2 .C_ON=1'b0;
    defparam \quad_counter0.i4_2_lut_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_2_lut_LC_6_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i4_2_lut_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__27338),
            .in2(_gnd_net_),
            .in3(N__27326),
            .lcout(\quad_counter0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_LC_6_12_3 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_LC_6_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter0.i3_4_lut_LC_6_12_3  (
            .in0(N__28064),
            .in1(N__28137),
            .in2(N__28090),
            .in3(N__27315),
            .lcout(count_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_2052_LC_6_12_4 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_2052_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_2052_LC_6_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_2052_LC_6_12_4  (
            .in0(N__27309),
            .in1(N__27293),
            .in2(N__27282),
            .in3(N__27263),
            .lcout(),
            .ltout(\quad_counter0.n24_adj_4758_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_2053_LC_6_12_5 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_2053_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_2053_LC_6_12_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i12_4_lut_adj_2053_LC_6_12_5  (
            .in0(N__27674),
            .in1(N__27662),
            .in2(N__27651),
            .in3(N__27648),
            .lcout(\quad_counter0.n26_adj_4759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_85_2_lut_LC_6_13_0 .C_ON=1'b1;
    defparam \quad_counter0.add_85_2_lut_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_85_2_lut_LC_6_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_85_2_lut_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__27636),
            .in2(_gnd_net_),
            .in3(N__27612),
            .lcout(n39),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\quad_counter0.n19671 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i1_LC_6_13_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i1_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i1_LC_6_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i1_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__27609),
            .in2(_gnd_net_),
            .in3(N__27597),
            .lcout(\quad_counter0.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n19671 ),
            .carryout(\quad_counter0.n19672 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i2_LC_6_13_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i2_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i2_LC_6_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i2_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(N__27593),
            .in2(_gnd_net_),
            .in3(N__27579),
            .lcout(\quad_counter0.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n19672 ),
            .carryout(\quad_counter0.n19673 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i3_LC_6_13_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i3_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i3_LC_6_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i3_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__27576),
            .in2(_gnd_net_),
            .in3(N__27564),
            .lcout(\quad_counter0.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n19673 ),
            .carryout(\quad_counter0.n19674 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i4_LC_6_13_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i4_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i4_LC_6_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i4_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(N__27560),
            .in2(_gnd_net_),
            .in3(N__27546),
            .lcout(\quad_counter0.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n19674 ),
            .carryout(\quad_counter0.n19675 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i5_LC_6_13_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i5_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i5_LC_6_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i5_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(N__27543),
            .in2(_gnd_net_),
            .in3(N__27531),
            .lcout(\quad_counter0.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n19675 ),
            .carryout(\quad_counter0.n19676 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i6_LC_6_13_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i6_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i6_LC_6_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i6_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__27527),
            .in2(_gnd_net_),
            .in3(N__27513),
            .lcout(\quad_counter0.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n19676 ),
            .carryout(\quad_counter0.n19677 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i7_LC_6_13_7 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i7_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i7_LC_6_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i7_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__27798),
            .in2(_gnd_net_),
            .in3(N__27786),
            .lcout(\quad_counter0.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n19677 ),
            .carryout(\quad_counter0.n19678 ),
            .clk(N__78576),
            .ce(N__28025),
            .sr(N__28008));
    defparam \quad_counter0.a_delay_counter__i8_LC_6_14_0 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i8_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i8_LC_6_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i8_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__27783),
            .in2(_gnd_net_),
            .in3(N__27771),
            .lcout(\quad_counter0.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\quad_counter0.n19679 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i9_LC_6_14_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i9_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i9_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i9_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__27768),
            .in2(_gnd_net_),
            .in3(N__27756),
            .lcout(\quad_counter0.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n19679 ),
            .carryout(\quad_counter0.n19680 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i10_LC_6_14_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i10_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i10_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i10_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__27752),
            .in2(_gnd_net_),
            .in3(N__27738),
            .lcout(\quad_counter0.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n19680 ),
            .carryout(\quad_counter0.n19681 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i11_LC_6_14_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i11_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i11_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i11_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__27735),
            .in2(_gnd_net_),
            .in3(N__27723),
            .lcout(\quad_counter0.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n19681 ),
            .carryout(\quad_counter0.n19682 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i12_LC_6_14_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i12_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i12_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i12_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__27720),
            .in2(_gnd_net_),
            .in3(N__27708),
            .lcout(\quad_counter0.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n19682 ),
            .carryout(\quad_counter0.n19683 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i13_LC_6_14_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i13_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i13_LC_6_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i13_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(N__27705),
            .in2(_gnd_net_),
            .in3(N__27693),
            .lcout(\quad_counter0.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n19683 ),
            .carryout(\quad_counter0.n19684 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i14_LC_6_14_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i14_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i14_LC_6_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i14_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__27690),
            .in2(_gnd_net_),
            .in3(N__27678),
            .lcout(\quad_counter0.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n19684 ),
            .carryout(\quad_counter0.n19685 ),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.a_delay_counter__i15_LC_6_14_7 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i15_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i15_LC_6_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i15_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(N__28041),
            .in2(_gnd_net_),
            .in3(N__28044),
            .lcout(\quad_counter0.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78573),
            .ce(N__28024),
            .sr(N__28003));
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_6_15_4 .C_ON=1'b0;
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_6_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.quadA_I_0_73_2_lut_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__27921),
            .in2(_gnd_net_),
            .in3(N__27871),
            .lcout(a_delay_counter_15__N_4123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i21282_1_lut_LC_6_16_1 .C_ON=1'b0;
    defparam \c0.tx.i21282_1_lut_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i21282_1_lut_LC_6_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.i21282_1_lut_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28951),
            .lcout(\c0.tx.n25051 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1161_LC_6_16_4 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1161_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1161_LC_6_16_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1161_LC_6_16_4  (
            .in0(N__27984),
            .in1(N__27968),
            .in2(N__27957),
            .in3(N__27941),
            .lcout(\quad_counter1.n28_adj_4199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadA_delayed_61_LC_6_16_6 .C_ON=1'b0;
    defparam \quad_counter0.quadA_delayed_61_LC_6_16_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadA_delayed_61_LC_6_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.quadA_delayed_61_LC_6_16_6  (
            .in0(N__27919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadA_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78567),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1163_LC_6_17_6 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1163_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1163_LC_6_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1163_LC_6_17_6  (
            .in0(N__27854),
            .in1(N__27842),
            .in2(N__27831),
            .in3(N__27815),
            .lcout(\quad_counter1.n27_adj_4201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i13_LC_6_18_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_6_18_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_6_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_6_18_5  (
            .in0(_gnd_net_),
            .in1(N__29494),
            .in2(_gnd_net_),
            .in3(N__48978),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78568),
            .ce(),
            .sr(N__29472));
    defparam \c0.rx.n25068_bdd_4_lut_4_lut_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.rx.n25068_bdd_4_lut_4_lut_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.n25068_bdd_4_lut_4_lut_LC_6_21_6 .LUT_INIT=16'b1111110000000101;
    LogicCell40 \c0.rx.n25068_bdd_4_lut_4_lut_LC_6_21_6  (
            .in0(N__50825),
            .in1(N__39315),
            .in2(N__50177),
            .in3(N__28284),
            .lcout(n25071),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_7_11_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_7_11_0 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_7_11_0  (
            .in0(N__28101),
            .in1(N__38463),
            .in2(N__28686),
            .in3(N__28374),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78603),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1074_1_lut_2_lut_LC_7_12_0 .C_ON=1'b0;
    defparam \quad_counter0.i1074_1_lut_2_lut_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1074_1_lut_2_lut_LC_7_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter0.i1074_1_lut_2_lut_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__28060),
            .in2(_gnd_net_),
            .in3(N__28135),
            .lcout(\quad_counter0.n2313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_7_12_1 .C_ON=1'b0;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_7_12_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \quad_counter0.A_filtered_I_0_2_lut_LC_7_12_1  (
            .in0(N__28136),
            .in1(_gnd_net_),
            .in2(N__28065),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5179_4_lut_LC_7_12_3 .C_ON=1'b0;
    defparam \c0.tx.i5179_4_lut_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5179_4_lut_LC_7_12_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.tx.i5179_4_lut_LC_7_12_3  (
            .in0(N__29246),
            .in1(N__30577),
            .in2(N__28449),
            .in3(N__28372),
            .lcout(n8628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_7_12_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_7_12_5 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_7_12_5  (
            .in0(N__29247),
            .in1(N__28757),
            .in2(_gnd_net_),
            .in3(N__28539),
            .lcout(\c0.tx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_4_lut_LC_7_12_6 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_4_lut_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_4_lut_LC_7_12_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i2_3_lut_4_lut_LC_7_12_6  (
            .in0(N__28418),
            .in1(N__29245),
            .in2(N__30582),
            .in3(N__28666),
            .lcout(n9603),
            .ltout(n9603_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_7_12_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_7_12_7 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_7_12_7  (
            .in0(N__28559),
            .in1(N__30131),
            .in2(N__28095),
            .in3(N__28173),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__3__5450_LC_7_13_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__3__5450_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__3__5450_LC_7_13_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_9__3__5450_LC_7_13_4  (
            .in0(N__47994),
            .in1(N__46098),
            .in2(N__44781),
            .in3(N__28161),
            .lcout(data_out_frame_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5_1_lut_LC_7_14_1 .C_ON=1'b0;
    defparam \c0.tx.i5_1_lut_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5_1_lut_LC_7_14_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \c0.tx.i5_1_lut_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__28410),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n14374),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.B_delayed_68_LC_7_14_2 .C_ON=1'b0;
    defparam \quad_counter0.B_delayed_68_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_delayed_68_LC_7_14_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \quad_counter0.B_delayed_68_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__28091),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78577),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2062_LC_7_14_3.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2062_LC_7_14_3.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2062_LC_7_14_3.LUT_INIT=16'b1111110100001000;
    LogicCell40 i24_3_lut_4_lut_adj_2062_LC_7_14_3 (
            .in0(N__31197),
            .in1(N__28215),
            .in2(N__31329),
            .in3(N__28611),
            .lcout(n10_adj_4777),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21318_LC_7_14_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21318_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21318_LC_7_14_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_21318_LC_7_14_4  (
            .in0(N__30966),
            .in1(N__40816),
            .in2(N__30711),
            .in3(N__43219),
            .lcout(),
            .ltout(\c0.n25086_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25086_bdd_4_lut_LC_7_14_5 .C_ON=1'b0;
    defparam \c0.n25086_bdd_4_lut_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.n25086_bdd_4_lut_LC_7_14_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n25086_bdd_4_lut_LC_7_14_5  (
            .in0(N__40817),
            .in1(N__30003),
            .in2(N__28164),
            .in3(N__28160),
            .lcout(\c0.n25089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21035_4_lut_LC_7_14_6 .C_ON=1'b0;
    defparam \c0.i21035_4_lut_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i21035_4_lut_LC_7_14_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \c0.i21035_4_lut_LC_7_14_6  (
            .in0(N__32151),
            .in1(N__31323),
            .in2(N__31417),
            .in3(N__28197),
            .lcout(),
            .ltout(n24802_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2064_LC_7_14_7.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2064_LC_7_14_7.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2064_LC_7_14_7.LUT_INIT=16'b1111010010110000;
    LogicCell40 i24_3_lut_4_lut_adj_2064_LC_7_14_7 (
            .in0(N__31324),
            .in1(N__31198),
            .in2(N__28149),
            .in3(N__28143),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_7_15_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_7_15_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_7_15_0  (
            .in0(N__29241),
            .in1(N__28414),
            .in2(N__28683),
            .in3(N__28357),
            .lcout(\c0.tx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_7_15_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_7_15_3 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_7_15_3  (
            .in0(N__28508),
            .in1(N__28890),
            .in2(N__30146),
            .in3(N__30213),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_7_15_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_7_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_7_15_5  (
            .in0(N__30258),
            .in1(N__34935),
            .in2(_gnd_net_),
            .in3(N__43239),
            .lcout(),
            .ltout(\c0.n11_adj_4715_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21242_4_lut_LC_7_15_6 .C_ON=1'b0;
    defparam \c0.i21242_4_lut_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i21242_4_lut_LC_7_15_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.i21242_4_lut_LC_7_15_6  (
            .in0(N__40820),
            .in1(N__28260),
            .in2(N__28146),
            .in3(N__41046),
            .lcout(n25010),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_3_lut_3_lut_LC_7_16_0 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_3_lut_3_lut_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_3_lut_3_lut_LC_7_16_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.tx.i2_2_lut_3_lut_3_lut_LC_7_16_0  (
            .in0(N__28405),
            .in1(N__29240),
            .in2(_gnd_net_),
            .in3(N__28876),
            .lcout(),
            .ltout(\c0.tx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i21285_4_lut_LC_7_16_1 .C_ON=1'b0;
    defparam \c0.tx.i21285_4_lut_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i21285_4_lut_LC_7_16_1 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \c0.tx.i21285_4_lut_LC_7_16_1  (
            .in0(N__28406),
            .in1(N__28188),
            .in2(N__28227),
            .in3(N__28206),
            .lcout(\c0.tx.n17199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21249_4_lut_LC_7_16_2 .C_ON=1'b0;
    defparam \c0.i21249_4_lut_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21249_4_lut_LC_7_16_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i21249_4_lut_LC_7_16_2  (
            .in0(N__28224),
            .in1(N__40819),
            .in2(N__29154),
            .in3(N__41045),
            .lcout(n25018),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_LC_7_16_4 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_LC_7_16_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx.i2_4_lut_LC_7_16_4  (
            .in0(N__28669),
            .in1(N__29239),
            .in2(N__29004),
            .in3(N__28875),
            .lcout(\c0.tx.n23980 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_7_16_7 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_7_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.tx.i1_2_lut_LC_7_16_7  (
            .in0(N__28877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29003),
            .lcout(r_SM_Main_2_N_3751_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_7_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_7_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_7_17_0  (
            .in0(N__30339),
            .in1(N__28920),
            .in2(_gnd_net_),
            .in3(N__43181),
            .lcout(),
            .ltout(\c0.n5_adj_4712_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21033_4_lut_LC_7_17_1 .C_ON=1'b0;
    defparam \c0.i21033_4_lut_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21033_4_lut_LC_7_17_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.i21033_4_lut_LC_7_17_1  (
            .in0(N__28179),
            .in1(N__40818),
            .in2(N__28200),
            .in3(N__41034),
            .lcout(\c0.n24800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_7_17_5 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_7_17_5 .LUT_INIT=16'b0010010100000101;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_7_17_5  (
            .in0(N__50035),
            .in1(N__49941),
            .in2(N__50178),
            .in3(N__42027),
            .lcout(\c0.rx.n14277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_LC_7_18_3 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \c0.tx.i1_3_lut_LC_7_18_3  (
            .in0(N__28998),
            .in1(N__29220),
            .in2(_gnd_net_),
            .in3(N__28667),
            .lcout(\c0.tx.n5_adj_4207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21182_3_lut_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.i21182_3_lut_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21182_3_lut_LC_7_18_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i21182_3_lut_LC_7_18_4  (
            .in0(N__28251),
            .in1(N__41026),
            .in2(_gnd_net_),
            .in3(N__43171),
            .lcout(\c0.n24949 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21204_2_lut_4_lut_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.rx.i21204_2_lut_4_lut_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21204_2_lut_4_lut_LC_7_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i21204_2_lut_4_lut_LC_7_18_5  (
            .in0(N__49685),
            .in1(N__49656),
            .in2(N__47232),
            .in3(N__42018),
            .lcout(\c0.rx.n24875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i14334_2_lut_3_lut_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.tx.i14334_2_lut_3_lut_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i14334_2_lut_3_lut_LC_7_18_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.tx.i14334_2_lut_3_lut_LC_7_18_6  (
            .in0(N__28668),
            .in1(N__28999),
            .in2(_gnd_net_),
            .in3(N__28878),
            .lcout(n17951),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1859_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1859_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1859_LC_7_19_1 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i2_3_lut_adj_1859_LC_7_19_1  (
            .in0(N__40780),
            .in1(N__31177),
            .in2(_gnd_net_),
            .in3(N__41025),
            .lcout(n24682),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21333_LC_7_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21333_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21333_LC_7_19_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_21333_LC_7_19_2  (
            .in0(N__30240),
            .in1(N__40779),
            .in2(N__35166),
            .in3(N__43180),
            .lcout(),
            .ltout(\c0.n25104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25104_bdd_4_lut_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.n25104_bdd_4_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.n25104_bdd_4_lut_LC_7_19_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n25104_bdd_4_lut_LC_7_19_3  (
            .in0(N__40781),
            .in1(N__29109),
            .in2(N__28263),
            .in3(N__28308),
            .lcout(\c0.n25107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__7__5478_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__7__5478_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__7__5478_LC_7_20_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__7__5478_LC_7_20_6  (
            .in0(N__48067),
            .in1(N__46084),
            .in2(N__42618),
            .in3(N__28250),
            .lcout(data_out_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78578),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_7_21_0 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_7_21_0  (
            .in0(N__28236),
            .in1(N__49956),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1940_2_lut_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.rx.i1940_2_lut_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1940_2_lut_LC_7_21_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i1940_2_lut_LC_7_21_1  (
            .in0(N__47233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49658),
            .lcout(),
            .ltout(n3821_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_7_21_2 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_7_21_2  (
            .in0(N__49684),
            .in1(N__47103),
            .in2(N__28230),
            .in3(N__47150),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__7__5446_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__7__5446_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__7__5446_LC_7_21_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_9__7__5446_LC_7_21_4  (
            .in0(N__48068),
            .in1(N__45945),
            .in2(N__36711),
            .in3(N__28307),
            .lcout(data_out_frame_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_21_7 .LUT_INIT=16'b0111101000101010;
    LogicCell40 \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_21_7  (
            .in0(N__50000),
            .in1(N__42022),
            .in2(N__50162),
            .in3(N__28293),
            .lcout(\c0.rx.n25068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i26_LC_7_22_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_7_22_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_7_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_7_22_7  (
            .in0(_gnd_net_),
            .in1(N__31585),
            .in2(_gnd_net_),
            .in3(N__48960),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78595),
            .ce(),
            .sr(N__30495));
    defparam \c0.FRAME_MATCHER_state_i8_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_7_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_7_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__33466),
            .in2(_gnd_net_),
            .in3(N__48961),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78614),
            .ce(),
            .sr(N__33444));
    defparam \c0.FRAME_MATCHER_state_i14_LC_7_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_7_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_7_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_7_25_0  (
            .in0(_gnd_net_),
            .in1(N__29419),
            .in2(_gnd_net_),
            .in3(N__48962),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78628),
            .ce(),
            .sr(N__29400));
    defparam \quad_counter1.add_85_2_lut_LC_9_7_0 .C_ON=1'b1;
    defparam \quad_counter1.add_85_2_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_85_2_lut_LC_9_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_85_2_lut_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__29700),
            .in2(_gnd_net_),
            .in3(N__28278),
            .lcout(n39_adj_4770),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\quad_counter1.n19701 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i1_LC_9_7_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i1_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i1_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i1_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__29607),
            .in2(_gnd_net_),
            .in3(N__28275),
            .lcout(\quad_counter1.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n19701 ),
            .carryout(\quad_counter1.n19702 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i2_LC_9_7_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i2_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i2_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i2_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__29594),
            .in2(_gnd_net_),
            .in3(N__28272),
            .lcout(\quad_counter1.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n19702 ),
            .carryout(\quad_counter1.n19703 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i3_LC_9_7_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i3_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i3_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i3_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__29580),
            .in2(_gnd_net_),
            .in3(N__28269),
            .lcout(\quad_counter1.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n19703 ),
            .carryout(\quad_counter1.n19704 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i4_LC_9_7_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i4_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i4_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i4_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__29714),
            .in2(_gnd_net_),
            .in3(N__28266),
            .lcout(\quad_counter1.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n19704 ),
            .carryout(\quad_counter1.n19705 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i5_LC_9_7_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i5_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i5_LC_9_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i5_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__29739),
            .in2(_gnd_net_),
            .in3(N__28335),
            .lcout(\quad_counter1.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n19705 ),
            .carryout(\quad_counter1.n19706 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i6_LC_9_7_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i6_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i6_LC_9_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i6_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__29664),
            .in2(_gnd_net_),
            .in3(N__28332),
            .lcout(\quad_counter1.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n19706 ),
            .carryout(\quad_counter1.n19707 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i7_LC_9_7_7 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i7_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i7_LC_9_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i7_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__29550),
            .in2(_gnd_net_),
            .in3(N__28329),
            .lcout(\quad_counter1.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n19707 ),
            .carryout(\quad_counter1.n19708 ),
            .clk(N__78686),
            .ce(N__29789),
            .sr(N__29777));
    defparam \quad_counter1.a_delay_counter__i8_LC_9_8_0 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i8_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i8_LC_9_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i8_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__29619),
            .in2(_gnd_net_),
            .in3(N__28326),
            .lcout(\quad_counter1.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\quad_counter1.n19709 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i9_LC_9_8_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i9_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i9_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i9_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__29676),
            .in2(_gnd_net_),
            .in3(N__28323),
            .lcout(\quad_counter1.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n19709 ),
            .carryout(\quad_counter1.n19710 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i10_LC_9_8_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i10_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i10_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i10_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__29537),
            .in2(_gnd_net_),
            .in3(N__28320),
            .lcout(\quad_counter1.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n19710 ),
            .carryout(\quad_counter1.n19711 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i11_LC_9_8_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i11_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i11_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i11_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__29727),
            .in2(_gnd_net_),
            .in3(N__28317),
            .lcout(\quad_counter1.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n19711 ),
            .carryout(\quad_counter1.n19712 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i12_LC_9_8_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i12_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i12_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i12_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__29651),
            .in2(_gnd_net_),
            .in3(N__28314),
            .lcout(\quad_counter1.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n19712 ),
            .carryout(\quad_counter1.n19713 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i13_LC_9_8_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i13_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i13_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i13_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__29637),
            .in2(_gnd_net_),
            .in3(N__28311),
            .lcout(\quad_counter1.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n19713 ),
            .carryout(\quad_counter1.n19714 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i14_LC_9_8_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i14_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i14_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i14_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__29562),
            .in2(_gnd_net_),
            .in3(N__28428),
            .lcout(\quad_counter1.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n19714 ),
            .carryout(\quad_counter1.n19715 ),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.a_delay_counter__i15_LC_9_8_7 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i15_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i15_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i15_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__29523),
            .in2(_gnd_net_),
            .in3(N__28425),
            .lcout(\quad_counter1.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78669),
            .ce(N__29796),
            .sr(N__29778));
    defparam \quad_counter1.count_i0_i1_LC_9_9_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i1_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i1_LC_9_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i1_LC_9_9_2  (
            .in0(N__40411),
            .in1(N__32367),
            .in2(_gnd_net_),
            .in3(N__34737),
            .lcout(encoder1_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78654),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_delayed_68_LC_9_10_3 .C_ON=1'b0;
    defparam \quad_counter1.B_delayed_68_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_delayed_68_LC_9_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.B_delayed_68_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29906),
            .lcout(\quad_counter1.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78642),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i5_LC_9_11_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i5_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i5_LC_9_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i5_LC_9_11_0  (
            .in0(N__40412),
            .in1(N__32568),
            .in2(_gnd_net_),
            .in3(N__41139),
            .lcout(encoder1_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78629),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1962_2_lut_LC_9_11_4 .C_ON=1'b0;
    defparam \c0.tx.i1962_2_lut_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1962_2_lut_LC_9_11_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx.i1962_2_lut_LC_9_11_4  (
            .in0(N__28726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28774),
            .lcout(\c0.tx.n3843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_adj_1171_LC_9_11_5 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_adj_1171_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_adj_1171_LC_9_11_5 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.tx.i2_4_lut_adj_1171_LC_9_11_5  (
            .in0(N__29242),
            .in1(N__28679),
            .in2(N__28422),
            .in3(N__28373),
            .lcout(\c0.tx.n22949 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_9_12_0 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_9_12_0 .LUT_INIT=16'b1100000001001000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_9_12_0  (
            .in0(N__28341),
            .in1(N__28545),
            .in2(N__28467),
            .in3(N__28532),
            .lcout(\c0.tx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78615),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_12_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_12_1 .LUT_INIT=16'b1010101011011101;
    LogicCell40 \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_12_1  (
            .in0(N__29244),
            .in1(N__28485),
            .in2(_gnd_net_),
            .in3(N__28685),
            .lcout(),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_9_12_2 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_9_12_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_9_12_2  (
            .in0(N__28574),
            .in1(_gnd_net_),
            .in2(N__28602),
            .in3(N__38471),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78615),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_12_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_12_3 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_12_3  (
            .in0(N__28563),
            .in1(N__29970),
            .in2(N__28728),
            .in3(N__28766),
            .lcout(\c0.tx.n25080 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_adj_1172_LC_9_12_6 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_adj_1172_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_adj_1172_LC_9_12_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.tx.i1_3_lut_adj_1172_LC_9_12_6  (
            .in0(N__28439),
            .in1(N__29243),
            .in2(_gnd_net_),
            .in3(N__28530),
            .lcout(\c0.tx.n19492 ),
            .ltout(\c0.tx.n19492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_9_12_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_9_12_7 .LUT_INIT=16'b1001000011000000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_9_12_7  (
            .in0(N__28531),
            .in1(N__28727),
            .in2(N__28515),
            .in3(N__28767),
            .lcout(\c0.tx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78615),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n25080_bdd_4_lut_LC_9_13_0 .C_ON=1'b0;
    defparam \c0.tx.n25080_bdd_4_lut_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n25080_bdd_4_lut_LC_9_13_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.tx.n25080_bdd_4_lut_LC_9_13_0  (
            .in0(N__28720),
            .in1(N__28512),
            .in2(N__30039),
            .in3(N__28494),
            .lcout(),
            .ltout(\c0.tx.n25083_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1436221_i1_3_lut_LC_9_13_1 .C_ON=1'b0;
    defparam \c0.tx.i1436221_i1_3_lut_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1436221_i1_3_lut_LC_9_13_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.tx.i1436221_i1_3_lut_LC_9_13_1  (
            .in0(N__28463),
            .in1(_gnd_net_),
            .in2(N__28488),
            .in3(N__28794),
            .lcout(\c0.tx.o_Tx_Serial_N_3782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_9_13_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_9_13_2 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_9_13_2  (
            .in0(N__30202),
            .in1(N__28788),
            .in2(N__30138),
            .in3(N__28479),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_LC_9_13_3 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_LC_9_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i2_3_lut_LC_9_13_3  (
            .in0(N__28462),
            .in1(N__28722),
            .in2(_gnd_net_),
            .in3(N__28778),
            .lcout(\c0.tx.n17832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2065_LC_9_13_4.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2065_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2065_LC_9_13_4.LUT_INIT=16'b1111101101000000;
    LogicCell40 i24_3_lut_4_lut_adj_2065_LC_9_13_4 (
            .in0(N__31328),
            .in1(N__31200),
            .in2(N__30288),
            .in3(N__30351),
            .lcout(),
            .ltout(n10_adj_4776_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_9_13_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_9_13_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_9_13_5  (
            .in0(N__28803),
            .in1(N__30203),
            .in2(N__28806),
            .in3(N__30125),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n25074_bdd_4_lut_LC_9_13_6 .C_ON=1'b0;
    defparam \c0.tx.n25074_bdd_4_lut_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n25074_bdd_4_lut_LC_9_13_6 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.tx.n25074_bdd_4_lut_LC_9_13_6  (
            .in0(N__28721),
            .in1(N__28802),
            .in2(N__29871),
            .in3(N__28692),
            .lcout(\c0.tx.n25077 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_21308_LC_9_13_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_21308_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_21308_LC_9_13_7 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_21308_LC_9_13_7  (
            .in0(N__28787),
            .in1(N__29292),
            .in2(N__28779),
            .in3(N__28719),
            .lcout(\c0.tx.n25074 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_1174_LC_9_14_0 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_1174_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_1174_LC_9_14_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_1174_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__28684),
            .in2(_gnd_net_),
            .in3(N__30581),
            .lcout(\c0.tx.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__2__5483_LC_9_14_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__2__5483_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__2__5483_LC_9_14_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__2__5483_LC_9_14_1  (
            .in0(N__48379),
            .in1(N__46091),
            .in2(N__47316),
            .in3(N__29273),
            .lcout(data_out_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21192_3_lut_LC_9_14_2 .C_ON=1'b0;
    defparam \c0.i21192_3_lut_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21192_3_lut_LC_9_14_2 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i21192_3_lut_LC_9_14_2  (
            .in0(N__29139),
            .in1(N__41009),
            .in2(_gnd_net_),
            .in3(N__43061),
            .lcout(),
            .ltout(\c0.n24960_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21039_4_lut_LC_9_14_3 .C_ON=1'b0;
    defparam \c0.i21039_4_lut_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i21039_4_lut_LC_9_14_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i21039_4_lut_LC_9_14_3  (
            .in0(N__41010),
            .in1(N__32436),
            .in2(N__28617),
            .in3(N__40811),
            .lcout(),
            .ltout(\c0.n24806_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21041_4_lut_LC_9_14_4 .C_ON=1'b0;
    defparam \c0.i21041_4_lut_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21041_4_lut_LC_9_14_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.i21041_4_lut_LC_9_14_4  (
            .in0(N__31271),
            .in1(N__31415),
            .in2(N__28614),
            .in3(N__28902),
            .lcout(n24808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20990_4_lut_LC_9_14_5 .C_ON=1'b0;
    defparam \c0.i20990_4_lut_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20990_4_lut_LC_9_14_5 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \c0.i20990_4_lut_LC_9_14_5  (
            .in0(N__29307),
            .in1(N__31270),
            .in2(N__31419),
            .in3(N__34275),
            .lcout(n24757),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_9_14_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_9_14_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_9_14_7  (
            .in0(N__43060),
            .in1(_gnd_net_),
            .in2(N__37506),
            .in3(N__37698),
            .lcout(\c0.n26_adj_4645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_9_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_9_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_3_lut_3_lut_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__38174),
            .in2(_gnd_net_),
            .in3(N__38083),
            .lcout(\c0.data_out_frame_29__7__N_1143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2060_LC_9_15_2.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2060_LC_9_15_2.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2060_LC_9_15_2.LUT_INIT=16'b1010111010100010;
    LogicCell40 i24_3_lut_4_lut_adj_2060_LC_9_15_2 (
            .in0(N__28896),
            .in1(N__31176),
            .in2(N__31304),
            .in3(N__29163),
            .lcout(n10_adj_4779),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i2_LC_9_15_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i2_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i2_LC_9_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i2_LC_9_15_5  (
            .in0(N__40526),
            .in1(N__32607),
            .in2(_gnd_net_),
            .in3(N__46314),
            .lcout(encoder1_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_LC_9_15_6 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_LC_9_15_6 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \c0.tx.i1_4_lut_LC_9_15_6  (
            .in0(N__28835),
            .in1(N__29066),
            .in2(N__29088),
            .in3(N__28820),
            .lcout(),
            .ltout(\c0.tx.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i14291_4_lut_LC_9_15_7 .C_ON=1'b0;
    defparam \c0.tx.i14291_4_lut_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i14291_4_lut_LC_9_15_7 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx.i14291_4_lut_LC_9_15_7  (
            .in0(N__29051),
            .in1(N__29036),
            .in2(N__28881),
            .in3(N__29021),
            .lcout(\c0.tx.n17904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_9_16_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_9_16_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_2_lut_LC_9_16_0  (
            .in0(N__28848),
            .in1(N__38400),
            .in2(_gnd_net_),
            .in3(N__28839),
            .lcout(\c0.tx.n24889 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\c0.tx.n19723 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_9_16_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i1_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__28836),
            .in2(_gnd_net_),
            .in3(N__28824),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx.n19723 ),
            .carryout(\c0.tx.n19724 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i2_LC_9_16_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i2_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__28821),
            .in2(_gnd_net_),
            .in3(N__28809),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx.n19724 ),
            .carryout(\c0.tx.n19725 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i3_LC_9_16_3 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i3_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__29084),
            .in2(_gnd_net_),
            .in3(N__29070),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx.n19725 ),
            .carryout(\c0.tx.n19726 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i4_LC_9_16_4 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i4_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_9_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__29067),
            .in2(_gnd_net_),
            .in3(N__29055),
            .lcout(\c0.tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx.n19726 ),
            .carryout(\c0.tx.n19727 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i5_LC_9_16_5 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i5_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_9_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__29052),
            .in2(_gnd_net_),
            .in3(N__29040),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx.n19727 ),
            .carryout(\c0.tx.n19728 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i6_LC_9_16_6 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i6_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_9_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__29037),
            .in2(_gnd_net_),
            .in3(N__29025),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx.n19728 ),
            .carryout(\c0.tx.n19729 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i7_LC_9_16_7 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i7_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_9_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__29022),
            .in2(_gnd_net_),
            .in3(N__29010),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx.n19729 ),
            .carryout(\c0.tx.n19730 ),
            .clk(N__78579),
            .ce(N__38483),
            .sr(N__28964));
    defparam \c0.tx.r_Clock_Count__i8_LC_9_17_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_9_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__28987),
            .in2(_gnd_net_),
            .in3(N__29007),
            .lcout(\c0.tx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78570),
            .ce(N__38484),
            .sr(N__28965));
    defparam \c0.tx.i2_4_lut_adj_1169_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_adj_1169_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_adj_1169_LC_9_18_0 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \c0.tx.i2_4_lut_adj_1169_LC_9_18_0  (
            .in0(N__28935),
            .in1(N__29258),
            .in2(N__38478),
            .in3(N__29212),
            .lcout(),
            .ltout(\c0.tx.n14290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_9_18_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_9_18_1 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_9_18_1  (
            .in0(N__29213),
            .in1(_gnd_net_),
            .in2(N__28923),
            .in3(N__30520),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__7__5470_LC_9_18_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__7__5470_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__7__5470_LC_9_18_2 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__7__5470_LC_9_18_2  (
            .in0(N__48185),
            .in1(N__46089),
            .in2(N__44715),
            .in3(N__28916),
            .lcout(data_out_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_9_18_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_9_18_4 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_9_18_4  (
            .in0(N__31095),
            .in1(N__29291),
            .in2(N__30130),
            .in3(N__30217),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_5 .LUT_INIT=16'b1010000001000100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_5  (
            .in0(N__41038),
            .in1(N__30414),
            .in2(N__29277),
            .in3(N__43125),
            .lcout(\c0.n6_adj_4649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_9_18_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_9_18_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_9_18_6  (
            .in0(N__38467),
            .in1(N__29259),
            .in2(_gnd_net_),
            .in3(N__29214),
            .lcout(r_SM_Main_1_adj_4774),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21238_4_lut_LC_9_19_0 .C_ON=1'b0;
    defparam \c0.i21238_4_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21238_4_lut_LC_9_19_0 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i21238_4_lut_LC_9_19_0  (
            .in0(N__38274),
            .in1(N__40810),
            .in2(N__32454),
            .in3(N__41008),
            .lcout(n25006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_9_19_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_9_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_9_19_1  (
            .in0(N__29117),
            .in1(N__35085),
            .in2(_gnd_net_),
            .in3(N__43175),
            .lcout(\c0.n11_adj_4663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__1__5484_LC_9_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__1__5484_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__1__5484_LC_9_19_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_5__1__5484_LC_9_19_2  (
            .in0(N__46085),
            .in1(N__48376),
            .in2(N__47027),
            .in3(N__29135),
            .lcout(data_out_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__3__5418_LC_9_19_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__3__5418_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__3__5418_LC_9_19_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_frame_13__3__5418_LC_9_19_3  (
            .in0(N__48374),
            .in1(N__45505),
            .in2(N__29121),
            .in3(N__46088),
            .lcout(data_out_frame_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14240_4_lut_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.i14240_4_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14240_4_lut_LC_9_19_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \c0.i14240_4_lut_LC_9_19_4  (
            .in0(N__31157),
            .in1(N__29313),
            .in2(N__31303),
            .in3(N__29319),
            .lcout(\c0.n17846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__7__5454_LC_9_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__7__5454_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__7__5454_LC_9_19_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_8__7__5454_LC_9_19_5  (
            .in0(N__48375),
            .in1(N__46087),
            .in2(N__29108),
            .in3(N__39558),
            .lcout(data_out_frame_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__6__5423_LC_9_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__6__5423_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__6__5423_LC_9_19_7 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_12__6__5423_LC_9_19_7  (
            .in0(N__48373),
            .in1(N__46086),
            .in2(N__29334),
            .in3(N__33702),
            .lcout(data_out_frame_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78589),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1472_LC_9_20_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1472_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1472_LC_9_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1472_LC_9_20_2  (
            .in0(N__33471),
            .in1(N__29501),
            .in2(N__29433),
            .in3(N__49200),
            .lcout(\c0.n14_adj_4520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_20_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_20_3  (
            .in0(N__30018),
            .in1(N__43034),
            .in2(_gnd_net_),
            .in3(N__29330),
            .lcout(\c0.n11_adj_4703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21265_2_lut_3_lut_LC_9_20_4 .C_ON=1'b0;
    defparam \c0.i21265_2_lut_3_lut_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21265_2_lut_3_lut_LC_9_20_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.i21265_2_lut_3_lut_LC_9_20_4  (
            .in0(N__30565),
            .in1(N__30526),
            .in2(_gnd_net_),
            .in3(N__39441),
            .lcout(\c0.tx_transmit_N_3650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_9_20_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_9_20_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \c0.i1_3_lut_LC_9_20_5  (
            .in0(N__40648),
            .in1(N__43032),
            .in2(_gnd_net_),
            .in3(N__40929),
            .lcout(\c0.n5_adj_4334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1345_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1345_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1345_LC_9_20_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1345_LC_9_20_6  (
            .in0(N__30072),
            .in1(N__29357),
            .in2(_gnd_net_),
            .in3(N__29375),
            .lcout(\c0.n4_adj_4332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_9_20_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_9_20_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_9_20_7  (
            .in0(N__41805),
            .in1(N__43033),
            .in2(_gnd_net_),
            .in3(N__31004),
            .lcout(\c0.n26_adj_4662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1413__i0_LC_9_21_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i0_LC_9_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i0_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i0_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__43054),
            .in2(N__33215),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\c0.n19795 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i1_LC_9_21_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i1_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i1_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i1_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__40684),
            .in2(_gnd_net_),
            .in3(N__29295),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n19795 ),
            .carryout(\c0.n19796 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i2_LC_9_21_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i2_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i2_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i2_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__40995),
            .in2(_gnd_net_),
            .in3(N__29388),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(\c0.n19796 ),
            .carryout(\c0.n19797 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i3_LC_9_21_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i3_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i3_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i3_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__31156),
            .in2(_gnd_net_),
            .in3(N__29385),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(\c0.n19797 ),
            .carryout(\c0.n19798 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i4_LC_9_21_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i4_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i4_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i4_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__31266),
            .in2(_gnd_net_),
            .in3(N__29382),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(\c0.n19798 ),
            .carryout(\c0.n19799 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i5_LC_9_21_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i5_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i5_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i5_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__30090),
            .in2(_gnd_net_),
            .in3(N__29379),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(\c0.n19799 ),
            .carryout(\c0.n19800 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i6_LC_9_21_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1413__i6_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i6_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i6_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__29376),
            .in2(_gnd_net_),
            .in3(N__29364),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(\c0.n19800 ),
            .carryout(\c0.n19801 ),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.byte_transmit_counter_1413__i7_LC_9_21_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1413__i7_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1413__i7_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1413__i7_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__29358),
            .in2(_gnd_net_),
            .in3(N__29361),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78605),
            .ce(N__30471),
            .sr(N__30462));
    defparam \c0.FRAME_MATCHER_state_i17_LC_9_22_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_9_22_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_9_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__31559),
            .in2(_gnd_net_),
            .in3(N__48837),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78616),
            .ce(),
            .sr(N__29457));
    defparam \c0.i1_2_lut_4_lut_adj_1812_LC_9_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1812_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1812_LC_9_23_0 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1812_LC_9_23_0  (
            .in0(N__35784),
            .in1(N__44219),
            .in2(N__35463),
            .in3(N__38951),
            .lcout(\c0.n21611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i3_LC_9_23_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_9_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_9_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__35453),
            .in2(_gnd_net_),
            .in3(N__48825),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78630),
            .ce(),
            .sr(N__29346));
    defparam \c0.i1_2_lut_4_lut_adj_1845_LC_9_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1845_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1845_LC_9_23_2 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1845_LC_9_23_2  (
            .in0(N__35785),
            .in1(N__44220),
            .in2(N__33525),
            .in3(N__38952),
            .lcout(\c0.n21575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1846_LC_9_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1846_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1846_LC_9_23_4 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1846_LC_9_23_4  (
            .in0(N__35786),
            .in1(N__44221),
            .in2(N__29505),
            .in3(N__38953),
            .lcout(\c0.n21573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1909_LC_9_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1909_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1909_LC_9_23_7 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1909_LC_9_23_7  (
            .in0(N__38954),
            .in1(N__31558),
            .in2(N__44226),
            .in3(N__35787),
            .lcout(\c0.n21581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i9_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_9_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_9_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__33523),
            .in2(_gnd_net_),
            .in3(N__48838),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78643),
            .ce(),
            .sr(N__29445));
    defparam \c0.i1_2_lut_4_lut_adj_1858_LC_9_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1858_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1858_LC_9_25_3 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1858_LC_9_25_3  (
            .in0(N__35757),
            .in1(N__44225),
            .in2(N__29429),
            .in3(N__38955),
            .lcout(\c0.n21577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14287_2_lut_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.rx.i14287_2_lut_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14287_2_lut_LC_9_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i14287_2_lut_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__31899),
            .in2(_gnd_net_),
            .in3(N__31658),
            .lcout(\c0.rx.r_SM_Main_2_N_3680_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__36249),
            .in2(_gnd_net_),
            .in3(N__48991),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78685),
            .ce(),
            .sr(N__36225));
    defparam \quad_counter1.quadA_delayed_61_LC_10_6_0 .C_ON=1'b0;
    defparam \quad_counter1.quadA_delayed_61_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadA_delayed_61_LC_10_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.quadA_delayed_61_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29853),
            .lcout(quadA_delayed_adj_4767),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78701),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_10_6_1 .C_ON=1'b0;
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_10_6_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.quadA_I_0_73_2_lut_LC_10_6_1  (
            .in0(N__29852),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29815),
            .lcout(a_delay_counter_15__N_4123_adj_4772),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_LC_10_7_0 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_LC_10_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_LC_10_7_0  (
            .in0(N__29625),
            .in1(N__29511),
            .in2(N__29685),
            .in3(N__29568),
            .lcout(n9806),
            .ltout(n9806_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_63_LC_10_7_1 .C_ON=1'b0;
    defparam \quad_counter1.A_63_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_63_LC_10_7_1 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \quad_counter1.A_63_LC_10_7_1  (
            .in0(N__29846),
            .in1(N__29817),
            .in2(N__29856),
            .in3(N__30656),
            .lcout(A_filtered_adj_4763),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78688),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_10_7_3.C_ON=1'b0;
    defparam i1_3_lut_LC_10_7_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_10_7_3.LUT_INIT=16'b1111111101100110;
    LogicCell40 i1_3_lut_LC_10_7_3 (
            .in0(N__29845),
            .in1(N__29816),
            .in2(_gnd_net_),
            .in3(N__29802),
            .lcout(n14345),
            .ltout(n14345_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i0_LC_10_7_4 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i0_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i0_LC_10_7_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \quad_counter1.a_delay_counter__i0_LC_10_7_4  (
            .in0(N__29770),
            .in1(N__29699),
            .in2(N__29748),
            .in3(N__29745),
            .lcout(a_delay_counter_0_adj_4765),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78688),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_LC_10_7_6 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_LC_10_7_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter1.i9_4_lut_LC_10_7_6  (
            .in0(N__29738),
            .in1(N__29726),
            .in2(N__29715),
            .in3(N__29698),
            .lcout(\quad_counter1.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_LC_10_7_7 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_LC_10_7_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_LC_10_7_7  (
            .in0(N__29675),
            .in1(N__29663),
            .in2(N__29652),
            .in3(N__29636),
            .lcout(\quad_counter1.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_LC_10_8_5 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_LC_10_8_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter1.i12_4_lut_LC_10_8_5  (
            .in0(N__29618),
            .in1(N__29606),
            .in2(N__29595),
            .in3(N__29579),
            .lcout(\quad_counter1.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_LC_10_8_6 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_LC_10_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_LC_10_8_6  (
            .in0(N__29561),
            .in1(N__29549),
            .in2(N__29538),
            .in3(N__29522),
            .lcout(\quad_counter1.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_10_9_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_10_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_10_9_0  (
            .in0(N__31662),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31917),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78656),
            .ce(),
            .sr(N__49881));
    defparam CONSTANT_ONE_LUT4_LC_10_9_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_9_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_9_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_LC_10_10_1 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_LC_10_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter1.i3_4_lut_LC_10_10_1  (
            .in0(N__29877),
            .in1(N__30623),
            .in2(N__29907),
            .in3(N__30658),
            .lcout(count_enable_adj_4769),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_delayed_67_LC_10_10_3 .C_ON=1'b0;
    defparam \quad_counter1.A_delayed_67_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_delayed_67_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.A_delayed_67_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30659),
            .lcout(\quad_counter1.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78644),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1075_1_lut_2_lut_LC_10_10_5 .C_ON=1'b0;
    defparam \quad_counter1.i1075_1_lut_2_lut_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1075_1_lut_2_lut_LC_10_10_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter1.i1075_1_lut_2_lut_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__30622),
            .in2(_gnd_net_),
            .in3(N__30657),
            .lcout(\quad_counter1.n2226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_10_11_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_10_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_10_11_7  (
            .in0(N__30732),
            .in1(N__45540),
            .in2(_gnd_net_),
            .in3(N__43222),
            .lcout(\c0.n5_adj_4660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2017_LC_10_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2017_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2017_LC_10_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_2017_LC_10_12_0  (
            .in0(N__35112),
            .in1(N__32140),
            .in2(N__41779),
            .in3(N__34154),
            .lcout(\c0.data_out_frame_29__7__N_1148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_10_12_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_10_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_10_12_2  (
            .in0(N__33693),
            .in1(N__32201),
            .in2(N__33995),
            .in3(N__33855),
            .lcout(\c0.n12464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_10_12_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_10_12_3 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_10_12_3  (
            .in0(N__29870),
            .in1(N__29925),
            .in2(N__30147),
            .in3(N__30201),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1699_LC_10_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1699_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1699_LC_10_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1699_LC_10_12_4  (
            .in0(N__32706),
            .in1(N__33854),
            .in2(N__33700),
            .in3(N__32141),
            .lcout(\c0.n22291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_10_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_10_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_10_12_5  (
            .in0(N__38165),
            .in1(N__34609),
            .in2(_gnd_net_),
            .in3(N__38031),
            .lcout(\c0.n6_adj_4456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1680_LC_10_12_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1680_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1680_LC_10_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1680_LC_10_12_6  (
            .in0(N__32707),
            .in1(N__32200),
            .in2(N__33994),
            .in3(N__32142),
            .lcout(\c0.n21391 ),
            .ltout(\c0.n21391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1529_LC_10_12_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1529_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1529_LC_10_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1529_LC_10_12_7  (
            .in0(N__38164),
            .in1(N__38226),
            .in2(N__29916),
            .in3(N__38059),
            .lcout(\c0.n12539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1885_LC_10_13_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1885_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1885_LC_10_13_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i12_4_lut_adj_1885_LC_10_13_0  (
            .in0(N__34433),
            .in1(N__37287),
            .in2(N__35297),
            .in3(N__30941),
            .lcout(\c0.n28_adj_4698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i21252_3_lut_LC_10_13_2.C_ON=1'b0;
    defparam i21252_3_lut_LC_10_13_2.SEQ_MODE=4'b0000;
    defparam i21252_3_lut_LC_10_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 i21252_3_lut_LC_10_13_2 (
            .in0(N__32928),
            .in1(N__31199),
            .in2(_gnd_net_),
            .in3(N__32088),
            .lcout(n25021),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1205_LC_10_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1205_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1205_LC_10_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1205_LC_10_13_3  (
            .in0(N__38177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38228),
            .lcout(\c0.n21362 ),
            .ltout(\c0.n21362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1967_LC_10_13_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1967_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1967_LC_10_13_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1967_LC_10_13_4  (
            .in0(N__34765),
            .in1(N__41364),
            .in2(N__29913),
            .in3(N__37265),
            .lcout(\c0.n21244 ),
            .ltout(\c0.n21244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_2006_LC_10_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_2006_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_2006_LC_10_13_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_2006_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__37115),
            .in2(N__29910),
            .in3(N__41413),
            .lcout(\c0.n21309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i25_LC_10_13_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i25_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i25_LC_10_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i25_LC_10_13_6  (
            .in0(N__40467),
            .in1(N__32769),
            .in2(_gnd_net_),
            .in3(N__35344),
            .lcout(encoder1_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78607),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1841_LC_10_13_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1841_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1841_LC_10_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1841_LC_10_13_7  (
            .in0(N__38176),
            .in1(N__38227),
            .in2(_gnd_net_),
            .in3(N__46590),
            .lcout(\c0.n21475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__4__5297_LC_10_14_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__4__5297_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__4__5297_LC_10_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__4__5297_LC_10_14_0  (
            .in0(N__38090),
            .in1(N__32232),
            .in2(N__30810),
            .in3(N__46606),
            .lcout(\c0.data_out_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78598),
            .ce(N__45036),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1308_LC_10_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1308_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1308_LC_10_14_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1308_LC_10_14_1  (
            .in0(N__36707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37939),
            .lcout(\c0.n22163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1272_LC_10_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1272_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1272_LC_10_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1272_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__35040),
            .in2(_gnd_net_),
            .in3(N__32345),
            .lcout(),
            .ltout(\c0.n6_adj_4297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1274_LC_10_14_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1274_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1274_LC_10_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1274_LC_10_14_3  (
            .in0(N__29952),
            .in1(N__42147),
            .in2(N__29946),
            .in3(N__34155),
            .lcout(\c0.n12604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_10_14_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_10_14_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_10_14_4  (
            .in0(N__29943),
            .in1(N__45075),
            .in2(_gnd_net_),
            .in3(N__43220),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i21253_4_lut_LC_10_14_5.C_ON=1'b0;
    defparam i21253_4_lut_LC_10_14_5.SEQ_MODE=4'b0000;
    defparam i21253_4_lut_LC_10_14_5.LUT_INIT=16'b0111010100100000;
    LogicCell40 i21253_4_lut_LC_10_14_5 (
            .in0(N__31319),
            .in1(N__31418),
            .in2(N__29937),
            .in3(N__29934),
            .lcout(n25022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1765_LC_10_14_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1765_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1765_LC_10_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1765_LC_10_14_6  (
            .in0(N__37938),
            .in1(N__34650),
            .in2(_gnd_net_),
            .in3(N__36706),
            .lcout(\c0.n22593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1177_LC_10_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1177_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1177_LC_10_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1177_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__41430),
            .in2(_gnd_net_),
            .in3(N__38089),
            .lcout(\c0.n22757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1683_LC_10_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1683_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1683_LC_10_15_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1683_LC_10_15_1  (
            .in0(N__38254),
            .in1(N__46221),
            .in2(N__38189),
            .in3(N__32261),
            .lcout(\c0.n22544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1684_LC_10_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1684_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1684_LC_10_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1684_LC_10_15_2  (
            .in0(N__30844),
            .in1(N__38178),
            .in2(N__38265),
            .in3(N__46213),
            .lcout(\c0.n22478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1835_LC_10_15_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1835_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1835_LC_10_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1835_LC_10_15_3  (
            .in0(N__38179),
            .in1(N__50574),
            .in2(N__38263),
            .in3(N__41495),
            .lcout(\c0.n24033 ),
            .ltout(\c0.n24033_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1476_LC_10_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1476_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1476_LC_10_15_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1476_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__38180),
            .in2(N__29985),
            .in3(N__38025),
            .lcout(n21307),
            .ltout(n21307_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_10_15_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_10_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_LC_10_15_5  (
            .in0(N__32260),
            .in1(N__37721),
            .in2(N__29982),
            .in3(N__50651),
            .lcout(),
            .ltout(\c0.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1184_LC_10_15_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1184_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1184_LC_10_15_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1184_LC_10_15_6  (
            .in0(N__32233),
            .in1(N__30825),
            .in2(N__29979),
            .in3(N__29976),
            .lcout(\c0.n22475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1992_LC_10_15_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1992_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1992_LC_10_15_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1992_LC_10_15_7  (
            .in0(N__32259),
            .in1(N__46132),
            .in2(N__37138),
            .in3(N__30772),
            .lcout(\c0.n23918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_10_16_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_10_16_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i13_LC_10_16_0  (
            .in0(N__50436),
            .in1(N__37812),
            .in2(_gnd_net_),
            .in3(N__37872),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78582),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i22_LC_10_16_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i22_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i22_LC_10_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i22_LC_10_16_1  (
            .in0(N__40485),
            .in1(N__32790),
            .in2(_gnd_net_),
            .in3(N__34649),
            .lcout(encoder1_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78582),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__2__5475_LC_10_16_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__2__5475_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__2__5475_LC_10_16_4 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_frame_6__2__5475_LC_10_16_4  (
            .in0(N__30902),
            .in1(N__46083),
            .in2(N__37056),
            .in3(N__48362),
            .lcout(data_out_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78582),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_10_16_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_10_16_5 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_10_16_5  (
            .in0(N__29966),
            .in1(N__30139),
            .in2(N__30221),
            .in3(N__31038),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78582),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1734_LC_10_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1734_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1734_LC_10_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1734_LC_10_16_6  (
            .in0(N__38184),
            .in1(N__38010),
            .in2(N__40032),
            .in3(N__37209),
            .lcout(\c0.n20341 ),
            .ltout(\c0.n20341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2031_LC_10_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2031_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2031_LC_10_16_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2031_LC_10_16_7  (
            .in0(N__38011),
            .in1(N__38262),
            .in2(N__30261),
            .in3(N__46607),
            .lcout(\c0.n12514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__5__5432_LC_10_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__5__5432_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__5__5432_LC_10_17_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_11__5__5432_LC_10_17_1  (
            .in0(N__48348),
            .in1(N__46062),
            .in2(N__40278),
            .in3(N__30308),
            .lcout(data_out_frame_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__7__5414_LC_10_17_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__7__5414_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__7__5414_LC_10_17_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_13__7__5414_LC_10_17_2  (
            .in0(N__46060),
            .in1(N__34595),
            .in2(N__48378),
            .in3(N__30254),
            .lcout(data_out_frame_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__7__5438_LC_10_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__7__5438_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__7__5438_LC_10_17_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__7__5438_LC_10_17_3  (
            .in0(N__48347),
            .in1(N__46061),
            .in2(N__40335),
            .in3(N__30236),
            .lcout(data_out_frame_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_10_17_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_10_17_4 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_10_17_4  (
            .in0(N__30318),
            .in1(N__30032),
            .in2(N__30222),
            .in3(N__30129),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__1__5420_LC_10_17_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__1__5420_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__1__5420_LC_10_17_5 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_13__1__5420_LC_10_17_5  (
            .in0(N__48349),
            .in1(N__32468),
            .in2(N__34785),
            .in3(N__46063),
            .lcout(data_out_frame_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__6__5415_LC_10_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__6__5415_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__6__5415_LC_10_17_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_13__6__5415_LC_10_17_6  (
            .in0(N__46059),
            .in1(N__34437),
            .in2(N__48377),
            .in3(N__30017),
            .lcout(data_out_frame_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__3__5458_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__3__5458_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__3__5458_LC_10_18_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__3__5458_LC_10_18_0  (
            .in0(N__48345),
            .in1(N__46022),
            .in2(N__36564),
            .in3(N__29999),
            .lcout(data_out_frame_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21029_4_lut_LC_10_18_1 .C_ON=1'b0;
    defparam \c0.i21029_4_lut_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21029_4_lut_LC_10_18_1 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.i21029_4_lut_LC_10_18_1  (
            .in0(N__31313),
            .in1(N__30786),
            .in2(N__31416),
            .in3(N__31473),
            .lcout(n24796),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__7__5462_LC_10_18_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__7__5462_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__7__5462_LC_10_18_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_7__7__5462_LC_10_18_3  (
            .in0(N__46021),
            .in1(N__48346),
            .in2(N__42720),
            .in3(N__30335),
            .lcout(data_out_frame_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_10_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_10_18_5 .LUT_INIT=16'b1111010101000100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_10_18_5  (
            .in0(N__40996),
            .in1(N__30372),
            .in2(N__34860),
            .in3(N__43164),
            .lcout(\c0.n6_adj_4659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21038_4_lut_LC_10_18_6 .C_ON=1'b0;
    defparam \c0.i21038_4_lut_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i21038_4_lut_LC_10_18_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.i21038_4_lut_LC_10_18_6  (
            .in0(N__31071),
            .in1(N__34512),
            .in2(N__31318),
            .in3(N__31401),
            .lcout(),
            .ltout(n24805_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_LC_10_18_7.C_ON=1'b0;
    defparam i24_3_lut_4_lut_LC_10_18_7.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_LC_10_18_7.LUT_INIT=16'b1111010010110000;
    LogicCell40 i24_3_lut_4_lut_LC_10_18_7 (
            .in0(N__31314),
            .in1(N__31158),
            .in2(N__30321),
            .in3(N__30426),
            .lcout(n10_adj_4780),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21323_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21323_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21323_LC_10_19_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_21323_LC_10_19_0  (
            .in0(N__38648),
            .in1(N__40806),
            .in2(N__30312),
            .in3(N__43179),
            .lcout(),
            .ltout(\c0.n25092_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25092_bdd_4_lut_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.n25092_bdd_4_lut_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.n25092_bdd_4_lut_LC_10_19_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n25092_bdd_4_lut_LC_10_19_1  (
            .in0(N__40807),
            .in1(N__35403),
            .in2(N__30294),
            .in3(N__30269),
            .lcout(),
            .ltout(\c0.n25095_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21246_4_lut_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.i21246_4_lut_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21246_4_lut_LC_10_19_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.i21246_4_lut_LC_10_19_2  (
            .in0(N__41000),
            .in1(N__30420),
            .in2(N__30291),
            .in3(N__40809),
            .lcout(n25014),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__5__5448_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__5__5448_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__5__5448_LC_10_19_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_9__5__5448_LC_10_19_4  (
            .in0(N__48372),
            .in1(N__46026),
            .in2(N__30273),
            .in3(N__45399),
            .lcout(data_out_frame_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78590),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21240_4_lut_LC_10_19_5 .C_ON=1'b0;
    defparam \c0.i21240_4_lut_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21240_4_lut_LC_10_19_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.i21240_4_lut_LC_10_19_5  (
            .in0(N__40808),
            .in1(N__30978),
            .in2(N__30927),
            .in3(N__41001),
            .lcout(n25008),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_10_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_10_19_7  (
            .in0(N__43178),
            .in1(N__35148),
            .in2(_gnd_net_),
            .in3(N__30387),
            .lcout(\c0.n11_adj_4681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21185_4_lut_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.i21185_4_lut_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21185_4_lut_LC_10_20_0 .LUT_INIT=16'b1000110100000000;
    LogicCell40 \c0.i21185_4_lut_LC_10_20_0  (
            .in0(N__40949),
            .in1(N__30404),
            .in2(N__40685),
            .in3(N__43053),
            .lcout(\c0.n24953 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21222_2_lut_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.i21222_2_lut_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21222_2_lut_LC_10_20_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i21222_2_lut_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__40650),
            .in2(_gnd_net_),
            .in3(N__30395),
            .lcout(\c0.n24897 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__0__5485_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__0__5485_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__0__5485_LC_10_20_2 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__0__5485_LC_10_20_2  (
            .in0(N__48294),
            .in1(N__46025),
            .in2(N__45189),
            .in3(N__30405),
            .lcout(data_out_frame_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78599),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__2__5523_LC_10_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__2__5523_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__2__5523_LC_10_20_3 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \c0.data_out_frame_0__2__5523_LC_10_20_3  (
            .in0(N__33380),
            .in1(N__30396),
            .in2(N__43838),
            .in3(N__43925),
            .lcout(data_out_frame_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78599),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__5__5424_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__5__5424_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__5__5424_LC_10_20_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_12__5__5424_LC_10_20_4  (
            .in0(N__48293),
            .in1(N__46024),
            .in2(N__32715),
            .in3(N__30386),
            .lcout(data_out_frame_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78599),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21161_2_lut_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.i21161_2_lut_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21161_2_lut_LC_10_20_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.i21161_2_lut_LC_10_20_5  (
            .in0(N__30359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40649),
            .lcout(\c0.n24900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1579_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1579_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1579_LC_10_20_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i2_3_lut_adj_1579_LC_10_20_6  (
            .in0(N__30437),
            .in1(N__30456),
            .in2(_gnd_net_),
            .in3(N__39038),
            .lcout(n14247),
            .ltout(n14247_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__3__5522_LC_10_20_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__3__5522_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__3__5522_LC_10_20_7 .LUT_INIT=16'b0011101011111010;
    LogicCell40 \c0.data_out_frame_0__3__5522_LC_10_20_7  (
            .in0(N__30360),
            .in1(N__43829),
            .in2(N__30363),
            .in3(N__43926),
            .lcout(data_out_frame_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78599),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1946_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1946_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1946_LC_10_21_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \c0.i3_4_lut_adj_1946_LC_10_21_1  (
            .in0(N__33600),
            .in1(N__35963),
            .in2(N__31614),
            .in3(N__39111),
            .lcout(),
            .ltout(\c0.n8_adj_4740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19189_4_lut_LC_10_21_2 .C_ON=1'b0;
    defparam \c0.i19189_4_lut_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i19189_4_lut_LC_10_21_2 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \c0.i19189_4_lut_LC_10_21_2  (
            .in0(N__39112),
            .in1(N__35826),
            .in2(N__30477),
            .in3(N__35470),
            .lcout(\c0.n22952 ),
            .ltout(\c0.n22952_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1960_LC_10_21_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1960_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1960_LC_10_21_3 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \c0.i2_3_lut_adj_1960_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__30447),
            .in2(N__30474),
            .in3(N__43533),
            .lcout(\c0.n14380 ),
            .ltout(\c0.n14380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11327_2_lut_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.i11327_2_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11327_2_lut_LC_10_21_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.i11327_2_lut_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30465),
            .in3(N__44004),
            .lcout(\c0.n14942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2553_3_lut_4_lut_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.i2553_3_lut_4_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2553_3_lut_4_lut_LC_10_21_5 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \c0.i2553_3_lut_4_lut_LC_10_21_5  (
            .in0(N__39488),
            .in1(N__43830),
            .in2(N__48323),
            .in3(N__43923),
            .lcout(\c0.n4728 ),
            .ltout(\c0.n4728_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i75_3_lut_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.i75_3_lut_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i75_3_lut_LC_10_21_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.i75_3_lut_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__35719),
            .in2(N__30450),
            .in3(N__44003),
            .lcout(\c0.n58_adj_4742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_5282_LC_10_21_7 .C_ON=1'b0;
    defparam \c0.tx_transmit_5282_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_5282_LC_10_21_7 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \c0.tx_transmit_5282_LC_10_21_7  (
            .in0(N__35720),
            .in1(N__33198),
            .in2(N__48324),
            .in3(N__39039),
            .lcout(\c0.r_SM_Main_2_N_3754_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78608),
            .ce(),
            .sr(N__30441));
    defparam \c0.rx.i2_4_lut_adj_1167_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_adj_1167_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_adj_1167_LC_10_22_3 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \c0.rx.i2_4_lut_adj_1167_LC_10_22_3  (
            .in0(N__50025),
            .in1(N__42007),
            .in2(N__50157),
            .in3(N__49944),
            .lcout(n14484),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_10_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_10_22_5 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_10_22_5  (
            .in0(N__30555),
            .in1(N__30528),
            .in2(N__39458),
            .in3(N__39144),
            .lcout(\c0.n9_adj_4549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__4__5441_LC_10_22_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__4__5441_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__4__5441_LC_10_22_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__4__5441_LC_10_22_6  (
            .in0(N__48271),
            .in1(N__46030),
            .in2(N__39990),
            .in3(N__33254),
            .lcout(data_out_frame_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78619),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13932_2_lut_LC_10_22_7 .C_ON=1'b0;
    defparam \c0.i13932_2_lut_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13932_2_lut_LC_10_22_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i13932_2_lut_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__30554),
            .in2(_gnd_net_),
            .in3(N__30527),
            .lcout(\c0.n17533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1197_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1197_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1197_LC_10_23_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \c0.i1_4_lut_adj_1197_LC_10_23_0  (
            .in0(N__39114),
            .in1(N__48511),
            .in2(N__35691),
            .in3(N__30483),
            .lcout(\c0.n5 ),
            .ltout(\c0.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i22_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_10_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_10_23_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30498),
            .in3(N__35901),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78632),
            .ce(),
            .sr(N__31605));
    defparam \c0.i1_2_lut_4_lut_adj_1942_LC_10_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1942_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1942_LC_10_23_2 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1942_LC_10_23_2  (
            .in0(N__35780),
            .in1(N__44197),
            .in2(N__36171),
            .in3(N__38944),
            .lcout(\c0.n21595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1943_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1943_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1943_LC_10_23_3 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1943_LC_10_23_3  (
            .in0(N__38945),
            .in1(N__31593),
            .in2(N__44217),
            .in3(N__35781),
            .lcout(\c0.n21585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1947_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1947_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1947_LC_10_23_4 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1947_LC_10_23_4  (
            .in0(N__35782),
            .in1(N__44201),
            .in2(N__33610),
            .in3(N__38946),
            .lcout(\c0.n21587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1958_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1958_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1958_LC_10_23_5 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1958_LC_10_23_5  (
            .in0(N__38947),
            .in1(N__31692),
            .in2(N__44218),
            .in3(N__35783),
            .lcout(\c0.n21597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_2037_LC_10_23_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_2037_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_2037_LC_10_23_7 .LUT_INIT=16'b0011000100000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_2037_LC_10_23_7  (
            .in0(N__39451),
            .in1(N__39143),
            .in2(N__39392),
            .in3(N__39113),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i30_LC_10_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_10_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_10_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__31691),
            .in2(_gnd_net_),
            .in3(N__48824),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78645),
            .ce(),
            .sr(N__30600));
    defparam \c0.FRAME_MATCHER_state_i16_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_10_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_10_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__35545),
            .in2(_gnd_net_),
            .in3(N__48870),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78655),
            .ce(),
            .sr(N__33633));
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_10_26_0  (
            .in0(_gnd_net_),
            .in1(N__33592),
            .in2(_gnd_net_),
            .in3(N__48882),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78671),
            .ce(),
            .sr(N__30594));
    defparam \c0.FRAME_MATCHER_state_i23_LC_11_7_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_11_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_11_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__49103),
            .in2(_gnd_net_),
            .in3(N__48984),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78703),
            .ce(),
            .sr(N__31845));
    defparam \c0.i6_4_lut_adj_1385_LC_11_8_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1385_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1385_LC_11_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1385_LC_11_8_3  (
            .in0(N__32099),
            .in1(N__30681),
            .in2(N__45613),
            .in3(N__39797),
            .lcout(\c0.n14_adj_4368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i4_LC_11_8_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i4_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i4_LC_11_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i4_LC_11_8_4  (
            .in0(N__47648),
            .in1(N__36282),
            .in2(_gnd_net_),
            .in3(N__45228),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78690),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1600_LC_11_8_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1600_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1600_LC_11_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1600_LC_11_8_5  (
            .in0(N__46357),
            .in1(N__45506),
            .in2(N__34780),
            .in3(N__34610),
            .lcout(\c0.n22218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i1_LC_11_8_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i1_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i1_LC_11_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i1_LC_11_8_6  (
            .in0(N__47647),
            .in1(N__36315),
            .in2(_gnd_net_),
            .in3(N__36349),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78690),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1282_LC_11_9_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1282_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1282_LC_11_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1282_LC_11_9_0  (
            .in0(N__34091),
            .in1(N__38809),
            .in2(N__33911),
            .in3(N__33884),
            .lcout(),
            .ltout(\c0.n10_adj_4303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_2002_LC_11_9_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_2002_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_2002_LC_11_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_2002_LC_11_9_1  (
            .in0(N__45612),
            .in1(N__39549),
            .in2(N__30585),
            .in3(N__39626),
            .lcout(\c0.n21399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1367_LC_11_9_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1367_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1367_LC_11_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1367_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__36788),
            .in2(_gnd_net_),
            .in3(N__36870),
            .lcout(\c0.n22531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i29_LC_11_9_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i29_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i29_LC_11_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i29_LC_11_9_5  (
            .in0(N__36843),
            .in1(N__47598),
            .in2(_gnd_net_),
            .in3(N__36871),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78673),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i13_LC_11_9_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i13_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i13_LC_11_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i13_LC_11_9_7  (
            .in0(N__40440),
            .in1(N__32661),
            .in2(_gnd_net_),
            .in3(N__32694),
            .lcout(encoder1_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78673),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i14_LC_11_10_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i14_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i14_LC_11_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i14_LC_11_10_0  (
            .in0(N__40409),
            .in1(N__32643),
            .in2(_gnd_net_),
            .in3(N__33671),
            .lcout(encoder1_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1355_LC_11_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1355_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1355_LC_11_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1355_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__36801),
            .in2(_gnd_net_),
            .in3(N__30680),
            .lcout(\c0.n22800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1281_LC_11_10_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1281_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1281_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1281_LC_11_10_4  (
            .in0(N__36489),
            .in1(N__30609),
            .in2(_gnd_net_),
            .in3(N__44409),
            .lcout(\c0.n22611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1352_LC_11_10_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1352_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1352_LC_11_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1352_LC_11_10_5  (
            .in0(N__36951),
            .in1(N__39625),
            .in2(_gnd_net_),
            .in3(N__44707),
            .lcout(\c0.n13741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1307_LC_11_10_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1307_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1307_LC_11_10_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1307_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__32684),
            .in2(_gnd_net_),
            .in3(N__32139),
            .lcout(\c0.n22294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1349_LC_11_10_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1349_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1349_LC_11_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1349_LC_11_10_7  (
            .in0(N__30608),
            .in1(N__30743),
            .in2(N__38685),
            .in3(N__36490),
            .lcout(\c0.n13121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.encoder0_position_27__I_0_2_lut_LC_11_11_0 .C_ON=1'b0;
    defparam \c0.encoder0_position_27__I_0_2_lut_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.encoder0_position_27__I_0_2_lut_LC_11_11_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.encoder0_position_27__I_0_2_lut_LC_11_11_0  (
            .in0(N__37034),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45598),
            .lcout(\c0.data_out_frame_29__7__N_849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i11_LC_11_11_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i11_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i11_LC_11_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i11_LC_11_11_2  (
            .in0(N__40410),
            .in1(N__32745),
            .in2(_gnd_net_),
            .in3(N__35116),
            .lcout(encoder1_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_2005_LC_11_11_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_2005_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_2005_LC_11_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_2005_LC_11_11_3  (
            .in0(N__36540),
            .in1(N__37033),
            .in2(N__42611),
            .in3(N__41326),
            .lcout(\c0.n22246 ),
            .ltout(\c0.n22246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1368_LC_11_11_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1368_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1368_LC_11_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1368_LC_11_11_4  (
            .in0(N__36488),
            .in1(N__42658),
            .in2(N__30684),
            .in3(N__36597),
            .lcout(\c0.n22846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i9_LC_11_11_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i9_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i9_LC_11_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i9_LC_11_11_5  (
            .in0(N__40413),
            .in1(N__32523),
            .in2(_gnd_net_),
            .in3(N__40064),
            .lcout(encoder1_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78646),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i10_LC_11_11_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i10_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i10_LC_11_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i10_LC_11_11_7  (
            .in0(N__36598),
            .in1(N__47597),
            .in2(_gnd_net_),
            .in3(N__36579),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1306_LC_11_12_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1306_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1306_LC_11_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1306_LC_11_12_0  (
            .in0(N__43292),
            .in1(N__30717),
            .in2(_gnd_net_),
            .in3(N__43416),
            .lcout(\c0.n20379 ),
            .ltout(\c0.n20379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1578_LC_11_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1578_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1578_LC_11_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1578_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__41753),
            .in2(N__30666),
            .in3(N__32138),
            .lcout(\c0.n13938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_11_12_3 .C_ON=1'b0;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_11_12_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.A_filtered_I_0_2_lut_LC_11_12_3  (
            .in0(N__30663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30630),
            .lcout(\quad_counter1.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1235_LC_11_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1235_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1235_LC_11_12_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1235_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__37116),
            .in2(_gnd_net_),
            .in3(N__41412),
            .lcout(n21484),
            .ltout(n21484_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1816_LC_11_12_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1816_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1816_LC_11_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1816_LC_11_12_6  (
            .in0(N__41232),
            .in1(N__30753),
            .in2(N__30747),
            .in3(N__41491),
            .lcout(\c0.n22452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1252_LC_11_12_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1252_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1252_LC_11_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1252_LC_11_12_7  (
            .in0(N__39982),
            .in1(N__34320),
            .in2(_gnd_net_),
            .in3(N__30744),
            .lcout(\c0.n13384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__0__5469_LC_11_13_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__0__5469_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__0__5469_LC_11_13_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_7__0__5469_LC_11_13_0  (
            .in0(N__48189),
            .in1(N__46095),
            .in2(N__32502),
            .in3(N__36802),
            .lcout(data_out_frame_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__3__5466_LC_11_13_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__3__5466_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__3__5466_LC_11_13_2 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_7__3__5466_LC_11_13_2  (
            .in0(N__48190),
            .in1(N__46096),
            .in2(N__42408),
            .in3(N__30731),
            .lcout(data_out_frame_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1305_LC_11_13_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1305_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1305_LC_11_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1305_LC_11_13_4  (
            .in0(N__42818),
            .in1(N__42497),
            .in2(N__38367),
            .in3(N__42263),
            .lcout(\c0.n10_adj_4313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1682_LC_11_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1682_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1682_LC_11_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1682_LC_11_13_5  (
            .in0(N__38185),
            .in1(N__46220),
            .in2(N__38264),
            .in3(N__50621),
            .lcout(\c0.n22617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__3__5434_LC_11_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__3__5434_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__3__5434_LC_11_13_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \c0.data_out_frame_11__3__5434_LC_11_13_6  (
            .in0(N__32853),
            .in1(N__30704),
            .in2(N__48269),
            .in3(N__46097),
            .lcout(data_out_frame_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_11_13_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_11_13_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_11_13_7  (
            .in0(N__34263),
            .in1(N__38029),
            .in2(N__38190),
            .in3(N__37605),
            .lcout(\c0.n22668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1187_LC_11_14_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1187_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1187_LC_11_14_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1187_LC_11_14_0  (
            .in0(N__30690),
            .in1(N__30759),
            .in2(N__41952),
            .in3(N__50620),
            .lcout(\c0.n10_adj_4214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1186_LC_11_14_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1186_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1186_LC_11_14_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1186_LC_11_14_1  (
            .in0(N__50588),
            .in1(N__34344),
            .in2(N__32318),
            .in3(N__38092),
            .lcout(\c0.n22534 ),
            .ltout(\c0.n22534_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__2__5299_LC_11_14_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__2__5299_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__2__5299_LC_11_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__2__5299_LC_11_14_2  (
            .in0(N__30824),
            .in1(N__41657),
            .in2(N__30831),
            .in3(N__30855),
            .lcout(\c0.data_out_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78609),
            .ce(N__45042),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1180_LC_11_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1180_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1180_LC_11_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1180_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__46883),
            .in2(_gnd_net_),
            .in3(N__41564),
            .lcout(\c0.n20415 ),
            .ltout(\c0.n20415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_11_14_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_11_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_LC_11_14_5  (
            .in0(N__37137),
            .in1(N__41370),
            .in2(N__30828),
            .in3(N__34367),
            .lcout(\c0.n24530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1661_LC_11_14_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1661_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1661_LC_11_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1661_LC_11_14_6  (
            .in0(N__30823),
            .in1(N__32028),
            .in2(N__33996),
            .in3(N__32349),
            .lcout(\c0.n22414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1188_LC_11_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1188_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1188_LC_11_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1188_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__38091),
            .in2(_gnd_net_),
            .in3(N__46599),
            .lcout(\c0.n20384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__5__5296_LC_11_15_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__5__5296_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__5__5296_LC_11_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__5__5296_LC_11_15_0  (
            .in0(N__30774),
            .in1(N__30809),
            .in2(N__46140),
            .in3(N__41639),
            .lcout(\c0.data_out_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78600),
            .ce(N__45043),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_11_15_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_11_15_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_11_15_1  (
            .in0(N__43233),
            .in1(_gnd_net_),
            .in2(N__30795),
            .in3(N__34467),
            .lcout(\c0.n26_adj_4680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1633_LC_11_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1633_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1633_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1633_LC_11_15_2  (
            .in0(N__37139),
            .in1(N__41431),
            .in2(_gnd_net_),
            .in3(N__30845),
            .lcout(\c0.n21496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1226_LC_11_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1226_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1226_LC_11_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1226_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__46134),
            .in2(_gnd_net_),
            .in3(N__30773),
            .lcout(n22735),
            .ltout(n22735_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i21229_4_lut_LC_11_15_4.C_ON=1'b0;
    defparam i21229_4_lut_LC_11_15_4.SEQ_MODE=4'b0000;
    defparam i21229_4_lut_LC_11_15_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 i21229_4_lut_LC_11_15_4 (
            .in0(N__30861),
            .in1(N__37535),
            .in2(N__30876),
            .in3(N__34345),
            .lcout(n24904),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1825_LC_11_15_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1825_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1825_LC_11_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1825_LC_11_15_5  (
            .in0(N__30846),
            .in1(N__46135),
            .in2(N__30873),
            .in3(N__32301),
            .lcout(),
            .ltout(\c0.n20_adj_4699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__0__5293_LC_11_15_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__0__5293_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__0__5293_LC_11_15_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.data_out_frame_29__0__5293_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__50505),
            .in2(N__30864),
            .in3(N__41850),
            .lcout(\c0.data_out_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78600),
            .ce(N__45043),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1229_LC_11_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1229_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1229_LC_11_16_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1229_LC_11_16_0  (
            .in0(N__46609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41562),
            .lcout(n22285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_11_16_1 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_11_16_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_11_16_1  (
            .in0(N__47179),
            .in1(N__47098),
            .in2(_gnd_net_),
            .in3(N__47149),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78591),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1601_LC_11_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1601_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1601_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1601_LC_11_16_3  (
            .in0(N__50650),
            .in1(N__38093),
            .in2(_gnd_net_),
            .in3(N__46608),
            .lcout(\c0.n22330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i7_LC_11_16_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i7_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i7_LC_11_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i7_LC_11_16_4  (
            .in0(N__40567),
            .in1(N__32535),
            .in2(_gnd_net_),
            .in3(N__34594),
            .lcout(encoder1_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78591),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_2035_LC_11_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_2035_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_2035_LC_11_16_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_2035_LC_11_16_5  (
            .in0(N__41563),
            .in1(N__41432),
            .in2(_gnd_net_),
            .in3(N__38094),
            .lcout(\c0.n6_adj_4210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1808_LC_11_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1808_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1808_LC_11_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1808_LC_11_16_7  (
            .in0(N__46800),
            .in1(N__41366),
            .in2(_gnd_net_),
            .in3(N__46391),
            .lcout(\c0.n13683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i15_LC_11_17_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i15_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i15_LC_11_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i15_LC_11_17_0  (
            .in0(N__40535),
            .in1(N__32625),
            .in2(_gnd_net_),
            .in3(N__34963),
            .lcout(encoder1_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__3__5442_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__3__5442_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__3__5442_LC_11_17_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__3__5442_LC_11_17_1  (
            .in0(N__48319),
            .in1(N__46056),
            .in2(N__34899),
            .in3(N__30962),
            .lcout(data_out_frame_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1185_LC_11_17_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1185_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1185_LC_11_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1185_LC_11_17_2  (
            .in0(N__41230),
            .in1(N__41429),
            .in2(N__30948),
            .in3(N__37742),
            .lcout(\c0.n20641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i3_LC_11_17_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i3_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i3_LC_11_17_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i3_LC_11_17_3  (
            .in0(N__32595),
            .in1(N__40536),
            .in2(_gnd_net_),
            .in3(N__45479),
            .lcout(encoder1_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__6__5431_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__6__5431_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__6__5431_LC_11_17_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_11__6__5431_LC_11_17_4  (
            .in0(N__46055),
            .in1(N__48322),
            .in2(N__34655),
            .in3(N__31532),
            .lcout(data_out_frame_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__2__5459_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__2__5459_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__2__5459_LC_11_17_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__2__5459_LC_11_17_5  (
            .in0(N__48321),
            .in1(N__46057),
            .in2(N__36622),
            .in3(N__31058),
            .lcout(data_out_frame_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_17_6  (
            .in0(N__33185),
            .in1(N__30911),
            .in2(_gnd_net_),
            .in3(N__43234),
            .lcout(\c0.n11_adj_4572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__0__5421_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__0__5421_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__0__5421_LC_11_17_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_frame_13__0__5421_LC_11_17_7  (
            .in0(N__48320),
            .in1(N__33953),
            .in2(N__30915),
            .in3(N__46058),
            .lcout(data_out_frame_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_11_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_11_18_0  (
            .in0(N__34548),
            .in1(N__30903),
            .in2(_gnd_net_),
            .in3(N__43216),
            .lcout(),
            .ltout(\c0.n5_adj_4650_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21042_4_lut_LC_11_18_1 .C_ON=1'b0;
    defparam \c0.i21042_4_lut_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21042_4_lut_LC_11_18_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.i21042_4_lut_LC_11_18_1  (
            .in0(N__40773),
            .in1(N__41019),
            .in2(N__30888),
            .in3(N__30885),
            .lcout(\c0.n24809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21036_4_lut_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.i21036_4_lut_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21036_4_lut_LC_11_18_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i21036_4_lut_LC_11_18_2  (
            .in0(N__41020),
            .in1(N__32487),
            .in2(N__31083),
            .in3(N__40774),
            .lcout(\c0.n24803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25056_bdd_4_lut_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.n25056_bdd_4_lut_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.n25056_bdd_4_lut_LC_11_18_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n25056_bdd_4_lut_LC_11_18_3  (
            .in0(N__40775),
            .in1(N__33342),
            .in2(N__31059),
            .in3(N__30972),
            .lcout(),
            .ltout(\c0.n25059_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21236_4_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.i21236_4_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21236_4_lut_LC_11_18_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.i21236_4_lut_LC_11_18_4  (
            .in0(N__41021),
            .in1(N__32427),
            .in2(N__31044),
            .in3(N__40776),
            .lcout(),
            .ltout(n25004_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2061_LC_11_18_5.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2061_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2061_LC_11_18_5.LUT_INIT=16'b1100110011100100;
    LogicCell40 i24_3_lut_4_lut_adj_2061_LC_11_18_5 (
            .in0(N__31189),
            .in1(N__31023),
            .in2(N__31041),
            .in3(N__31317),
            .lcout(n10_adj_4778),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21044_4_lut_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.i21044_4_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21044_4_lut_LC_11_19_0 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.i21044_4_lut_LC_11_19_0  (
            .in0(N__32409),
            .in1(N__31029),
            .in2(N__31395),
            .in3(N__31312),
            .lcout(n24811),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__3__5298_LC_11_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__3__5298_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__3__5298_LC_11_19_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_28__3__5298_LC_11_19_1  (
            .in0(N__46019),
            .in1(N__48252),
            .in2(N__31005),
            .in3(N__31017),
            .lcout(data_out_frame_28_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21338_LC_11_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21338_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21338_LC_11_19_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_21338_LC_11_19_2  (
            .in0(N__33269),
            .in1(N__40772),
            .in2(N__31446),
            .in3(N__43176),
            .lcout(),
            .ltout(\c0.n25110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25110_bdd_4_lut_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.n25110_bdd_4_lut_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.n25110_bdd_4_lut_LC_11_19_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n25110_bdd_4_lut_LC_11_19_3  (
            .in0(N__35226),
            .in1(N__34695),
            .in2(N__30981),
            .in3(N__40805),
            .lcout(\c0.n25113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21313_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21313_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21313_LC_11_19_5 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_21313_LC_11_19_5  (
            .in0(N__43177),
            .in1(N__31457),
            .in2(N__32913),
            .in3(N__40804),
            .lcout(\c0.n25056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__2__5443_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__2__5443_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__2__5443_LC_11_19_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_10__2__5443_LC_11_19_6  (
            .in0(N__48250),
            .in1(N__31458),
            .in2(N__38366),
            .in3(N__46020),
            .lcout(data_out_frame_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__0__5437_LC_11_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__0__5437_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__0__5437_LC_11_19_7 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_11__0__5437_LC_11_19_7  (
            .in0(N__46018),
            .in1(N__48251),
            .in2(N__34073),
            .in3(N__31445),
            .lcout(data_out_frame_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78601),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i12_LC_11_20_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i12_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i12_LC_11_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i12_LC_11_20_1  (
            .in0(N__47653),
            .in1(N__36453),
            .in2(_gnd_net_),
            .in3(N__36487),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78610),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__5__5480_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__5__5480_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__5__5480_LC_11_20_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_out_frame_5__5__5480_LC_11_20_2  (
            .in0(N__47064),
            .in1(N__46023),
            .in2(N__31497),
            .in3(N__48256),
            .lcout(data_out_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78610),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21244_4_lut_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.i21244_4_lut_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i21244_4_lut_LC_11_20_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.i21244_4_lut_LC_11_20_3  (
            .in0(N__40778),
            .in1(N__31515),
            .in2(N__31434),
            .in3(N__41023),
            .lcout(n25012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21178_3_lut_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.i21178_3_lut_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21178_3_lut_LC_11_20_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \c0.i21178_3_lut_LC_11_20_4  (
            .in0(N__41022),
            .in1(N__34995),
            .in2(_gnd_net_),
            .in3(N__43217),
            .lcout(),
            .ltout(\c0.n24945_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21030_4_lut_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.i21030_4_lut_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21030_4_lut_LC_11_20_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i21030_4_lut_LC_11_20_5  (
            .in0(N__40777),
            .in1(N__31464),
            .in2(N__31422),
            .in3(N__41024),
            .lcout(),
            .ltout(\c0.n24797_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21032_4_lut_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.i21032_4_lut_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i21032_4_lut_LC_11_20_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i21032_4_lut_LC_11_20_6  (
            .in0(N__31405),
            .in1(N__41601),
            .in2(N__31332),
            .in3(N__31315),
            .lcout(),
            .ltout(n24799_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2063_LC_11_20_7.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2063_LC_11_20_7.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2063_LC_11_20_7.LUT_INIT=16'b1111010010110000;
    LogicCell40 i24_3_lut_4_lut_adj_2063_LC_11_20_7 (
            .in0(N__31316),
            .in1(N__31190),
            .in2(N__31104),
            .in3(N__31101),
            .lcout(n10_adj_4775),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21328_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21328_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_21328_LC_11_21_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_21328_LC_11_21_0  (
            .in0(N__40769),
            .in1(N__35319),
            .in2(N__31536),
            .in3(N__43085),
            .lcout(),
            .ltout(\c0.n25098_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25098_bdd_4_lut_LC_11_21_1 .C_ON=1'b0;
    defparam \c0.n25098_bdd_4_lut_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.n25098_bdd_4_lut_LC_11_21_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n25098_bdd_4_lut_LC_11_21_1  (
            .in0(N__45699),
            .in1(N__33413),
            .in2(N__31518),
            .in3(N__40771),
            .lcout(\c0.n25101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_21_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_21_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_21_2  (
            .in0(N__35385),
            .in1(N__31505),
            .in2(_gnd_net_),
            .in3(N__43084),
            .lcout(\c0.n5_adj_4679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__5__5472_LC_11_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__5__5472_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__5__5472_LC_11_21_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_6__5__5472_LC_11_21_3  (
            .in0(N__48363),
            .in1(N__45936),
            .in2(N__31509),
            .in3(N__36897),
            .lcout(data_out_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78621),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21247_4_lut_LC_11_21_4 .C_ON=1'b0;
    defparam \c0.i21247_4_lut_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21247_4_lut_LC_11_21_4 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \c0.i21247_4_lut_LC_11_21_4  (
            .in0(N__40768),
            .in1(N__43087),
            .in2(N__41033),
            .in3(N__31493),
            .lcout(),
            .ltout(\c0.n25016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21027_4_lut_LC_11_21_5 .C_ON=1'b0;
    defparam \c0.i21027_4_lut_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21027_4_lut_LC_11_21_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i21027_4_lut_LC_11_21_5  (
            .in0(N__40994),
            .in1(N__31482),
            .in2(N__31476),
            .in3(N__40770),
            .lcout(\c0.n24794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_11_21_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_11_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_11_21_7  (
            .in0(N__43086),
            .in1(N__35487),
            .in2(_gnd_net_),
            .in3(N__33398),
            .lcout(\c0.n5_adj_4700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1849_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1849_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1849_LC_11_22_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1849_LC_11_22_0  (
            .in0(N__39257),
            .in1(N__43825),
            .in2(N__43708),
            .in3(N__43654),
            .lcout(\c0.n4_adj_4678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_11_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_11_22_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i23_LC_11_22_1  (
            .in0(N__50466),
            .in1(N__44499),
            .in2(_gnd_net_),
            .in3(N__38868),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78633),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21170_3_lut_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.rx.i21170_3_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21170_3_lut_LC_11_22_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i21170_3_lut_LC_11_22_4  (
            .in0(N__50044),
            .in1(N__31907),
            .in2(_gnd_net_),
            .in3(N__31654),
            .lcout(n24922),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_105_i4_2_lut_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.rx.equal_105_i4_2_lut_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_105_i4_2_lut_LC_11_22_5 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \c0.rx.equal_105_i4_2_lut_LC_11_22_5  (
            .in0(N__49722),
            .in1(N__49634),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n4_adj_4761),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1944_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1944_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1944_LC_11_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_1944_LC_11_22_6  (
            .in0(N__39756),
            .in1(N__33552),
            .in2(N__36099),
            .in3(N__49047),
            .lcout(\c0.n24255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1936_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1936_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1936_LC_11_23_1 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1936_LC_11_23_1  (
            .in0(N__35779),
            .in1(N__44196),
            .in2(N__35908),
            .in3(N__38934),
            .lcout(\c0.n21583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1842_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1842_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1842_LC_11_23_2 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1842_LC_11_23_2  (
            .in0(N__44056),
            .in1(N__44087),
            .in2(N__43997),
            .in3(N__43526),
            .lcout(\c0.n13056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1956_LC_11_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1956_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1956_LC_11_23_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1956_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__31592),
            .in2(_gnd_net_),
            .in3(N__31563),
            .lcout(\c0.n14530 ),
            .ltout(\c0.n14530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_1964_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1964_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1964_LC_11_23_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1964_LC_11_23_4  (
            .in0(N__35897),
            .in1(N__36265),
            .in2(N__31539),
            .in3(N__36003),
            .lcout(\c0.n6_adj_4495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2004_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2004_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2004_LC_11_23_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_2004_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__33593),
            .in2(_gnd_net_),
            .in3(N__33543),
            .lcout(\c0.n14784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_2_lut_3_lut_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.rx.i3_2_lut_3_lut_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_2_lut_3_lut_LC_11_24_0 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \c0.rx.i3_2_lut_3_lut_LC_11_24_0  (
            .in0(N__31976),
            .in1(_gnd_net_),
            .in2(N__32007),
            .in3(N__31900),
            .lcout(),
            .ltout(\c0.rx.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5_4_lut_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.rx.i5_4_lut_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5_4_lut_LC_11_24_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.rx.i5_4_lut_LC_11_24_1  (
            .in0(N__31776),
            .in1(N__31953),
            .in2(N__31695),
            .in3(N__31812),
            .lcout(\c0.rx.r_SM_Main_2_N_3686_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1957_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1957_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1957_LC_11_24_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1957_LC_11_24_2  (
            .in0(N__36212),
            .in1(N__48420),
            .in2(_gnd_net_),
            .in3(N__31687),
            .lcout(\c0.n22131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2007_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2007_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2007_LC_11_24_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_2007_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__36170),
            .in2(_gnd_net_),
            .in3(N__35544),
            .lcout(\c0.n14721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13988_2_lut_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.rx.i13988_2_lut_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13988_2_lut_LC_11_24_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.i13988_2_lut_LC_11_24_4  (
            .in0(N__31749),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31775),
            .lcout(\c0.rx.n17590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13930_2_lut_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.rx.i13930_2_lut_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13930_2_lut_LC_11_24_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i13930_2_lut_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__31975),
            .in2(_gnd_net_),
            .in3(N__32003),
            .lcout(),
            .ltout(\c0.rx.n17531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_11_24_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \c0.rx.i2_4_lut_LC_11_24_6  (
            .in0(N__31722),
            .in1(N__31948),
            .in2(N__31671),
            .in3(N__31668),
            .lcout(\c0.rx.n17848 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5_3_lut_LC_11_24_7 .C_ON=1'b0;
    defparam \c0.rx.i5_3_lut_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5_3_lut_LC_11_24_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.rx.i5_3_lut_LC_11_24_7  (
            .in0(N__31949),
            .in1(N__31977),
            .in2(_gnd_net_),
            .in3(N__31805),
            .lcout(\c0.rx.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i20933_3_lut_LC_11_25_0 .C_ON=1'b0;
    defparam \c0.rx.i20933_3_lut_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i20933_3_lut_LC_11_25_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.rx.i20933_3_lut_LC_11_25_0  (
            .in0(N__39300),
            .in1(N__50865),
            .in2(_gnd_net_),
            .in3(N__31894),
            .lcout(),
            .ltout(\c0.rx.n24697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21217_4_lut_LC_11_25_1 .C_ON=1'b0;
    defparam \c0.rx.i21217_4_lut_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21217_4_lut_LC_11_25_1 .LUT_INIT=16'b0101110101010101;
    LogicCell40 \c0.rx.i21217_4_lut_LC_11_25_1  (
            .in0(N__50042),
            .in1(N__31626),
            .in2(N__31620),
            .in3(N__31818),
            .lcout(),
            .ltout(\c0.rx.n24914_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_11_25_2 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \c0.rx.i1_4_lut_LC_11_25_2  (
            .in0(N__50106),
            .in1(N__49957),
            .in2(N__31617),
            .in3(N__42017),
            .lcout(n14895),
            .ltout(n14895_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_11_25_3 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_11_25_3  (
            .in0(N__31804),
            .in1(N__31785),
            .in2(N__31833),
            .in3(N__39275),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21223_3_lut_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.rx.i21223_3_lut_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21223_3_lut_LC_11_25_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.rx.i21223_3_lut_LC_11_25_4  (
            .in0(N__39301),
            .in1(N__50043),
            .in2(_gnd_net_),
            .in3(N__50866),
            .lcout(),
            .ltout(n24921_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_11_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_11_25_5 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_11_25_5  (
            .in0(N__49958),
            .in1(N__50107),
            .in2(N__31830),
            .in3(N__31827),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21234_4_lut_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.rx.i21234_4_lut_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21234_4_lut_LC_11_25_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.rx.i21234_4_lut_LC_11_25_6  (
            .in0(N__31747),
            .in1(N__31773),
            .in2(N__31721),
            .in3(N__32001),
            .lcout(\c0.rx.n24916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_11_25_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.rx.i2_3_lut_LC_11_25_7  (
            .in0(N__31803),
            .in1(N__31713),
            .in2(_gnd_net_),
            .in3(N__31746),
            .lcout(\c0.rx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_11_26_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_11_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_2_lut_LC_11_26_0  (
            .in0(_gnd_net_),
            .in1(N__31806),
            .in2(_gnd_net_),
            .in3(N__31779),
            .lcout(n226),
            .ltout(),
            .carryin(bfn_11_26_0_),
            .carryout(\c0.rx.n19716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_11_26_1 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i1_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_11_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_11_26_1  (
            .in0(_gnd_net_),
            .in1(N__31774),
            .in2(_gnd_net_),
            .in3(N__31752),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.rx.n19716 ),
            .carryout(\c0.rx.n19717 ),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.rx.r_Clock_Count__i2_LC_11_26_2 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i2_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_11_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_11_26_2  (
            .in0(_gnd_net_),
            .in1(N__31748),
            .in2(_gnd_net_),
            .in3(N__31725),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.rx.n19717 ),
            .carryout(\c0.rx.n19718 ),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.rx.r_Clock_Count__i3_LC_11_26_3 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i3_LC_11_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_11_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__31720),
            .in2(_gnd_net_),
            .in3(N__32010),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.rx.n19718 ),
            .carryout(\c0.rx.n19719 ),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.rx.r_Clock_Count__i4_LC_11_26_4 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i4_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_11_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_11_26_4  (
            .in0(_gnd_net_),
            .in1(N__32002),
            .in2(_gnd_net_),
            .in3(N__31980),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.rx.n19719 ),
            .carryout(\c0.rx.n19720 ),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.rx.r_Clock_Count__i5_LC_11_26_5 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i5_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_11_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(N__31974),
            .in2(_gnd_net_),
            .in3(N__31956),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.rx.n19720 ),
            .carryout(\c0.rx.n19721 ),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.rx.r_Clock_Count__i6_LC_11_26_6 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i6_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_11_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_11_26_6  (
            .in0(_gnd_net_),
            .in1(N__31947),
            .in2(_gnd_net_),
            .in3(N__31923),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.rx.n19721 ),
            .carryout(\c0.rx.n19722 ),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.rx.r_Clock_Count__i7_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_11_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(N__31898),
            .in2(_gnd_net_),
            .in3(N__31920),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78689),
            .ce(N__39279),
            .sr(N__31857));
    defparam \c0.FRAME_MATCHER_state_i4_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_11_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_11_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_11_27_0  (
            .in0(_gnd_net_),
            .in1(N__36031),
            .in2(_gnd_net_),
            .in3(N__48992),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78702),
            .ce(),
            .sr(N__33480));
    defparam \c0.i1_2_lut_adj_1986_LC_12_7_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1986_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1986_LC_12_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1986_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__49102),
            .in2(_gnd_net_),
            .in3(N__47836),
            .lcout(\c0.n21645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1351_LC_12_8_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1351_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1351_LC_12_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1351_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__36421),
            .in2(_gnd_net_),
            .in3(N__36341),
            .lcout(\c0.n22638 ),
            .ltout(\c0.n22638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1760_LC_12_8_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1760_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1760_LC_12_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1760_LC_12_8_5  (
            .in0(N__36964),
            .in1(N__39613),
            .in2(N__31836),
            .in3(N__44708),
            .lcout(\c0.n6_adj_4336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1254_LC_12_8_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1254_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1254_LC_12_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1254_LC_12_8_7  (
            .in0(N__33891),
            .in1(N__33869),
            .in2(_gnd_net_),
            .in3(N__34028),
            .lcout(\c0.n20333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.encoder0_position_29__I_0_2_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \c0.encoder0_position_29__I_0_2_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.encoder0_position_29__I_0_2_lut_LC_12_9_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.encoder0_position_29__I_0_2_lut_LC_12_9_1  (
            .in0(N__36874),
            .in1(_gnd_net_),
            .in2(N__36975),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_frame_29__7__N_855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1404_LC_12_9_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1404_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1404_LC_12_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1404_LC_12_9_2  (
            .in0(N__34011),
            .in1(N__33852),
            .in2(_gnd_net_),
            .in3(N__42330),
            .lcout(\c0.n21323 ),
            .ltout(\c0.n21323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1266_LC_12_9_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1266_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1266_LC_12_9_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1266_LC_12_9_3  (
            .in0(N__34746),
            .in1(_gnd_net_),
            .in2(N__32052),
            .in3(N__38122),
            .lcout(\c0.n21406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1314_LC_12_9_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1314_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1314_LC_12_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1314_LC_12_9_4  (
            .in0(N__32848),
            .in1(N__36342),
            .in2(_gnd_net_),
            .in3(N__36872),
            .lcout(\c0.n22608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1386_LC_12_9_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1386_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1386_LC_12_9_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1386_LC_12_9_5  (
            .in0(N__44382),
            .in1(N__37899),
            .in2(N__36974),
            .in3(N__32049),
            .lcout(\c0.n12488 ),
            .ltout(\c0.n12488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1750_LC_12_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1750_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1750_LC_12_9_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1750_LC_12_9_6  (
            .in0(N__45591),
            .in1(_gnd_net_),
            .in2(N__32043),
            .in3(N__36873),
            .lcout(\c0.n20449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1354_LC_12_9_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1354_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1354_LC_12_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1354_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__35188),
            .in2(_gnd_net_),
            .in3(N__36422),
            .lcout(\c0.n22791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_2015_LC_12_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_2015_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_2015_LC_12_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_2015_LC_12_10_1  (
            .in0(N__35111),
            .in1(N__32040),
            .in2(_gnd_net_),
            .in3(N__34136),
            .lcout(\c0.n13531 ),
            .ltout(\c0.n13531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1332_LC_12_10_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1332_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1332_LC_12_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1332_LC_12_10_2  (
            .in0(N__41752),
            .in1(N__38551),
            .in2(N__32031),
            .in3(N__32021),
            .lcout(\c0.n29_adj_4329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1322_LC_12_10_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1322_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1322_LC_12_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1322_LC_12_10_3  (
            .in0(N__36697),
            .in1(N__35353),
            .in2(_gnd_net_),
            .in3(N__42552),
            .lcout(),
            .ltout(\c0.n14_adj_4317_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1324_LC_12_10_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1324_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1324_LC_12_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1324_LC_12_10_4  (
            .in0(N__44349),
            .in1(N__32073),
            .in2(N__32067),
            .in3(N__32064),
            .lcout(\c0.n20388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1323_LC_12_10_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1323_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1323_LC_12_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1323_LC_12_10_5  (
            .in0(N__34181),
            .in1(N__39553),
            .in2(N__42174),
            .in3(N__34027),
            .lcout(\c0.n15_adj_4318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1334_LC_12_10_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1334_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1334_LC_12_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1334_LC_12_10_6  (
            .in0(N__34137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38552),
            .lcout(\c0.n6_adj_4330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1335_LC_12_11_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1335_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1335_LC_12_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1335_LC_12_11_0  (
            .in0(N__39915),
            .in1(N__32058),
            .in2(N__44432),
            .in3(N__42400),
            .lcout(\c0.n20348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_2010_LC_12_11_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_2010_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_2010_LC_12_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_2010_LC_12_11_1  (
            .in0(N__39875),
            .in1(N__37035),
            .in2(_gnd_net_),
            .in3(N__41318),
            .lcout(\c0.n20_adj_4321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i19_LC_12_11_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i19_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i19_LC_12_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i19_LC_12_11_2  (
            .in0(N__32847),
            .in1(N__32820),
            .in2(_gnd_net_),
            .in3(N__40528),
            .lcout(encoder1_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78658),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i11_LC_12_11_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i11_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i11_LC_12_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i11_LC_12_11_3  (
            .in0(N__47654),
            .in1(N__36522),
            .in2(_gnd_net_),
            .in3(N__36547),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78658),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i28_LC_12_11_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i28_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i28_LC_12_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i28_LC_12_11_4  (
            .in0(N__36957),
            .in1(N__36912),
            .in2(_gnd_net_),
            .in3(N__47656),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78658),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i12_LC_12_11_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i12_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i12_LC_12_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i12_LC_12_11_5  (
            .in0(N__40527),
            .in1(N__32730),
            .in2(_gnd_net_),
            .in3(N__41760),
            .lcout(encoder1_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78658),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i26_LC_12_11_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i26_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i26_LC_12_11_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \quad_counter0.count_i0_i26_LC_12_11_6  (
            .in0(N__37008),
            .in1(_gnd_net_),
            .in2(N__37045),
            .in3(N__47655),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78658),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i4_LC_12_12_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i4_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i4_LC_12_12_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i4_LC_12_12_1  (
            .in0(N__32580),
            .in1(N__40543),
            .in2(_gnd_net_),
            .in3(N__35268),
            .lcout(encoder1_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1303_LC_12_12_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1303_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1303_LC_12_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1303_LC_12_12_2  (
            .in0(N__34895),
            .in1(N__34316),
            .in2(_gnd_net_),
            .in3(N__42498),
            .lcout(\c0.n20367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1353_LC_12_12_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1353_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1353_LC_12_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1353_LC_12_12_3  (
            .in0(N__32112),
            .in1(N__47485),
            .in2(N__32889),
            .in3(N__32103),
            .lcout(\c0.n13395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25062_bdd_4_lut_4_lut_LC_12_12_4 .C_ON=1'b0;
    defparam \c0.n25062_bdd_4_lut_4_lut_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.n25062_bdd_4_lut_4_lut_LC_12_12_4 .LUT_INIT=16'b1100110010011000;
    LogicCell40 \c0.n25062_bdd_4_lut_4_lut_LC_12_12_4  (
            .in0(N__41053),
            .in1(N__40599),
            .in2(N__33369),
            .in3(N__43238),
            .lcout(n25065),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i6_LC_12_12_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i6_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i6_LC_12_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i6_LC_12_12_5  (
            .in0(N__40541),
            .in1(N__32550),
            .in2(_gnd_net_),
            .in3(N__34421),
            .lcout(encoder1_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78647),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i20_LC_12_12_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i20_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i20_LC_12_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i20_LC_12_12_6  (
            .in0(N__40542),
            .in1(N__32805),
            .in2(_gnd_net_),
            .in3(N__33798),
            .lcout(encoder1_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78647),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i0_LC_12_12_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i0_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i0_LC_12_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i0_LC_12_12_7  (
            .in0(N__40540),
            .in1(N__32382),
            .in2(_gnd_net_),
            .in3(N__33942),
            .lcout(encoder1_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1524_LC_12_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1524_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1524_LC_12_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1524_LC_12_13_0  (
            .in0(N__44626),
            .in1(N__35261),
            .in2(N__41172),
            .in3(N__34814),
            .lcout(\c0.n10500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_4_lut_LC_12_13_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_4_lut_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_4_lut_LC_12_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_3_lut_4_lut_LC_12_13_1  (
            .in0(N__34815),
            .in1(N__46877),
            .in2(N__35283),
            .in3(N__44627),
            .lcout(\c0.n9_adj_4562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1811_LC_12_13_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1811_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1811_LC_12_13_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1811_LC_12_13_2  (
            .in0(N__32234),
            .in1(N__32344),
            .in2(N__32319),
            .in3(N__32274),
            .lcout(\c0.n12_adj_4688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1815_LC_12_13_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1815_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1815_LC_12_13_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1815_LC_12_13_3  (
            .in0(N__32297),
            .in1(N__46696),
            .in2(N__46395),
            .in3(N__34449),
            .lcout(),
            .ltout(\c0.n10_adj_4690_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1814_LC_12_13_4 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1814_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1814_LC_12_13_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_adj_1814_LC_12_13_4  (
            .in0(N__32286),
            .in1(N__34352),
            .in2(N__32277),
            .in3(N__37091),
            .lcout(\c0.n22710 ),
            .ltout(\c0.n22710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1793_LC_12_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1793_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1793_LC_12_13_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1793_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32268),
            .in3(N__32265),
            .lcout(),
            .ltout(\c0.n6_adj_4683_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__6__5287_LC_12_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__6__5287_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__6__5287_LC_12_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_29__6__5287_LC_12_13_6  (
            .in0(N__32235),
            .in1(N__37779),
            .in2(N__32208),
            .in3(N__32175),
            .lcout(\c0.data_out_frame_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78634),
            .ce(N__45054),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1810_LC_12_14_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1810_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1810_LC_12_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1810_LC_12_14_0  (
            .in0(N__32168),
            .in1(N__46557),
            .in2(N__32205),
            .in3(N__32181),
            .lcout(\c0.n20360 ),
            .ltout(\c0.n20360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__7__5286_LC_12_14_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__7__5286_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__7__5286_LC_12_14_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.data_out_frame_29__7__5286_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__32169),
            .in2(N__32160),
            .in3(N__38030),
            .lcout(\c0.data_out_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78622),
            .ce(N__45035),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_12_14_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_12_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_12_14_2  (
            .in0(N__43231),
            .in1(N__32157),
            .in2(_gnd_net_),
            .in3(N__41472),
            .lcout(\c0.n26_adj_4713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_12_14_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_12_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_12_14_3  (
            .in0(N__33234),
            .in1(N__32498),
            .in2(_gnd_net_),
            .in3(N__43229),
            .lcout(\c0.n5_adj_4567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_12_14_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_12_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_12_14_4  (
            .in0(N__43227),
            .in1(N__32475),
            .in2(_gnd_net_),
            .in3(N__33171),
            .lcout(\c0.n11_adj_4646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_12_14_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_12_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_12_14_5  (
            .in0(N__34842),
            .in1(N__41283),
            .in2(_gnd_net_),
            .in3(N__43230),
            .lcout(\c0.n5_adj_4644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_12_14_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_12_14_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_12_14_6  (
            .in0(N__43232),
            .in1(_gnd_net_),
            .in2(N__35064),
            .in3(N__33315),
            .lcout(\c0.n11_adj_4652 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_12_14_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_12_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_12_14_7  (
            .in0(N__41262),
            .in1(N__32415),
            .in2(_gnd_net_),
            .in3(N__43228),
            .lcout(\c0.n26_adj_4651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_1_LC_12_15_0 .C_ON=1'b1;
    defparam \quad_counter1.add_613_1_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_1_LC_12_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter1.add_613_1_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__32995),
            .in2(N__33074),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\quad_counter1.n19731 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_2_lut_LC_12_15_1 .C_ON=1'b1;
    defparam \quad_counter1.add_613_2_lut_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_2_lut_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_2_lut_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__33946),
            .in2(N__32394),
            .in3(N__32370),
            .lcout(n2291),
            .ltout(),
            .carryin(\quad_counter1.n19731 ),
            .carryout(\quad_counter1.n19732 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_3_lut_LC_12_15_2 .C_ON=1'b1;
    defparam \quad_counter1.add_613_3_lut_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_3_lut_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_3_lut_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__34775),
            .in2(N__33075),
            .in3(N__32352),
            .lcout(n2290),
            .ltout(),
            .carryin(\quad_counter1.n19732 ),
            .carryout(\quad_counter1.n19733 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_4_lut_LC_12_15_3 .C_ON=1'b1;
    defparam \quad_counter1.add_613_4_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_4_lut_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_4_lut_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__46329),
            .in2(N__33071),
            .in3(N__32598),
            .lcout(n2289),
            .ltout(),
            .carryin(\quad_counter1.n19733 ),
            .carryout(\quad_counter1.n19734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_5_lut_LC_12_15_4 .C_ON=1'b1;
    defparam \quad_counter1.add_613_5_lut_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_5_lut_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_5_lut_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__45493),
            .in2(N__33076),
            .in3(N__32583),
            .lcout(n2288),
            .ltout(),
            .carryin(\quad_counter1.n19734 ),
            .carryout(\quad_counter1.n19735 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_6_lut_LC_12_15_5 .C_ON=1'b1;
    defparam \quad_counter1.add_613_6_lut_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_6_lut_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_6_lut_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__35284),
            .in2(N__33072),
            .in3(N__32571),
            .lcout(n2287),
            .ltout(),
            .carryin(\quad_counter1.n19735 ),
            .carryout(\quad_counter1.n19736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_7_lut_LC_12_15_6 .C_ON=1'b1;
    defparam \quad_counter1.add_613_7_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_7_lut_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_7_lut_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__41185),
            .in2(N__33077),
            .in3(N__32553),
            .lcout(n2286),
            .ltout(),
            .carryin(\quad_counter1.n19736 ),
            .carryout(\quad_counter1.n19737 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_8_lut_LC_12_15_7 .C_ON=1'b1;
    defparam \quad_counter1.add_613_8_lut_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_8_lut_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_8_lut_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__34425),
            .in2(N__33073),
            .in3(N__32538),
            .lcout(n2285),
            .ltout(),
            .carryin(\quad_counter1.n19737 ),
            .carryout(\quad_counter1.n19738 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_9_lut_LC_12_16_0 .C_ON=1'b1;
    defparam \quad_counter1.add_613_9_lut_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_9_lut_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_9_lut_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__34593),
            .in2(N__33129),
            .in3(N__32529),
            .lcout(n2284),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\quad_counter1.n19739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_10_lut_LC_12_16_1 .C_ON=1'b1;
    defparam \quad_counter1.add_613_10_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_10_lut_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_10_lut_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__33081),
            .in2(N__40174),
            .in3(N__32526),
            .lcout(n2283),
            .ltout(),
            .carryin(\quad_counter1.n19739 ),
            .carryout(\quad_counter1.n19740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_11_lut_LC_12_16_2 .C_ON=1'b1;
    defparam \quad_counter1.add_613_11_lut_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_11_lut_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_11_lut_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__40084),
            .in2(N__33130),
            .in3(N__32508),
            .lcout(n2282),
            .ltout(),
            .carryin(\quad_counter1.n19740 ),
            .carryout(\quad_counter1.n19741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_12_lut_LC_12_16_3 .C_ON=1'b1;
    defparam \quad_counter1.add_613_12_lut_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_12_lut_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_12_lut_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__33085),
            .in2(N__35038),
            .in3(N__32505),
            .lcout(n2281),
            .ltout(),
            .carryin(\quad_counter1.n19741 ),
            .carryout(\quad_counter1.n19742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_13_lut_LC_12_16_4 .C_ON=1'b1;
    defparam \quad_counter1.add_613_13_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_13_lut_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_13_lut_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__35132),
            .in2(N__33131),
            .in3(N__32733),
            .lcout(n2280),
            .ltout(),
            .carryin(\quad_counter1.n19742 ),
            .carryout(\quad_counter1.n19743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_14_lut_LC_12_16_5 .C_ON=1'b1;
    defparam \quad_counter1.add_613_14_lut_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_14_lut_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_14_lut_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__33089),
            .in2(N__41780),
            .in3(N__32718),
            .lcout(n2279),
            .ltout(),
            .carryin(\quad_counter1.n19743 ),
            .carryout(\quad_counter1.n19744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_15_lut_LC_12_16_6 .C_ON=1'b1;
    defparam \quad_counter1.add_613_15_lut_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_15_lut_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_15_lut_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__32711),
            .in2(N__33132),
            .in3(N__32646),
            .lcout(n2278),
            .ltout(),
            .carryin(\quad_counter1.n19744 ),
            .carryout(\quad_counter1.n19745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_16_lut_LC_12_16_7 .C_ON=1'b1;
    defparam \quad_counter1.add_613_16_lut_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_16_lut_LC_12_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_16_lut_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__33093),
            .in2(N__33701),
            .in3(N__32628),
            .lcout(n2277),
            .ltout(),
            .carryin(\quad_counter1.n19745 ),
            .carryout(\quad_counter1.n19746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_17_lut_LC_12_17_0 .C_ON=1'b1;
    defparam \quad_counter1.add_613_17_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_17_lut_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_17_lut_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__34959),
            .in2(N__33133),
            .in3(N__32619),
            .lcout(n2276),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\quad_counter1.n19747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_18_lut_LC_12_17_1 .C_ON=1'b1;
    defparam \quad_counter1.add_613_18_lut_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_18_lut_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_18_lut_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__33097),
            .in2(N__34083),
            .in3(N__32616),
            .lcout(n2275),
            .ltout(),
            .carryin(\quad_counter1.n19747 ),
            .carryout(\quad_counter1.n19748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_19_lut_LC_12_17_2 .C_ON=1'b1;
    defparam \quad_counter1.add_613_19_lut_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_19_lut_LC_12_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_19_lut_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__35207),
            .in2(N__33134),
            .in3(N__32613),
            .lcout(n2274),
            .ltout(),
            .carryin(\quad_counter1.n19748 ),
            .carryout(\quad_counter1.n19749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_20_lut_LC_12_17_3 .C_ON=1'b1;
    defparam \quad_counter1.add_613_20_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_20_lut_LC_12_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_20_lut_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__33101),
            .in2(N__32888),
            .in3(N__32610),
            .lcout(n2273),
            .ltout(),
            .carryin(\quad_counter1.n19749 ),
            .carryout(\quad_counter1.n19750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_21_lut_LC_12_17_4 .C_ON=1'b1;
    defparam \quad_counter1.add_613_21_lut_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_21_lut_LC_12_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_21_lut_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__32849),
            .in2(N__33135),
            .in3(N__32808),
            .lcout(n2272),
            .ltout(),
            .carryin(\quad_counter1.n19750 ),
            .carryout(\quad_counter1.n19751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_22_lut_LC_12_17_5 .C_ON=1'b1;
    defparam \quad_counter1.add_613_22_lut_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_22_lut_LC_12_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_22_lut_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__33105),
            .in2(N__33806),
            .in3(N__32796),
            .lcout(n2271),
            .ltout(),
            .carryin(\quad_counter1.n19751 ),
            .carryout(\quad_counter1.n19752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_23_lut_LC_12_17_6 .C_ON=1'b1;
    defparam \quad_counter1.add_613_23_lut_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_23_lut_LC_12_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_23_lut_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__40264),
            .in2(N__33136),
            .in3(N__32793),
            .lcout(n2270),
            .ltout(),
            .carryin(\quad_counter1.n19752 ),
            .carryout(\quad_counter1.n19753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_24_lut_LC_12_17_7 .C_ON=1'b1;
    defparam \quad_counter1.add_613_24_lut_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_24_lut_LC_12_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_24_lut_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__33109),
            .in2(N__34659),
            .in3(N__32778),
            .lcout(n2269),
            .ltout(),
            .carryin(\quad_counter1.n19753 ),
            .carryout(\quad_counter1.n19754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_25_lut_LC_12_18_0 .C_ON=1'b1;
    defparam \quad_counter1.add_613_25_lut_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_25_lut_LC_12_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_25_lut_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__38542),
            .in2(N__33137),
            .in3(N__32775),
            .lcout(n2268),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\quad_counter1.n19755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_26_lut_LC_12_18_1 .C_ON=1'b1;
    defparam \quad_counter1.add_613_26_lut_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_26_lut_LC_12_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_26_lut_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__33113),
            .in2(N__37946),
            .in3(N__32772),
            .lcout(n2267),
            .ltout(),
            .carryin(\quad_counter1.n19755 ),
            .carryout(\quad_counter1.n19756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_27_lut_LC_12_18_2 .C_ON=1'b1;
    defparam \quad_counter1.add_613_27_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_27_lut_LC_12_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_27_lut_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__35360),
            .in2(N__33138),
            .in3(N__32754),
            .lcout(n2266),
            .ltout(),
            .carryin(\quad_counter1.n19756 ),
            .carryout(\quad_counter1.n19757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_28_lut_LC_12_18_3 .C_ON=1'b1;
    defparam \quad_counter1.add_613_28_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_28_lut_LC_12_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_28_lut_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__33117),
            .in2(N__38365),
            .in3(N__32751),
            .lcout(n2265),
            .ltout(),
            .carryin(\quad_counter1.n19757 ),
            .carryout(\quad_counter1.n19758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_29_lut_LC_12_18_4 .C_ON=1'b1;
    defparam \quad_counter1.add_613_29_lut_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_29_lut_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_29_lut_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__34884),
            .in2(N__33139),
            .in3(N__32748),
            .lcout(n2264),
            .ltout(),
            .carryin(\quad_counter1.n19758 ),
            .carryout(\quad_counter1.n19759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_30_lut_LC_12_18_5 .C_ON=1'b1;
    defparam \quad_counter1.add_613_30_lut_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_30_lut_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_30_lut_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__33121),
            .in2(N__39972),
            .in3(N__33150),
            .lcout(n2263),
            .ltout(),
            .carryin(\quad_counter1.n19759 ),
            .carryout(\quad_counter1.n19760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_31_lut_LC_12_18_6 .C_ON=1'b1;
    defparam \quad_counter1.add_613_31_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_31_lut_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_31_lut_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__38673),
            .in2(N__33140),
            .in3(N__33147),
            .lcout(n2262),
            .ltout(),
            .carryin(\quad_counter1.n19760 ),
            .carryout(\quad_counter1.n19761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_32_lut_LC_12_18_7 .C_ON=1'b1;
    defparam \quad_counter1.add_613_32_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_32_lut_LC_12_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_613_32_lut_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__33125),
            .in2(N__38811),
            .in3(N__33144),
            .lcout(n2261),
            .ltout(),
            .carryin(\quad_counter1.n19761 ),
            .carryout(\quad_counter1.n19762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_613_33_lut_LC_12_19_0 .C_ON=1'b0;
    defparam \quad_counter1.add_613_33_lut_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_613_33_lut_LC_12_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter1.add_613_33_lut_LC_12_19_0  (
            .in0(N__40331),
            .in1(N__33141),
            .in2(_gnd_net_),
            .in3(N__32934),
            .lcout(n2260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__1__5452_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__1__5452_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__1__5452_LC_12_19_1 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_frame_9__1__5452_LC_12_19_1  (
            .in0(N__38288),
            .in1(N__48249),
            .in2(N__36363),
            .in3(N__45991),
            .lcout(data_out_frame_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21017_4_lut_LC_12_19_2 .C_ON=1'b0;
    defparam \c0.i21017_4_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21017_4_lut_LC_12_19_2 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.i21017_4_lut_LC_12_19_2  (
            .in0(N__41017),
            .in1(N__35409),
            .in2(N__40815),
            .in3(N__33240),
            .lcout(),
            .ltout(\c0.n24784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21250_4_lut_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.i21250_4_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i21250_4_lut_LC_12_19_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.i21250_4_lut_LC_12_19_3  (
            .in0(N__42891),
            .in1(N__40767),
            .in2(N__32931),
            .in3(N__41018),
            .lcout(n25019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__2__5435_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__2__5435_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__2__5435_LC_12_19_4 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_frame_11__2__5435_LC_12_19_4  (
            .in0(N__45989),
            .in1(N__32912),
            .in2(N__32884),
            .in3(N__48248),
            .lcout(data_out_frame_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78611),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i18_LC_12_19_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i18_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i18_LC_12_19_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \quad_counter1.count_i0_i18_LC_12_19_5  (
            .in0(N__32898),
            .in1(N__32877),
            .in2(_gnd_net_),
            .in3(N__40545),
            .lcout(encoder1_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78611),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i16_LC_12_19_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i16_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i16_LC_12_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i16_LC_12_19_6  (
            .in0(N__40544),
            .in1(N__33282),
            .in2(_gnd_net_),
            .in3(N__34074),
            .lcout(encoder1_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__0__5445_LC_12_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__0__5445_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__0__5445_LC_12_19_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__0__5445_LC_12_19_7  (
            .in0(N__48247),
            .in1(N__45990),
            .in2(N__37950),
            .in3(N__33270),
            .lcout(data_out_frame_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14062_2_lut_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.i14062_2_lut_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14062_2_lut_LC_12_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i14062_2_lut_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__43796),
            .in2(_gnd_net_),
            .in3(N__43901),
            .lcout(\c0.data_out_frame_29_7_N_1482_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21016_3_lut_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.i21016_3_lut_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21016_3_lut_LC_12_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i21016_3_lut_LC_12_20_2  (
            .in0(N__43206),
            .in1(N__33326),
            .in2(_gnd_net_),
            .in3(N__33258),
            .lcout(\c0.n24783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__0__5477_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__0__5477_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__0__5477_LC_12_20_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_6__0__5477_LC_12_20_3  (
            .in0(N__45882),
            .in1(N__48255),
            .in2(N__42567),
            .in3(N__33233),
            .lcout(data_out_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78623),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21165_4_lut_LC_12_20_4 .C_ON=1'b0;
    defparam \c0.i21165_4_lut_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i21165_4_lut_LC_12_20_4 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \c0.i21165_4_lut_LC_12_20_4  (
            .in0(N__43516),
            .in1(N__43998),
            .in2(N__33219),
            .in3(N__39495),
            .lcout(\c0.n24888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__0__5429_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__0__5429_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__0__5429_LC_12_20_5 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_12__0__5429_LC_12_20_5  (
            .in0(N__45880),
            .in1(N__48253),
            .in2(N__40179),
            .in3(N__33186),
            .lcout(data_out_frame_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78623),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_12_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i19_LC_12_20_6  (
            .in0(N__50391),
            .in1(N__38718),
            .in2(_gnd_net_),
            .in3(N__43329),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78623),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__1__5428_LC_12_20_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__1__5428_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__1__5428_LC_12_20_7 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_12__1__5428_LC_12_20_7  (
            .in0(N__45881),
            .in1(N__48254),
            .in2(N__40098),
            .in3(N__33164),
            .lcout(data_out_frame_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78623),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__6__5447_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__6__5447_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__6__5447_LC_12_21_0 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_9__6__5447_LC_12_21_0  (
            .in0(N__45873),
            .in1(N__48246),
            .in2(N__42789),
            .in3(N__33414),
            .lcout(data_out_frame_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__6__5471_LC_12_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__6__5471_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__6__5471_LC_12_21_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__6__5471_LC_12_21_1  (
            .in0(N__48243),
            .in1(N__45875),
            .in2(N__39645),
            .in3(N__33399),
            .lcout(data_out_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__4__5521_LC_12_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__4__5521_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__4__5521_LC_12_21_3 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \c0.data_out_frame_0__4__5521_LC_12_21_3  (
            .in0(N__33387),
            .in1(N__43824),
            .in2(N__33362),
            .in3(N__43911),
            .lcout(data_out_frame_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__2__5451_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__2__5451_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__2__5451_LC_12_21_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_9__2__5451_LC_12_21_4  (
            .in0(N__45872),
            .in1(N__48245),
            .in2(N__39861),
            .in3(N__33341),
            .lcout(data_out_frame_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__4__5433_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__4__5433_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__4__5433_LC_12_21_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_11__4__5433_LC_12_21_5  (
            .in0(N__48242),
            .in1(N__45874),
            .in2(N__33810),
            .in3(N__33327),
            .lcout(data_out_frame_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__2__5419_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__2__5419_LC_12_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__2__5419_LC_12_21_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_13__2__5419_LC_12_21_6  (
            .in0(N__45871),
            .in1(N__48244),
            .in2(N__33311),
            .in3(N__46356),
            .lcout(data_out_frame_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1985_LC_12_21_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1985_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1985_LC_12_21_7 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1985_LC_12_21_7  (
            .in0(N__35964),
            .in1(N__33291),
            .in2(N__43431),
            .in3(N__39110),
            .lcout(\c0.n4_adj_4212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1687_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1687_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1687_LC_12_22_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1687_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__43491),
            .in2(_gnd_net_),
            .in3(N__39412),
            .lcout(\c0.n12976 ),
            .ltout(\c0.n12976_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1237_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1237_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1237_LC_12_22_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \c0.i2_4_lut_adj_1237_LC_12_22_1  (
            .in0(N__35982),
            .in1(N__39089),
            .in2(N__33285),
            .in3(N__48443),
            .lcout(\c0.n63_adj_4249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1175_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1175_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1175_LC_12_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1175_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__36213),
            .in2(_gnd_net_),
            .in3(N__47787),
            .lcout(\c0.n21649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1972_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1972_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1972_LC_12_22_3 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1972_LC_12_22_3  (
            .in0(N__43968),
            .in1(N__44086),
            .in2(_gnd_net_),
            .in3(N__44262),
            .lcout(\c0.n58_adj_4706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14178_2_lut_3_lut_4_lut_LC_12_22_4 .C_ON=1'b0;
    defparam \c0.i14178_2_lut_3_lut_4_lut_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14178_2_lut_3_lut_4_lut_LC_12_22_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.i14178_2_lut_3_lut_4_lut_LC_12_22_4  (
            .in0(N__35616),
            .in1(N__43816),
            .in2(N__44142),
            .in3(N__35664),
            .lcout(\c0.data_out_frame_29_7_N_1482_0 ),
            .ltout(\c0.data_out_frame_29_7_N_1482_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1725_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1725_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1725_LC_12_22_5 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1725_LC_12_22_5  (
            .in0(N__33612),
            .in1(N__39088),
            .in2(N__33435),
            .in3(N__33551),
            .lcout(\c0.n13052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_12_22_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i15_LC_12_22_7  (
            .in0(N__44548),
            .in1(N__50453),
            .in2(_gnd_net_),
            .in3(N__38875),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1670_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1670_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1670_LC_12_23_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1670_LC_12_23_0  (
            .in0(N__35614),
            .in1(_gnd_net_),
            .in2(N__43834),
            .in3(N__35662),
            .lcout(\c0.n9706 ),
            .ltout(\c0.n9706_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14180_4_lut_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.i14180_4_lut_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14180_4_lut_LC_12_23_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i14180_4_lut_LC_12_23_1  (
            .in0(N__33432),
            .in1(N__33426),
            .in2(N__33420),
            .in3(N__49043),
            .lcout(\c0.n9248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1545_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1545_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1545_LC_12_23_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1545_LC_12_23_2  (
            .in0(N__35615),
            .in1(N__43698),
            .in2(N__43835),
            .in3(N__35663),
            .lcout(\c0.n9587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1771_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1771_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1771_LC_12_23_3 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1771_LC_12_23_3  (
            .in0(N__49793),
            .in1(N__33620),
            .in2(N__35814),
            .in3(N__38913),
            .lcout(\c0.n6 ),
            .ltout(\c0.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1916_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1916_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1916_LC_12_23_4 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \c0.i1_2_lut_adj_1916_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__33501),
            .in2(N__33417),
            .in3(_gnd_net_),
            .lcout(\c0.n21625 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1868_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1868_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1868_LC_12_23_5 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1868_LC_12_23_5  (
            .in0(N__35756),
            .in1(N__44195),
            .in2(N__35562),
            .in3(N__38914),
            .lcout(\c0.n21579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1772_LC_12_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1772_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1772_LC_12_23_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1772_LC_12_23_6  (
            .in0(N__33621),
            .in1(N__35813),
            .in2(_gnd_net_),
            .in3(N__49794),
            .lcout(\c0.n17682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19210_3_lut_4_lut_LC_12_23_7 .C_ON=1'b0;
    defparam \c0.i19210_3_lut_4_lut_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i19210_3_lut_4_lut_LC_12_23_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i19210_3_lut_4_lut_LC_12_23_7  (
            .in0(N__35975),
            .in1(N__39071),
            .in2(N__33611),
            .in3(N__33544),
            .lcout(\c0.n22907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1474_LC_12_24_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1474_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1474_LC_12_24_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_1474_LC_12_24_0  (
            .in0(N__33524),
            .in1(N__39202),
            .in2(N__39705),
            .in3(N__33499),
            .lcout(\c0.n9_adj_4522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i5_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_12_24_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_12_24_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_12_24_1  (
            .in0(N__33500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48941),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78674),
            .ce(),
            .sr(N__33486));
    defparam \c0.i1_2_lut_adj_1912_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1912_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1912_LC_12_24_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1912_LC_12_24_4  (
            .in0(N__36041),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47788),
            .lcout(\c0.n8_adj_4561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1922_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1922_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1922_LC_12_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1922_LC_12_24_5  (
            .in0(N__47789),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36080),
            .lcout(\c0.n21637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1934_LC_12_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1934_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1934_LC_12_24_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1934_LC_12_24_7  (
            .in0(N__47790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33470),
            .lcout(\c0.n8_adj_4558 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i10_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_12_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_12_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__39206),
            .in2(_gnd_net_),
            .in3(N__48928),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78691),
            .ce(),
            .sr(N__39186));
    defparam \c0.FRAME_MATCHER_state_i6_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_12_26_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_12_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_12_26_7  (
            .in0(_gnd_net_),
            .in1(N__36076),
            .in2(_gnd_net_),
            .in3(N__48969),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78704),
            .ce(),
            .sr(N__33759));
    defparam \c0.i2_3_lut_adj_1387_LC_13_8_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1387_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1387_LC_13_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1387_LC_13_8_1  (
            .in0(N__36976),
            .in1(N__45602),
            .in2(_gnd_net_),
            .in3(N__33717),
            .lcout(),
            .ltout(\c0.n22831_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1325_LC_13_8_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1325_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1325_LC_13_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1325_LC_13_8_2  (
            .in0(N__33747),
            .in1(N__42307),
            .in2(N__33741),
            .in3(N__36688),
            .lcout(\c0.n14_adj_4319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1326_LC_13_8_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1326_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1326_LC_13_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1326_LC_13_8_4  (
            .in0(N__45229),
            .in1(N__39835),
            .in2(N__44762),
            .in3(N__39914),
            .lcout(),
            .ltout(\c0.n13_adj_4320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1327_LC_13_8_5 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1327_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1327_LC_13_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1327_LC_13_8_5  (
            .in0(N__33738),
            .in1(N__42822),
            .in2(N__33729),
            .in3(N__33726),
            .lcout(),
            .ltout(\c0.n28_adj_4322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1331_LC_13_8_6 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1331_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1331_LC_13_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1331_LC_13_8_6  (
            .in0(N__34090),
            .in1(N__40266),
            .in2(N__33720),
            .in3(N__39927),
            .lcout(\c0.n34_adj_4328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_13_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_13_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1751_LC_13_9_0  (
            .in0(N__40324),
            .in1(N__47497),
            .in2(_gnd_net_),
            .in3(N__33715),
            .lcout(\c0.n22656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1359_LC_13_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1359_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1359_LC_13_9_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1359_LC_13_9_1  (
            .in0(N__33716),
            .in1(_gnd_net_),
            .in2(N__47502),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n20318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1309_LC_13_9_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1309_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1309_LC_13_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1309_LC_13_9_2  (
            .in0(N__33686),
            .in1(N__34976),
            .in2(N__33636),
            .in3(N__38810),
            .lcout(\c0.n22466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1392_LC_13_9_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1392_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1392_LC_13_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1392_LC_13_9_3  (
            .in0(N__34977),
            .in1(N__34205),
            .in2(N__34098),
            .in3(N__34029),
            .lcout(\c0.n10_adj_4374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21196_2_lut_LC_13_9_5 .C_ON=1'b0;
    defparam \c0.i21196_2_lut_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21196_2_lut_LC_13_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i21196_2_lut_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__34677),
            .in2(_gnd_net_),
            .in3(N__43182),
            .lcout(\c0.n24901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1253_LC_13_9_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1253_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1253_LC_13_9_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1253_LC_13_9_6  (
            .in0(N__34002),
            .in1(N__33993),
            .in2(N__33954),
            .in3(N__33915),
            .lcout(\c0.n10_adj_4274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i16_LC_13_9_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i16_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i16_LC_13_9_7 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \quad_counter0.count_i0_i16_LC_13_9_7  (
            .in0(N__36753),
            .in1(N__47726),
            .in2(N__36803),
            .in3(_gnd_net_),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78705),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_1758_LC_13_10_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1758_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1758_LC_13_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1758_LC_13_10_0  (
            .in0(N__47312),
            .in1(N__44862),
            .in2(N__33885),
            .in3(N__47028),
            .lcout(\c0.n10_adj_4339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1329_LC_13_10_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1329_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1329_LC_13_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1329_LC_13_10_2  (
            .in0(N__40127),
            .in1(N__33870),
            .in2(N__33771),
            .in3(N__45437),
            .lcout(),
            .ltout(\c0.n30_adj_4326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1333_LC_13_10_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1333_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1333_LC_13_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1333_LC_13_10_3  (
            .in0(N__33853),
            .in1(N__33828),
            .in2(N__33819),
            .in3(N__33816),
            .lcout(\c0.n22408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1310_LC_13_10_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1310_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1310_LC_13_10_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1310_LC_13_10_4  (
            .in0(N__33799),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39623),
            .lcout(\c0.n22788 ),
            .ltout(\c0.n22788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1297_LC_13_10_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1297_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1297_LC_13_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1297_LC_13_10_5  (
            .in0(N__44861),
            .in1(N__39841),
            .in2(N__33762),
            .in3(N__36784),
            .lcout(\c0.n22149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i17_LC_13_10_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i17_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i17_LC_13_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i17_LC_13_10_6  (
            .in0(N__40479),
            .in1(N__34233),
            .in2(_gnd_net_),
            .in3(N__35194),
            .lcout(encoder1_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78692),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i8_LC_13_11_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i8_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i8_LC_13_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i8_LC_13_11_0  (
            .in0(N__40144),
            .in1(N__40565),
            .in2(_gnd_net_),
            .in3(N__34218),
            .lcout(encoder1_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1356_LC_13_11_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1356_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1356_LC_13_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1356_LC_13_11_1  (
            .in0(N__45336),
            .in1(N__34206),
            .in2(N__34191),
            .in3(N__39780),
            .lcout(),
            .ltout(\c0.n14_adj_4338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1358_LC_13_11_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1358_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1358_LC_13_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1358_LC_13_11_2  (
            .in0(N__34170),
            .in1(N__34805),
            .in2(N__34161),
            .in3(N__42351),
            .lcout(\c0.n20455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1295_LC_13_11_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1295_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1295_LC_13_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1295_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__40143),
            .in2(_gnd_net_),
            .in3(N__34109),
            .lcout(\c0.n20461 ),
            .ltout(\c0.n20461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1778_LC_13_11_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1778_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1778_LC_13_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1778_LC_13_11_4  (
            .in0(N__40267),
            .in1(N__44773),
            .in2(N__34158),
            .in3(N__44370),
            .lcout(\c0.n22327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i25_LC_13_11_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i25_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i25_LC_13_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i25_LC_13_11_5  (
            .in0(N__41325),
            .in1(N__37065),
            .in2(_gnd_net_),
            .in3(N__47657),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78675),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i27_LC_13_11_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i27_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i27_LC_13_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i27_LC_13_11_6  (
            .in0(N__47658),
            .in1(N__36993),
            .in2(_gnd_net_),
            .in3(N__45587),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1339_LC_13_12_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1339_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1339_LC_13_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1339_LC_13_12_0  (
            .in0(N__37188),
            .in1(N__34150),
            .in2(N__34614),
            .in3(N__34113),
            .lcout(\c0.n21364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i6_LC_13_12_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i6_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i6_LC_13_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i6_LC_13_12_2  (
            .in0(N__42770),
            .in1(N__36723),
            .in2(_gnd_net_),
            .in3(N__47610),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78659),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1770_LC_13_12_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1770_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1770_LC_13_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1770_LC_13_12_4  (
            .in0(N__41317),
            .in1(N__43415),
            .in2(N__36623),
            .in3(N__42535),
            .lcout(\c0.n22268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1761_LC_13_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1761_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1761_LC_13_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1761_LC_13_12_5  (
            .in0(N__45519),
            .in1(N__46440),
            .in2(N__46361),
            .in3(N__45436),
            .lcout(\c0.n10497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20988_4_lut_LC_13_12_6 .C_ON=1'b0;
    defparam \c0.i20988_4_lut_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20988_4_lut_LC_13_12_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.i20988_4_lut_LC_13_12_6  (
            .in0(N__40835),
            .in1(N__41054),
            .in2(N__34305),
            .in3(N__34287),
            .lcout(\c0.n24755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i24_LC_13_12_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i24_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i24_LC_13_12_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i24_LC_13_12_7  (
            .in0(N__37074),
            .in1(_gnd_net_),
            .in2(N__47652),
            .in3(N__42537),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78659),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1821_LC_13_13_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1821_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1821_LC_13_13_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1821_LC_13_13_0  (
            .in0(N__41365),
            .in1(N__34262),
            .in2(N__44631),
            .in3(N__34448),
            .lcout(),
            .ltout(\c0.n19_adj_4693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1819_LC_13_13_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1819_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1819_LC_13_13_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1819_LC_13_13_1  (
            .in0(N__46179),
            .in1(N__37218),
            .in2(N__34245),
            .in3(N__34239),
            .lcout(),
            .ltout(\c0.n6_adj_4691_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1818_LC_13_13_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1818_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1818_LC_13_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1818_LC_13_13_2  (
            .in0(N__41229),
            .in1(N__41943),
            .in2(N__34242),
            .in3(N__34455),
            .lcout(\c0.n20404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1820_LC_13_13_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1820_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1820_LC_13_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1820_LC_13_13_3  (
            .in0(N__50584),
            .in1(N__41535),
            .in2(N__46448),
            .in3(N__45440),
            .lcout(\c0.n21_adj_4692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1312_LC_13_13_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1312_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1312_LC_13_13_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1312_LC_13_13_4  (
            .in0(N__35033),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40079),
            .lcout(\c0.n22372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1420_LC_13_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1420_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1420_LC_13_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1420_LC_13_13_5  (
            .in0(N__40080),
            .in1(N__35034),
            .in2(_gnd_net_),
            .in3(N__37201),
            .lcout(\c0.n20766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1791_LC_13_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1791_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1791_LC_13_13_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1791_LC_13_13_6  (
            .in0(N__41536),
            .in1(_gnd_net_),
            .in2(N__37170),
            .in3(N__41104),
            .lcout(\c0.n21457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1817_LC_13_13_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1817_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1817_LC_13_13_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1817_LC_13_13_7  (
            .in0(N__41179),
            .in1(N__37164),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n21489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1341_LC_13_14_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1341_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1341_LC_13_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1341_LC_13_14_0  (
            .in0(N__44901),
            .in1(N__34377),
            .in2(N__34432),
            .in3(N__34389),
            .lcout(\c0.n21330 ),
            .ltout(\c0.n21330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1342_LC_13_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1342_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1342_LC_13_14_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1342_LC_13_14_1  (
            .in0(N__41107),
            .in1(_gnd_net_),
            .in2(N__34380),
            .in3(_gnd_net_),
            .lcout(\c0.n20511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1340_LC_13_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1340_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1340_LC_13_14_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1340_LC_13_14_3  (
            .in0(N__37577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45123),
            .lcout(\c0.n6_adj_4331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1990_LC_13_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1990_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1990_LC_13_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1990_LC_13_14_5  (
            .in0(N__41108),
            .in1(N__34371),
            .in2(_gnd_net_),
            .in3(N__37169),
            .lcout(),
            .ltout(\c0.n6_adj_4215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__0__5301_LC_13_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__0__5301_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__0__5301_LC_13_14_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__0__5301_LC_13_14_6  (
            .in0(N__38021),
            .in1(N__34356),
            .in2(N__34323),
            .in3(N__37601),
            .lcout(\c0.data_out_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78636),
            .ce(N__45050),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_13_14_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_13_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_13_14_7  (
            .in0(N__34530),
            .in1(N__34518),
            .in2(_gnd_net_),
            .in3(N__43218),
            .lcout(\c0.n26_adj_4570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_13_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_13_15_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_13_15_0  (
            .in0(N__45439),
            .in1(N__34781),
            .in2(N__45517),
            .in3(N__37258),
            .lcout(\c0.n10529 ),
            .ltout(\c0.n10529_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1293_LC_13_15_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1293_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1293_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1293_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__46789),
            .in2(N__34500),
            .in3(N__46247),
            .lcout(\c0.n21437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_13_15_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_13_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_13_15_2  (
            .in0(N__46790),
            .in1(N__34476),
            .in2(_gnd_net_),
            .in3(N__46752),
            .lcout(\c0.n21393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1285_LC_13_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1285_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1285_LC_13_15_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1285_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__35285),
            .in2(_gnd_net_),
            .in3(N__45438),
            .lcout(\c0.n22489 ),
            .ltout(\c0.n22489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1289_LC_13_15_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1289_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1289_LC_13_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1289_LC_13_15_4  (
            .in0(N__45507),
            .in1(N__41911),
            .in2(N__34497),
            .in3(N__34816),
            .lcout(\c0.n21416 ),
            .ltout(\c0.n21416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_2051_LC_13_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_2051_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_2051_LC_13_15_5 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_2051_LC_13_15_5  (
            .in0(N__46522),
            .in1(N__41912),
            .in2(N__34494),
            .in3(_gnd_net_),
            .lcout(\c0.n22671 ),
            .ltout(\c0.n22671_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_2044_LC_13_15_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_2044_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_2044_LC_13_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_2044_LC_13_15_6  (
            .in0(N__35286),
            .in1(N__34491),
            .in2(N__34479),
            .in3(N__34817),
            .lcout(\c0.n20230 ),
            .ltout(\c0.n20230_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__5__5288_LC_13_15_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__5__5288_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__5__5288_LC_13_15_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__5__5288_LC_13_15_7  (
            .in0(N__46884),
            .in1(N__46791),
            .in2(N__34470),
            .in3(N__45105),
            .lcout(\c0.data_out_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78624),
            .ce(N__45060),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__1__5468_LC_13_16_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__1__5468_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__1__5468_LC_13_16_0 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_7__1__5468_LC_13_16_0  (
            .in0(N__45994),
            .in1(N__48132),
            .in2(N__40227),
            .in3(N__34841),
            .lcout(data_out_frame_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78612),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i21_LC_13_16_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i21_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i21_LC_13_16_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter1.count_i0_i21_LC_13_16_1  (
            .in0(N__34827),
            .in1(_gnd_net_),
            .in2(N__40575),
            .in3(N__40265),
            .lcout(encoder1_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78612),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1291_LC_13_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1291_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1291_LC_13_16_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1291_LC_13_16_2  (
            .in0(N__35287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34821),
            .lcout(\c0.n22722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1823_LC_13_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1823_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1823_LC_13_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1823_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__34776),
            .in2(_gnd_net_),
            .in3(N__46348),
            .lcout(\c0.n22797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__0__5453_LC_13_16_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__0__5453_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__0__5453_LC_13_16_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_9__0__5453_LC_13_16_4  (
            .in0(N__45995),
            .in1(N__48133),
            .in2(N__36432),
            .in3(N__34691),
            .lcout(data_out_frame_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78612),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__4__5481_LC_13_16_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__4__5481_LC_13_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__4__5481_LC_13_16_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__4__5481_LC_13_16_5  (
            .in0(N__48131),
            .in1(N__45996),
            .in2(N__43296),
            .in3(N__34673),
            .lcout(data_out_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78612),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1337_LC_13_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1337_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1337_LC_13_16_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1337_LC_13_16_6  (
            .in0(N__34654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34602),
            .lcout(\c0.n22366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_8_i3_2_lut_LC_13_16_7 .C_ON=1'b0;
    defparam \c0.select_367_Select_8_i3_2_lut_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_8_i3_2_lut_LC_13_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_8_i3_2_lut_LC_13_16_7  (
            .in0(N__52695),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71543),
            .lcout(\c0.n3_adj_4420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__2__5467_LC_13_17_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__2__5467_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__2__5467_LC_13_17_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_frame_7__2__5467_LC_13_17_0  (
            .in0(N__34544),
            .in1(N__46050),
            .in2(N__44871),
            .in3(N__48142),
            .lcout(data_out_frame_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__3__5426_LC_13_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__3__5426_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__3__5426_LC_13_17_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_out_frame_12__3__5426_LC_13_17_1  (
            .in0(N__46047),
            .in1(N__35078),
            .in2(N__48240),
            .in3(N__35133),
            .lcout(data_out_frame_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__2__5427_LC_13_17_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__2__5427_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__2__5427_LC_13_17_2 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_frame_12__2__5427_LC_13_17_2  (
            .in0(N__35060),
            .in1(N__48134),
            .in2(N__35039),
            .in3(N__46051),
            .lcout(data_out_frame_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78597),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i10_LC_13_17_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i10_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i10_LC_13_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i10_LC_13_17_3  (
            .in0(N__40568),
            .in1(N__35046),
            .in2(_gnd_net_),
            .in3(N__35032),
            .lcout(encoder1_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__6__5479_LC_13_17_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__6__5479_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__6__5479_LC_13_17_5 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_out_frame_5__6__5479_LC_13_17_5  (
            .in0(N__46048),
            .in1(N__34991),
            .in2(N__48241),
            .in3(N__43408),
            .lcout(data_out_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__7__5422_LC_13_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__7__5422_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__7__5422_LC_13_17_6 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_frame_12__7__5422_LC_13_17_6  (
            .in0(N__34928),
            .in1(N__46049),
            .in2(N__34975),
            .in3(N__48141),
            .lcout(data_out_frame_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1214_LC_13_17_7 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1214_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1214_LC_13_17_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i10_4_lut_adj_1214_LC_13_17_7  (
            .in0(N__37833),
            .in1(N__41682),
            .in2(N__37827),
            .in3(N__38734),
            .lcout(\c0.n63_adj_4238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i28_LC_13_18_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i28_LC_13_18_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i28_LC_13_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i28_LC_13_18_0  (
            .in0(N__40563),
            .in1(N__34914),
            .in2(_gnd_net_),
            .in3(N__39962),
            .lcout(encoder1_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78613),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i27_LC_13_18_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i27_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i27_LC_13_18_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \quad_counter1.count_i0_i27_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__40562),
            .in2(N__34908),
            .in3(N__34888),
            .lcout(encoder1_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78613),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__3__5482_LC_13_18_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__3__5482_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__3__5482_LC_13_18_2 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_5__3__5482_LC_13_18_2  (
            .in0(N__48239),
            .in1(N__45993),
            .in2(N__46962),
            .in3(N__34856),
            .lcout(data_out_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78613),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i29_LC_13_18_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i29_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i29_LC_13_18_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i29_LC_13_18_3  (
            .in0(N__38674),
            .in1(N__35325),
            .in2(_gnd_net_),
            .in3(N__40564),
            .lcout(encoder1_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78613),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__6__5439_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__6__5439_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__6__5439_LC_13_18_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_10__6__5439_LC_13_18_4  (
            .in0(N__48238),
            .in1(N__45992),
            .in2(N__35318),
            .in3(N__38808),
            .lcout(data_out_frame_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78613),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1209_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1209_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1209_LC_13_18_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i6_4_lut_adj_1209_LC_13_18_5  (
            .in0(N__38612),
            .in1(N__48632),
            .in2(N__44492),
            .in3(N__49242),
            .lcout(\c0.n16_adj_4233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__4__5417_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__4__5417_LC_13_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__4__5417_LC_13_19_0 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_13__4__5417_LC_13_19_0  (
            .in0(N__45983),
            .in1(N__48205),
            .in2(N__35298),
            .in3(N__35418),
            .lcout(data_out_frame_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__0__5461_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__0__5461_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__0__5461_LC_13_19_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__0__5461_LC_13_19_1  (
            .in0(N__48204),
            .in1(N__45988),
            .in2(N__42882),
            .in3(N__35225),
            .lcout(data_out_frame_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__4__5465_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__4__5465_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__4__5465_LC_13_19_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_7__4__5465_LC_13_19_2  (
            .in0(N__45985),
            .in1(N__45348),
            .in2(N__48381),
            .in3(N__35507),
            .lcout(data_out_frame_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__1__5436_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__1__5436_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__1__5436_LC_13_19_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_11__1__5436_LC_13_19_3  (
            .in0(N__48202),
            .in1(N__45986),
            .in2(N__35211),
            .in3(N__38306),
            .lcout(data_out_frame_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1211_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1211_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1211_LC_13_19_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i9_4_lut_adj_1211_LC_13_19_4  (
            .in0(N__39171),
            .in1(N__38568),
            .in2(N__41838),
            .in3(N__35172),
            .lcout(\c0.n63_adj_4235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__7__5430_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__7__5430_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__7__5430_LC_13_19_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_11__7__5430_LC_13_19_5  (
            .in0(N__48203),
            .in1(N__45987),
            .in2(N__38553),
            .in3(N__35162),
            .lcout(data_out_frame_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__5__5416_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__5__5416_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__5__5416_LC_13_19_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_frame_13__5__5416_LC_13_19_6  (
            .in0(N__45984),
            .in1(N__41190),
            .in2(N__48380),
            .in3(N__35147),
            .lcout(data_out_frame_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_13_19_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_13_19_7  (
            .in0(N__35417),
            .in1(N__43160),
            .in2(_gnd_net_),
            .in3(N__41718),
            .lcout(\c0.n11_adj_4669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__4__5457_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__4__5457_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__4__5457_LC_13_20_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_8__4__5457_LC_13_20_0  (
            .in0(N__48207),
            .in1(N__45878),
            .in2(N__36500),
            .in3(N__42905),
            .lcout(data_out_frame_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78637),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_13_20_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i32_LC_13_20_1  (
            .in0(N__76384),
            .in1(N__50482),
            .in2(_gnd_net_),
            .in3(N__38761),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78637),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_13_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i6_LC_13_20_2  (
            .in0(N__50481),
            .in1(N__42436),
            .in2(_gnd_net_),
            .in3(N__38847),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78637),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14067_3_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.i14067_3_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14067_3_lut_LC_13_20_3 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \c0.i14067_3_lut_LC_13_20_3  (
            .in0(N__35637),
            .in1(N__43623),
            .in2(_gnd_net_),
            .in3(N__35603),
            .lcout(data_out_frame_29_7_N_2878_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__5__5456_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__5__5456_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__5__5456_LC_13_20_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_8__5__5456_LC_13_20_4  (
            .in0(N__48208),
            .in1(N__35399),
            .in2(N__42329),
            .in3(N__45879),
            .lcout(data_out_frame_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78637),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__5__5464_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__5__5464_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__5__5464_LC_13_20_5 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_7__5__5464_LC_13_20_5  (
            .in0(N__45876),
            .in1(N__48209),
            .in2(N__45672),
            .in3(N__35381),
            .lcout(data_out_frame_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78637),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__1__5444_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__1__5444_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__1__5444_LC_13_20_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_10__1__5444_LC_13_20_6  (
            .in0(N__48206),
            .in1(N__45877),
            .in2(N__35367),
            .in3(N__38319),
            .lcout(data_out_frame_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78637),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1950_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1950_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1950_LC_13_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1950_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__39704),
            .in2(_gnd_net_),
            .in3(N__47814),
            .lcout(\c0.n8_adj_4555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__4__5473_LC_13_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__4__5473_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__4__5473_LC_13_21_0 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \c0.data_out_frame_6__4__5473_LC_13_21_0  (
            .in0(N__48364),
            .in1(N__35520),
            .in2(N__45997),
            .in3(N__36984),
            .lcout(data_out_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78649),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1688_LC_13_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1688_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1688_LC_13_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1688_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__35602),
            .in2(_gnd_net_),
            .in3(N__35651),
            .lcout(\c0.n7570 ),
            .ltout(\c0.n7570_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1671_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1671_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1671_LC_13_21_2 .LUT_INIT=16'b1011001111111111;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1671_LC_13_21_2  (
            .in0(N__35471),
            .in1(N__43752),
            .in2(N__35523),
            .in3(N__43899),
            .lcout(\c0.n4_adj_4654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_13_21_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_13_21_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_13_21_3  (
            .in0(N__35519),
            .in1(N__43062),
            .in2(_gnd_net_),
            .in3(N__35511),
            .lcout(\c0.n5_adj_4217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1437_LC_13_21_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1437_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1437_LC_13_21_4 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \c0.i1_4_lut_adj_1437_LC_13_21_4  (
            .in0(N__39240),
            .in1(N__43753),
            .in2(N__35430),
            .in3(N__43900),
            .lcout(\c0.n13055 ),
            .ltout(\c0.n13055_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1781_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1781_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1781_LC_13_21_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1781_LC_13_21_5  (
            .in0(N__43967),
            .in1(N__44104),
            .in2(N__35493),
            .in3(N__43515),
            .lcout(n13058),
            .ltout(n13058_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__6__5463_LC_13_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__6__5463_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__6__5463_LC_13_21_6 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.data_out_frame_7__6__5463_LC_13_21_6  (
            .in0(N__48365),
            .in1(N__42267),
            .in2(N__35490),
            .in3(N__35486),
            .lcout(data_out_frame_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78649),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1531_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1531_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1531_LC_13_22_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_1531_LC_13_22_0  (
            .in0(N__44045),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43513),
            .lcout(\c0.n12992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1539_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1539_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1539_LC_13_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1539_LC_13_22_1  (
            .in0(N__35472),
            .in1(N__43611),
            .in2(N__47895),
            .in3(N__35953),
            .lcout(\c0.n5_adj_4477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_13_22_4 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_13_22_4 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_13_22_4  (
            .in0(N__47235),
            .in1(N__47102),
            .in2(N__49638),
            .in3(N__47142),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1905_LC_13_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1905_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1905_LC_13_23_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i1_2_lut_adj_1905_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__43655),
            .in2(_gnd_net_),
            .in3(N__39333),
            .lcout(),
            .ltout(\c0.n14_adj_4727_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1907_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1907_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1907_LC_13_23_1 .LUT_INIT=16'b1100000011101110;
    LogicCell40 \c0.i2_4_lut_adj_1907_LC_13_23_1  (
            .in0(N__48510),
            .in1(N__35721),
            .in2(N__35694),
            .in3(N__35690),
            .lcout(\c0.n6_adj_4728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1894_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1894_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1894_LC_13_23_3 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \c0.i2_4_lut_adj_1894_LC_13_23_3  (
            .in0(N__39334),
            .in1(N__35689),
            .in2(N__48515),
            .in3(N__43865),
            .lcout(\c0.n24386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_13_23_4 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_13_23_4  (
            .in0(N__35604),
            .in1(N__43809),
            .in2(N__43452),
            .in3(N__35652),
            .lcout(\c0.data_out_frame_29_7_N_1482_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1245_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1245_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1245_LC_13_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i4_4_lut_adj_1245_LC_13_23_6  (
            .in0(N__39120),
            .in1(N__47366),
            .in2(N__45998),
            .in3(N__53807),
            .lcout(\c0.n2004 ),
            .ltout(\c0.n2004_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1572_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1572_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1572_LC_13_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1572_LC_13_23_7  (
            .in0(N__35653),
            .in1(N__35605),
            .in2(N__35574),
            .in3(N__43820),
            .lcout(\c0.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20970_4_lut_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.i20970_4_lut_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20970_4_lut_LC_13_24_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i20970_4_lut_LC_13_24_0  (
            .in0(N__44327),
            .in1(N__36009),
            .in2(N__35571),
            .in3(N__39090),
            .lcout(\c0.n24736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1530_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1530_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1530_LC_13_24_1 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1530_LC_13_24_1  (
            .in0(N__39755),
            .in1(_gnd_net_),
            .in2(N__35561),
            .in3(N__36159),
            .lcout(\c0.n28_adj_4565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1658_LC_13_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1658_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1658_LC_13_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1658_LC_13_24_2  (
            .in0(N__44325),
            .in1(N__35554),
            .in2(N__36166),
            .in3(N__39754),
            .lcout(\c0.n16919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1557_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1557_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1557_LC_13_24_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1557_LC_13_24_3  (
            .in0(N__47894),
            .in1(N__43610),
            .in2(_gnd_net_),
            .in3(N__44326),
            .lcout(\c0.n6_adj_4583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1475_LC_13_24_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1475_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1475_LC_13_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_1475_LC_13_24_4  (
            .in0(N__36081),
            .in1(N__36054),
            .in2(N__36042),
            .in3(N__36015),
            .lcout(\c0.n22145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1533_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1533_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1533_LC_13_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1533_LC_13_24_5  (
            .in0(N__36259),
            .in1(N__49036),
            .in2(N__35915),
            .in3(N__35849),
            .lcout(\c0.n20_adj_4265 ),
            .ltout(\c0.n20_adj_4265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1248_LC_13_24_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1248_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1248_LC_13_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_1248_LC_13_24_6  (
            .in0(N__47893),
            .in1(N__35999),
            .in2(N__35985),
            .in3(N__35922),
            .lcout(\c0.n22148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1247_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1247_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1247_LC_13_24_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1247_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__43609),
            .in2(_gnd_net_),
            .in3(N__35943),
            .lcout(\c0.n6_adj_4264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_1963_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1963_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1963_LC_13_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1963_LC_13_25_0  (
            .in0(N__35916),
            .in1(N__36266),
            .in2(N__35871),
            .in3(N__35853),
            .lcout(\c0.n7_adj_4741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2003_LC_13_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2003_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2003_LC_13_25_1 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2003_LC_13_25_1  (
            .in0(N__49829),
            .in1(N__39250),
            .in2(N__53916),
            .in3(N__43836),
            .lcout(\c0.n9683 ),
            .ltout(\c0.n9683_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_13_25_2 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \c0.i1_4_lut_LC_13_25_2  (
            .in0(N__35799),
            .in1(N__48475),
            .in2(N__35790),
            .in3(N__44276),
            .lcout(\c0.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1981_LC_13_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1981_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1981_LC_13_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1981_LC_13_25_3  (
            .in0(N__47817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49073),
            .lcout(\c0.n21643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2008_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2008_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2008_LC_13_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_2008_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(N__36267),
            .in2(_gnd_net_),
            .in3(N__47818),
            .lcout(\c0.n21653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1971_LC_13_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1971_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1971_LC_13_25_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1971_LC_13_25_6  (
            .in0(N__39744),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47815),
            .lcout(\c0.n21639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1976_LC_13_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1976_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1976_LC_13_25_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.i1_2_lut_adj_1976_LC_13_25_7  (
            .in0(N__47816),
            .in1(_gnd_net_),
            .in2(N__49139),
            .in3(_gnd_net_),
            .lcout(\c0.n21641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i29_LC_13_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_13_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_13_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__36205),
            .in2(_gnd_net_),
            .in3(N__48985),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78716),
            .ce(),
            .sr(N__36183));
    defparam \c0.FRAME_MATCHER_state_i24_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_13_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_13_27_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_13_27_0  (
            .in0(N__48987),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36155),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78728),
            .ce(),
            .sr(N__36126));
    defparam \c0.FRAME_MATCHER_state_i21_LC_13_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_13_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_13_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_13_28_0  (
            .in0(_gnd_net_),
            .in1(N__49069),
            .in2(_gnd_net_),
            .in3(N__48989),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78741),
            .ce(),
            .sr(N__36111));
    defparam \quad_counter0.count_i0_i2_LC_14_8_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i2_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i2_LC_14_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i2_LC_14_8_0  (
            .in0(N__47728),
            .in1(N__36300),
            .in2(_gnd_net_),
            .in3(N__39840),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78730),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i3_LC_14_8_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i3_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i3_LC_14_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i3_LC_14_8_1  (
            .in0(N__44755),
            .in1(N__36291),
            .in2(_gnd_net_),
            .in3(N__47730),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78730),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i7_LC_14_8_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i7_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i7_LC_14_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i7_LC_14_8_3  (
            .in0(N__36689),
            .in1(N__36645),
            .in2(_gnd_net_),
            .in3(N__47731),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78730),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i30_LC_14_8_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i30_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i30_LC_14_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i30_LC_14_8_5  (
            .in0(N__39612),
            .in1(N__36825),
            .in2(_gnd_net_),
            .in3(N__47729),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78730),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i0_LC_14_8_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i0_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i0_LC_14_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i0_LC_14_8_6  (
            .in0(N__47727),
            .in1(N__36372),
            .in2(_gnd_net_),
            .in3(N__36414),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78730),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_1_LC_14_9_0 .C_ON=1'b1;
    defparam \quad_counter0.add_647_1_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_1_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter0.add_647_1_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__37384),
            .in2(N__37447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\quad_counter0.n19763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_2_lut_LC_14_9_1 .C_ON=1'b1;
    defparam \quad_counter0.add_647_2_lut_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_2_lut_LC_14_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_2_lut_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__36413),
            .in2(N__36387),
            .in3(N__36366),
            .lcout(n2357),
            .ltout(),
            .carryin(\quad_counter0.n19763 ),
            .carryout(\quad_counter0.n19764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_3_lut_LC_14_9_2 .C_ON=1'b1;
    defparam \quad_counter0.add_647_3_lut_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_3_lut_LC_14_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_3_lut_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__36356),
            .in2(N__37448),
            .in3(N__36303),
            .lcout(n2356),
            .ltout(),
            .carryin(\quad_counter0.n19764 ),
            .carryout(\quad_counter0.n19765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_4_lut_LC_14_9_3 .C_ON=1'b1;
    defparam \quad_counter0.add_647_4_lut_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_4_lut_LC_14_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_4_lut_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__39836),
            .in2(N__37444),
            .in3(N__36294),
            .lcout(n2355),
            .ltout(),
            .carryin(\quad_counter0.n19765 ),
            .carryout(\quad_counter0.n19766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_5_lut_LC_14_9_4 .C_ON=1'b1;
    defparam \quad_counter0.add_647_5_lut_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_5_lut_LC_14_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_5_lut_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__44774),
            .in2(N__37449),
            .in3(N__36285),
            .lcout(n2354),
            .ltout(),
            .carryin(\quad_counter0.n19766 ),
            .carryout(\quad_counter0.n19767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_6_lut_LC_14_9_5 .C_ON=1'b1;
    defparam \quad_counter0.add_647_6_lut_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_6_lut_LC_14_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_6_lut_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__45263),
            .in2(N__37445),
            .in3(N__36270),
            .lcout(n2353),
            .ltout(),
            .carryin(\quad_counter0.n19767 ),
            .carryout(\quad_counter0.n19768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_7_lut_LC_14_9_6 .C_ON=1'b1;
    defparam \quad_counter0.add_647_7_lut_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_7_lut_LC_14_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_7_lut_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__45380),
            .in2(N__37450),
            .in3(N__36726),
            .lcout(n2352),
            .ltout(),
            .carryin(\quad_counter0.n19768 ),
            .carryout(\quad_counter0.n19769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_8_lut_LC_14_9_7 .C_ON=1'b1;
    defparam \quad_counter0.add_647_8_lut_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_8_lut_LC_14_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_8_lut_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__42771),
            .in2(N__37446),
            .in3(N__36714),
            .lcout(n2351),
            .ltout(),
            .carryin(\quad_counter0.n19769 ),
            .carryout(\quad_counter0.n19770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_9_lut_LC_14_10_0 .C_ON=1'b1;
    defparam \quad_counter0.add_647_9_lut_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_9_lut_LC_14_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_9_lut_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__36693),
            .in2(N__37484),
            .in3(N__36636),
            .lcout(n2350),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\quad_counter0.n19771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_10_lut_LC_14_10_1 .C_ON=1'b1;
    defparam \quad_counter0.add_647_10_lut_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_10_lut_LC_14_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_10_lut_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__37454),
            .in2(N__42881),
            .in3(N__36633),
            .lcout(n2349),
            .ltout(),
            .carryin(\quad_counter0.n19771 ),
            .carryout(\quad_counter0.n19772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_11_lut_LC_14_10_2 .C_ON=1'b1;
    defparam \quad_counter0.add_647_11_lut_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_11_lut_LC_14_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_11_lut_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__42656),
            .in2(N__37485),
            .in3(N__36630),
            .lcout(n2348),
            .ltout(),
            .carryin(\quad_counter0.n19772 ),
            .carryout(\quad_counter0.n19773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_12_lut_LC_14_10_3 .C_ON=1'b1;
    defparam \quad_counter0.add_647_12_lut_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_12_lut_LC_14_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_12_lut_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__37458),
            .in2(N__36627),
            .in3(N__36567),
            .lcout(n2347),
            .ltout(),
            .carryin(\quad_counter0.n19773 ),
            .carryout(\quad_counter0.n19774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_13_lut_LC_14_10_4 .C_ON=1'b1;
    defparam \quad_counter0.add_647_13_lut_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_13_lut_LC_14_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_13_lut_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(N__36554),
            .in2(N__37486),
            .in3(N__36507),
            .lcout(n2346),
            .ltout(),
            .carryin(\quad_counter0.n19774 ),
            .carryout(\quad_counter0.n19775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_14_lut_LC_14_10_5 .C_ON=1'b1;
    defparam \quad_counter0.add_647_14_lut_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_14_lut_LC_14_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_14_lut_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__37462),
            .in2(N__36504),
            .in3(N__36435),
            .lcout(n2345),
            .ltout(),
            .carryin(\quad_counter0.n19775 ),
            .carryout(\quad_counter0.n19776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_15_lut_LC_14_10_6 .C_ON=1'b1;
    defparam \quad_counter0.add_647_15_lut_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_15_lut_LC_14_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_15_lut_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__42328),
            .in2(N__37487),
            .in3(N__36813),
            .lcout(n2344),
            .ltout(),
            .carryin(\quad_counter0.n19776 ),
            .carryout(\quad_counter0.n19777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_16_lut_LC_14_10_7 .C_ON=1'b1;
    defparam \quad_counter0.add_647_16_lut_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_16_lut_LC_14_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_16_lut_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__37466),
            .in2(N__47501),
            .in3(N__36810),
            .lcout(n2343),
            .ltout(),
            .carryin(\quad_counter0.n19777 ),
            .carryout(\quad_counter0.n19778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_17_lut_LC_14_11_0 .C_ON=1'b1;
    defparam \quad_counter0.add_647_17_lut_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_17_lut_LC_14_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_17_lut_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__39554),
            .in2(N__37488),
            .in3(N__36807),
            .lcout(n2342),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\quad_counter0.n19779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_18_lut_LC_14_11_1 .C_ON=1'b1;
    defparam \quad_counter0.add_647_18_lut_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_18_lut_LC_14_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_18_lut_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__37470),
            .in2(N__36804),
            .in3(N__36744),
            .lcout(n2341),
            .ltout(),
            .carryin(\quad_counter0.n19779 ),
            .carryout(\quad_counter0.n19780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_19_lut_LC_14_11_2 .C_ON=1'b1;
    defparam \quad_counter0.add_647_19_lut_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_19_lut_LC_14_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_19_lut_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__40213),
            .in2(N__37489),
            .in3(N__36741),
            .lcout(n2340),
            .ltout(),
            .carryin(\quad_counter0.n19780 ),
            .carryout(\quad_counter0.n19781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_20_lut_LC_14_11_3 .C_ON=1'b1;
    defparam \quad_counter0.add_647_20_lut_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_20_lut_LC_14_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_20_lut_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__37474),
            .in2(N__44863),
            .in3(N__36738),
            .lcout(n2339),
            .ltout(),
            .carryin(\quad_counter0.n19781 ),
            .carryout(\quad_counter0.n19782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_21_lut_LC_14_11_4 .C_ON=1'b1;
    defparam \quad_counter0.add_647_21_lut_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_21_lut_LC_14_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_21_lut_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__42401),
            .in2(N__37490),
            .in3(N__36735),
            .lcout(n2338),
            .ltout(),
            .carryin(\quad_counter0.n19782 ),
            .carryout(\quad_counter0.n19783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_22_lut_LC_14_11_5 .C_ON=1'b1;
    defparam \quad_counter0.add_647_22_lut_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_22_lut_LC_14_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_22_lut_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__37478),
            .in2(N__45344),
            .in3(N__36732),
            .lcout(n2337),
            .ltout(),
            .carryin(\quad_counter0.n19783 ),
            .carryout(\quad_counter0.n19784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_23_lut_LC_14_11_6 .C_ON=1'b1;
    defparam \quad_counter0.add_647_23_lut_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_23_lut_LC_14_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_23_lut_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__37479),
            .in2(N__45656),
            .in3(N__36729),
            .lcout(n2336),
            .ltout(),
            .carryin(\quad_counter0.n19784 ),
            .carryout(\quad_counter0.n19785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_24_lut_LC_14_11_7 .C_ON=1'b1;
    defparam \quad_counter0.add_647_24_lut_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_24_lut_LC_14_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_24_lut_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__42257),
            .in2(N__37491),
            .in3(N__37080),
            .lcout(n2335),
            .ltout(),
            .carryin(\quad_counter0.n19785 ),
            .carryout(\quad_counter0.n19786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_25_lut_LC_14_12_0 .C_ON=1'b1;
    defparam \quad_counter0.add_647_25_lut_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_25_lut_LC_14_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_25_lut_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__37337),
            .in2(N__42716),
            .in3(N__37077),
            .lcout(n2334),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\quad_counter0.n19787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_26_lut_LC_14_12_1 .C_ON=1'b1;
    defparam \quad_counter0.add_647_26_lut_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_26_lut_LC_14_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_26_lut_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__42536),
            .in2(N__37380),
            .in3(N__37068),
            .lcout(n2333),
            .ltout(),
            .carryin(\quad_counter0.n19787 ),
            .carryout(\quad_counter0.n19788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_27_lut_LC_14_12_2 .C_ON=1'b1;
    defparam \quad_counter0.add_647_27_lut_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_27_lut_LC_14_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_27_lut_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__37341),
            .in2(N__41327),
            .in3(N__37059),
            .lcout(n2332),
            .ltout(),
            .carryin(\quad_counter0.n19788 ),
            .carryout(\quad_counter0.n19789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_28_lut_LC_14_12_3 .C_ON=1'b1;
    defparam \quad_counter0.add_647_28_lut_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_28_lut_LC_14_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_28_lut_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__37052),
            .in2(N__37381),
            .in3(N__36996),
            .lcout(n2331),
            .ltout(),
            .carryin(\quad_counter0.n19789 ),
            .carryout(\quad_counter0.n19790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_29_lut_LC_14_12_4 .C_ON=1'b1;
    defparam \quad_counter0.add_647_29_lut_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_29_lut_LC_14_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_29_lut_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__37345),
            .in2(N__45614),
            .in3(N__36987),
            .lcout(n2330),
            .ltout(),
            .carryin(\quad_counter0.n19790 ),
            .carryout(\quad_counter0.n19791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_30_lut_LC_14_12_5 .C_ON=1'b1;
    defparam \quad_counter0.add_647_30_lut_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_30_lut_LC_14_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_30_lut_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__36977),
            .in2(N__37382),
            .in3(N__36900),
            .lcout(n2329),
            .ltout(),
            .carryin(\quad_counter0.n19791 ),
            .carryout(\quad_counter0.n19792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_31_lut_LC_14_12_6 .C_ON=1'b1;
    defparam \quad_counter0.add_647_31_lut_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_31_lut_LC_14_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_31_lut_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__37349),
            .in2(N__36893),
            .in3(N__36828),
            .lcout(n2328),
            .ltout(),
            .carryin(\quad_counter0.n19792 ),
            .carryout(\quad_counter0.n19793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_32_lut_LC_14_12_7 .C_ON=1'b1;
    defparam \quad_counter0.add_647_32_lut_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_32_lut_LC_14_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_647_32_lut_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__39624),
            .in2(N__37383),
            .in3(N__36816),
            .lcout(n2327),
            .ltout(),
            .carryin(\quad_counter0.n19793 ),
            .carryout(\quad_counter0.n19794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_647_33_lut_LC_14_13_0 .C_ON=1'b0;
    defparam \quad_counter0.add_647_33_lut_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_647_33_lut_LC_14_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.add_647_33_lut_LC_14_13_0  (
            .in0(N__44684),
            .in1(N__37483),
            .in2(_gnd_net_),
            .in3(N__37293),
            .lcout(),
            .ltout(n2326_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i31_LC_14_13_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i31_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i31_LC_14_13_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter0.count_i0_i31_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__44685),
            .in2(N__37290),
            .in3(N__47696),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1364_LC_14_13_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1364_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1364_LC_14_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1364_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__44683),
            .in2(_gnd_net_),
            .in3(N__45174),
            .lcout(\c0.n10427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1822_LC_14_13_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1822_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1822_LC_14_13_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1822_LC_14_13_3  (
            .in0(N__37637),
            .in1(N__37283),
            .in2(N__37266),
            .in3(N__37227),
            .lcout(\c0.n20_adj_4694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1782_LC_14_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1782_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1782_LC_14_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1782_LC_14_13_5  (
            .in0(N__37208),
            .in1(N__50528),
            .in2(N__40022),
            .in3(N__41102),
            .lcout(\c0.n21355 ),
            .ltout(\c0.n21355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1790_LC_14_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1790_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1790_LC_14_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1790_LC_14_13_6  (
            .in0(N__41103),
            .in1(N__37168),
            .in2(N__37146),
            .in3(N__41537),
            .lcout(\c0.n21327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_1799_LC_14_13_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_1799_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_1799_LC_14_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_1799_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__37143),
            .in2(_gnd_net_),
            .in3(N__37092),
            .lcout(\c0.n15_adj_4686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1219_LC_14_14_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1219_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1219_LC_14_14_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i7_4_lut_adj_1219_LC_14_14_0  (
            .in0(N__38493),
            .in1(N__41820),
            .in2(N__44485),
            .in3(N__48606),
            .lcout(\c0.n13046 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_14_14_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_14_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_0___i18_LC_14_14_1  (
            .in0(N__41821),
            .in1(_gnd_net_),
            .in2(N__49314),
            .in3(N__50438),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1784_LC_14_14_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1784_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1784_LC_14_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1784_LC_14_14_2  (
            .in0(N__37638),
            .in1(N__46610),
            .in2(N__46873),
            .in3(N__37597),
            .lcout(\c0.n24028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1792_LC_14_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1792_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1792_LC_14_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1792_LC_14_14_3  (
            .in0(N__41106),
            .in1(N__46854),
            .in2(_gnd_net_),
            .in3(N__50526),
            .lcout(\c0.n13268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i22_LC_14_14_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i22_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i22_LC_14_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i22_LC_14_14_4  (
            .in0(N__47711),
            .in1(N__37626),
            .in2(_gnd_net_),
            .in3(N__42247),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1301_LC_14_14_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1301_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1301_LC_14_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1301_LC_14_14_5  (
            .in0(N__44433),
            .in1(N__45261),
            .in2(N__37617),
            .in3(N__37556),
            .lcout(\c0.n21360 ),
            .ltout(\c0.n21360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1296_LC_14_14_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1296_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1296_LC_14_14_6 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \c0.i1_2_lut_adj_1296_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__41105),
            .in2(N__37608),
            .in3(_gnd_net_),
            .lcout(\c0.n10504 ),
            .ltout(\c0.n10504_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1299_LC_14_14_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1299_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1299_LC_14_14_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1299_LC_14_14_7  (
            .in0(N__37581),
            .in1(N__44699),
            .in2(N__37560),
            .in3(N__37557),
            .lcout(\c0.n12_adj_4312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1880_LC_14_15_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1880_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1880_LC_14_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1880_LC_14_15_0  (
            .in0(N__37545),
            .in1(N__41589),
            .in2(N__41189),
            .in3(N__46671),
            .lcout(),
            .ltout(\c0.n25_adj_4695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__1__5292_LC_14_15_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__1__5292_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__1__5292_LC_14_15_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__1__5292_LC_14_15_1  (
            .in0(N__37521),
            .in1(N__37671),
            .in2(N__37509),
            .in3(N__37752),
            .lcout(\c0.data_out_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78638),
            .ce(N__45059),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1884_LC_14_15_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1884_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1884_LC_14_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1884_LC_14_15_2  (
            .in0(N__37785),
            .in1(N__37778),
            .in2(N__37761),
            .in3(N__41448),
            .lcout(\c0.n26_adj_4697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__1__5300_LC_14_15_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__1__5300_LC_14_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__1__5300_LC_14_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_frame_28__1__5300_LC_14_15_4  (
            .in0(N__37743),
            .in1(N__37725),
            .in2(_gnd_net_),
            .in3(N__37710),
            .lcout(\c0.data_out_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78638),
            .ce(N__45059),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1834_LC_14_15_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1834_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1834_LC_14_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1834_LC_14_15_5  (
            .in0(N__38006),
            .in1(N__41067),
            .in2(N__37683),
            .in3(N__46155),
            .lcout(\c0.n27_adj_4696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_14_16_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_14_16_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i8_LC_14_16_0  (
            .in0(N__48628),
            .in1(N__50429),
            .in2(_gnd_net_),
            .in3(N__38988),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78626),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_14_16_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_14_16_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i5_LC_14_16_2  (
            .in0(N__37652),
            .in1(N__50428),
            .in2(_gnd_net_),
            .in3(N__37826),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78626),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_14_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_14_16_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i1_LC_14_16_3  (
            .in0(N__42063),
            .in1(_gnd_net_),
            .in2(N__50465),
            .in3(N__37665),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78626),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1215_LC_14_16_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1215_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1215_LC_14_16_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i4_4_lut_adj_1215_LC_14_16_4  (
            .in0(N__43363),
            .in1(N__37664),
            .in2(N__37653),
            .in3(N__38987),
            .lcout(\c0.n10_adj_4239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1221_LC_14_16_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1221_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1221_LC_14_16_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i6_4_lut_adj_1221_LC_14_16_5  (
            .in0(N__37860),
            .in1(N__44525),
            .in2(N__42066),
            .in3(N__37878),
            .lcout(),
            .ltout(\c0.n15_adj_4242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1222_LC_14_16_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1222_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1222_LC_14_16_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i8_4_lut_adj_1222_LC_14_16_6  (
            .in0(N__41698),
            .in1(N__38736),
            .in2(N__37641),
            .in3(N__37791),
            .lcout(\c0.n12898 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1806_LC_14_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1806_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1806_LC_14_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1806_LC_14_16_7  (
            .in0(N__38258),
            .in1(N__38175),
            .in2(_gnd_net_),
            .in3(N__38082),
            .lcout(\c0.n21464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i24_LC_14_17_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i24_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i24_LC_14_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i24_LC_14_17_0  (
            .in0(N__37962),
            .in1(N__40573),
            .in2(_gnd_net_),
            .in3(N__37926),
            .lcout(encoder1_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_14_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_14_17_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i21_LC_14_17_1  (
            .in0(N__37865),
            .in1(N__50426),
            .in2(_gnd_net_),
            .in3(N__42092),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i174_LC_14_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i174_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i174_LC_14_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i174_LC_14_17_2  (
            .in0(N__75909),
            .in1(N__79786),
            .in2(_gnd_net_),
            .in3(N__67648),
            .lcout(data_in_frame_21_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1384_LC_14_17_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1384_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1384_LC_14_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1384_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__47014),
            .in2(_gnd_net_),
            .in3(N__42341),
            .lcout(\c0.n10_adj_4367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1216_LC_14_17_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1216_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1216_LC_14_17_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i5_3_lut_adj_1216_LC_14_17_4  (
            .in0(N__42091),
            .in1(N__39009),
            .in2(_gnd_net_),
            .in3(N__37884),
            .lcout(\c0.n13049 ),
            .ltout(\c0.n13049_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1212_LC_14_17_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1212_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1212_LC_14_17_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i7_4_lut_adj_1212_LC_14_17_5  (
            .in0(N__42438),
            .in1(N__37861),
            .in2(N__37839),
            .in3(N__38630),
            .lcout(),
            .ltout(\c0.n18_adj_4236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1213_LC_14_17_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1213_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1213_LC_14_17_6 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i9_4_lut_adj_1213_LC_14_17_6  (
            .in0(N__44526),
            .in1(N__49424),
            .in2(N__37836),
            .in3(N__38585),
            .lcout(\c0.n20_adj_4237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1220_LC_14_17_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1220_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1220_LC_14_17_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.i5_3_lut_adj_1220_LC_14_17_7  (
            .in0(N__42437),
            .in1(N__37822),
            .in2(_gnd_net_),
            .in3(N__49423),
            .lcout(\c0.n14_adj_4241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1210_LC_14_18_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1210_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1210_LC_14_18_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.i7_4_lut_adj_1210_LC_14_18_0  (
            .in0(N__46919),
            .in1(N__49310),
            .in2(N__38586),
            .in3(N__48679),
            .lcout(\c0.n17_adj_4234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i23_LC_14_18_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i23_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i23_LC_14_18_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i23_LC_14_18_1  (
            .in0(N__38562),
            .in1(N__40558),
            .in2(_gnd_net_),
            .in3(N__38535),
            .lcout(encoder1_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78627),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i13_LC_14_18_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i13_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i13_LC_14_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i13_LC_14_18_2  (
            .in0(N__47732),
            .in1(N__38508),
            .in2(_gnd_net_),
            .in3(N__42297),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78627),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1217_LC_14_18_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1217_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1217_LC_14_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_adj_1217_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__39170),
            .in2(_gnd_net_),
            .in3(N__46918),
            .lcout(\c0.n10_adj_4240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_14_18_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_14_18_4  (
            .in0(N__38393),
            .in1(N__38482),
            .in2(_gnd_net_),
            .in3(N__38415),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78627),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i26_LC_14_19_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i26_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i26_LC_14_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i26_LC_14_19_0  (
            .in0(N__40569),
            .in1(N__38379),
            .in2(_gnd_net_),
            .in3(N__38343),
            .lcout(encoder1_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78639),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_14_19_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_LC_14_19_1  (
            .in0(N__38318),
            .in1(N__40821),
            .in2(N__38307),
            .in3(N__43221),
            .lcout(),
            .ltout(\c0.n25116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n25116_bdd_4_lut_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.n25116_bdd_4_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.n25116_bdd_4_lut_LC_14_19_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n25116_bdd_4_lut_LC_14_19_2  (
            .in0(N__40822),
            .in1(N__38693),
            .in2(N__38292),
            .in3(N__38289),
            .lcout(\c0.n25119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1168_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1168_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1168_LC_14_19_3 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.rx.i1_2_lut_adj_1168_LC_14_19_3  (
            .in0(N__47227),
            .in1(N__46656),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n12981),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_14_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_14_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i11_LC_14_19_4  (
            .in0(N__50472),
            .in1(N__38735),
            .in2(_gnd_net_),
            .in3(N__49264),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78639),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__1__5460_LC_14_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__1__5460_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__1__5460_LC_14_19_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_8__1__5460_LC_14_19_5  (
            .in0(N__48200),
            .in1(N__46011),
            .in2(N__38697),
            .in3(N__42663),
            .lcout(data_out_frame_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78639),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__5__5440_LC_14_19_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__5__5440_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__5__5440_LC_14_19_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_10__5__5440_LC_14_19_6  (
            .in0(N__46010),
            .in1(N__48201),
            .in2(N__38649),
            .in3(N__38675),
            .lcout(data_out_frame_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78639),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1690_LC_14_20_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1690_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1690_LC_14_20_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i8_4_lut_adj_1690_LC_14_20_0  (
            .in0(N__38846),
            .in1(N__38631),
            .in2(N__42122),
            .in3(N__38616),
            .lcout(),
            .ltout(\c0.n20_adj_4308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1290_LC_14_20_1 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1290_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1290_LC_14_20_1 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \c0.i11_3_lut_adj_1290_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__38595),
            .in2(N__38598),
            .in3(N__38886),
            .lcout(n63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1691_LC_14_20_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1691_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1691_LC_14_20_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i7_4_lut_adj_1691_LC_14_20_2  (
            .in0(N__44558),
            .in1(N__42466),
            .in2(N__38762),
            .in3(N__38879),
            .lcout(\c0.n19_adj_4307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1206_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1206_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1206_LC_14_20_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i6_4_lut_adj_1206_LC_14_20_3  (
            .in0(N__42200),
            .in1(N__44557),
            .in2(N__42470),
            .in3(N__49260),
            .lcout(),
            .ltout(\c0.n16_adj_4231_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1208_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1208_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1208_LC_14_20_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i9_4_lut_adj_1208_LC_14_20_4  (
            .in0(N__38754),
            .in1(N__42114),
            .in2(N__38589),
            .in3(N__38829),
            .lcout(\c0.n12986 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20978_4_lut_LC_14_20_6 .C_ON=1'b0;
    defparam \c0.i20978_4_lut_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20978_4_lut_LC_14_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i20978_4_lut_LC_14_20_6  (
            .in0(N__43318),
            .in1(N__42201),
            .in2(N__49268),
            .in3(N__43346),
            .lcout(\c0.n24745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1207_LC_14_21_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1207_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1207_LC_14_21_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i7_4_lut_adj_1207_LC_14_21_0  (
            .in0(N__43345),
            .in1(N__43317),
            .in2(N__38880),
            .in3(N__38845),
            .lcout(\c0.n17_adj_4232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i192_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i192_LC_14_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i192_LC_14_21_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_in_frame_0__i192_LC_14_21_4  (
            .in0(N__80988),
            .in1(N__63965),
            .in2(N__76382),
            .in3(N__80429),
            .lcout(\c0.data_in_frame_23_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78662),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i30_LC_14_21_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i30_LC_14_21_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i30_LC_14_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i30_LC_14_21_6  (
            .in0(N__38823),
            .in1(N__40574),
            .in2(_gnd_net_),
            .in3(N__38787),
            .lcout(encoder1_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_14_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_14_21_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1742_LC_14_21_7  (
            .in0(N__44141),
            .in1(N__39109),
            .in2(_gnd_net_),
            .in3(N__44103),
            .lcout(\c0.n13001 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i88_LC_14_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i88_LC_14_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i88_LC_14_22_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i88_LC_14_22_0  (
            .in0(N__61719),
            .in1(N__73707),
            .in2(N__76383),
            .in3(N__69236),
            .lcout(\c0.data_in_frame_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_14_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_14_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_14_22_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i24_LC_14_22_1  (
            .in0(N__38763),
            .in1(N__50462),
            .in2(_gnd_net_),
            .in3(N__39007),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i213_LC_14_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i213_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i213_LC_14_22_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i213_LC_14_22_2  (
            .in0(N__79442),
            .in1(N__69237),
            .in2(N__77332),
            .in3(N__71887),
            .lcout(\c0.data_in_frame_26_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i212_LC_14_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i212_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i212_LC_14_22_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i212_LC_14_22_3  (
            .in0(N__69235),
            .in1(N__68349),
            .in2(N__76916),
            .in3(N__79443),
            .lcout(\c0.data_in_frame_26_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_14_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_14_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_14_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i30_LC_14_22_4  (
            .in0(N__50460),
            .in1(N__79648),
            .in2(_gnd_net_),
            .in3(N__39168),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_14_22_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i22_LC_14_22_5  (
            .in0(N__39169),
            .in1(N__50461),
            .in2(_gnd_net_),
            .in3(N__42462),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_14_22_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_14_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_14_22_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_14_22_6  (
            .in0(N__47429),
            .in1(N__76883),
            .in2(N__50908),
            .in3(N__50726),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i237_LC_14_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i237_LC_14_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i237_LC_14_22_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i237_LC_14_22_7  (
            .in0(N__56481),
            .in1(N__52013),
            .in2(N__71938),
            .in3(N__75397),
            .lcout(\c0.data_in_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_2046_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_2046_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_2046_LC_14_23_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_2046_LC_14_23_0  (
            .in0(N__43493),
            .in1(N__39370),
            .in2(N__44011),
            .in3(N__39421),
            .lcout(\c0.n13063 ),
            .ltout(\c0.n13063_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_2047_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_2047_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_2047_LC_14_23_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_2047_LC_14_23_1  (
            .in0(N__39422),
            .in1(N__39371),
            .in2(N__39123),
            .in3(N__39020),
            .lcout(\c0.n6_adj_4263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1979_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1979_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1979_LC_14_23_3 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.i3_4_lut_adj_1979_LC_14_23_3  (
            .in0(N__39108),
            .in1(N__38967),
            .in2(N__44331),
            .in3(N__39336),
            .lcout(\c0.n8_adj_4553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1265_2_lut_3_lut_LC_14_23_5 .C_ON=1'b0;
    defparam \c0.i1265_2_lut_3_lut_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1265_2_lut_3_lut_LC_14_23_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i1265_2_lut_3_lut_LC_14_23_5  (
            .in0(N__44131),
            .in1(N__39097),
            .in2(_gnd_net_),
            .in3(N__43492),
            .lcout(\c0.n3325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_14_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_14_23_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i16_LC_14_23_6  (
            .in0(N__50463),
            .in1(N__39008),
            .in2(_gnd_net_),
            .in3(N__38981),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1961_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1961_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1961_LC_14_23_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i1_3_lut_adj_1961_LC_14_23_7  (
            .in0(N__43605),
            .in1(N__38966),
            .in2(_gnd_net_),
            .in3(N__38933),
            .lcout(\c0.n21659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1779_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1779_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1779_LC_14_24_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1779_LC_14_24_0  (
            .in0(N__44002),
            .in1(N__44058),
            .in2(N__48519),
            .in3(N__44108),
            .lcout(\c0.n24422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_2041_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_2041_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_2041_LC_14_24_1 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_2041_LC_14_24_1  (
            .in0(N__39465),
            .in1(N__39423),
            .in2(N__39399),
            .in3(N__39375),
            .lcout(),
            .ltout(\c0.n24596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1287_LC_14_24_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1287_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1287_LC_14_24_2 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \c0.i1_4_lut_adj_1287_LC_14_24_2  (
            .in0(N__39348),
            .in1(N__43514),
            .in2(N__39339),
            .in3(N__39335),
            .lcout(\c0.n4_adj_4306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4626_2_lut_LC_14_24_3 .C_ON=1'b0;
    defparam \c0.i4626_2_lut_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4626_2_lut_LC_14_24_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i4626_2_lut_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__48270),
            .in2(_gnd_net_),
            .in3(N__45889),
            .lcout(\c0.n8162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_14_25_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.rx.i2_2_lut_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__50048),
            .in2(_gnd_net_),
            .in3(N__39314),
            .lcout(),
            .ltout(\c0.rx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21269_4_lut_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.rx.i21269_4_lut_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21269_4_lut_LC_14_25_1 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \c0.rx.i21269_4_lut_LC_14_25_1  (
            .in0(N__50161),
            .in1(N__49962),
            .in2(N__39282),
            .in3(N__50867),
            .lcout(n14439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1840_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1840_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1840_LC_14_25_2 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1840_LC_14_25_2  (
            .in0(N__43709),
            .in1(N__39258),
            .in2(N__43842),
            .in3(N__43445),
            .lcout(),
            .ltout(\c0.n24302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1896_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1896_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1896_LC_14_25_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \c0.i1_4_lut_adj_1896_LC_14_25_3  (
            .in0(N__43667),
            .in1(N__39219),
            .in2(N__39210),
            .in3(N__43531),
            .lcout(\c0.n4_adj_4721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1939_LC_14_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1939_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1939_LC_14_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1939_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__39207),
            .in2(_gnd_net_),
            .in3(N__47827),
            .lcout(\c0.n8_adj_4556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i18_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_14_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_14_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__39745),
            .in2(_gnd_net_),
            .in3(N__48986),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78729),
            .ce(),
            .sr(N__39717));
    defparam \c0.FRAME_MATCHER_state_i12_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_14_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_14_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_14_27_0  (
            .in0(_gnd_net_),
            .in1(N__48988),
            .in2(_gnd_net_),
            .in3(N__39694),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78742),
            .ce(),
            .sr(N__39672));
    defparam \c0.FRAME_MATCHER_state_i19_LC_14_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_14_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_14_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_14_28_0  (
            .in0(_gnd_net_),
            .in1(N__49129),
            .in2(_gnd_net_),
            .in3(N__48990),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78755),
            .ce(),
            .sr(N__39657));
    defparam \c0.i1_2_lut_3_lut_adj_1999_LC_15_8_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1999_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1999_LC_15_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1999_LC_15_8_7  (
            .in0(N__39529),
            .in1(N__39595),
            .in2(_gnd_net_),
            .in3(N__39779),
            .lcout(\c0.n22785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i15_LC_15_9_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i15_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i15_LC_15_9_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i15_LC_15_9_1  (
            .in0(N__39567),
            .in1(N__47724),
            .in2(_gnd_net_),
            .in3(N__39542),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78732),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i5_LC_15_9_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i5_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i5_LC_15_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i5_LC_15_9_3  (
            .in0(N__45381),
            .in1(N__39504),
            .in2(_gnd_net_),
            .in3(N__47725),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78732),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14227_2_lut_3_lut_LC_15_9_4 .C_ON=1'b0;
    defparam \c0.i14227_2_lut_3_lut_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14227_2_lut_3_lut_LC_15_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i14227_2_lut_3_lut_LC_15_9_4  (
            .in0(N__74279),
            .in1(N__74643),
            .in2(_gnd_net_),
            .in3(N__74441),
            .lcout(\c0.n17830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1915_LC_15_10_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1915_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1915_LC_15_10_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i13_4_lut_adj_1915_LC_15_10_0  (
            .in0(N__49155),
            .in1(N__51627),
            .in2(N__57159),
            .in3(N__61335),
            .lcout(),
            .ltout(\c0.n30_adj_4730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1931_LC_15_10_1 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1931_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1931_LC_15_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_1931_LC_15_10_1  (
            .in0(N__48570),
            .in1(N__44439),
            .in2(N__39498),
            .in3(N__51252),
            .lcout(\c0.n17539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_15_10_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_15_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_15_10_3  (
            .in0(N__40021),
            .in1(N__44345),
            .in2(N__39989),
            .in3(N__42655),
            .lcout(\c0.n31_adj_4325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_1_i3_2_lut_LC_15_10_4 .C_ON=1'b0;
    defparam \c0.select_367_Select_1_i3_2_lut_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_1_i3_2_lut_LC_15_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_1_i3_2_lut_LC_15_10_4  (
            .in0(N__74447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71538),
            .lcout(\c0.n3_adj_4434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1313_LC_15_11_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1313_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1313_LC_15_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1313_LC_15_11_0  (
            .in0(N__45382),
            .in1(N__45626),
            .in2(N__42788),
            .in3(N__43285),
            .lcout(\c0.n22775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i9_LC_15_11_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i9_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i9_LC_15_11_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter0.count_i0_i9_LC_15_11_1  (
            .in0(N__39891),
            .in1(_gnd_net_),
            .in2(N__47733),
            .in3(N__42657),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78706),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i21_LC_15_11_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i21_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i21_LC_15_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i21_LC_15_11_2  (
            .in0(N__45655),
            .in1(N__39885),
            .in2(_gnd_net_),
            .in3(N__47716),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1294_LC_15_11_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1294_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1294_LC_15_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1294_LC_15_11_4  (
            .in0(N__39879),
            .in1(N__39848),
            .in2(_gnd_net_),
            .in3(N__39798),
            .lcout(\c0.n13422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1756_LC_15_11_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1756_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1756_LC_15_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1756_LC_15_11_5  (
            .in0(N__44686),
            .in1(N__45173),
            .in2(_gnd_net_),
            .in3(N__40204),
            .lcout(\c0.n13630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i17_LC_15_11_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i17_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i17_LC_15_11_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i17_LC_15_11_6  (
            .in0(N__40205),
            .in1(N__47715),
            .in2(_gnd_net_),
            .in3(N__39762),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_15_12_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_15_12_0 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_15_12_0  (
            .in0(N__41055),
            .in1(N__40854),
            .in2(N__40836),
            .in3(N__40611),
            .lcout(\c0.n25062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1320_LC_15_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1320_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1320_LC_15_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1320_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__43275),
            .in2(_gnd_net_),
            .in3(N__42262),
            .lcout(\c0.n22635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1255_LC_15_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1255_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1255_LC_15_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1255_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__45116),
            .in2(_gnd_net_),
            .in3(N__42143),
            .lcout(\c0.n6_adj_4276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1317_LC_15_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1317_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1317_LC_15_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1317_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__42380),
            .in2(_gnd_net_),
            .in3(N__40206),
            .lcout(\c0.n13558 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i31_LC_15_12_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i31_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i31_LC_15_12_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \quad_counter1.count_i0_i31_LC_15_12_5  (
            .in0(N__40314),
            .in1(N__40590),
            .in2(N__40566),
            .in3(_gnd_net_),
            .lcout(encoder1_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78694),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i19_LC_15_12_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i19_LC_15_12_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i19_LC_15_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i19_LC_15_12_6  (
            .in0(N__47611),
            .in1(N__40284),
            .in2(_gnd_net_),
            .in3(N__42381),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78694),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i90_LC_15_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i90_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i90_LC_15_12_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i90_LC_15_12_7  (
            .in0(N__76613),
            .in1(N__73651),
            .in2(N__65286),
            .in3(N__75195),
            .lcout(\c0.data_in_frame_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78694),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1777_LC_15_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1777_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1777_LC_15_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1777_LC_15_13_1  (
            .in0(N__40274),
            .in1(N__42389),
            .in2(_gnd_net_),
            .in3(N__40214),
            .lcout(\c0.n22580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1256_LC_15_13_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1256_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1256_LC_15_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1256_LC_15_13_2  (
            .in0(N__40178),
            .in1(N__40128),
            .in2(N__40094),
            .in3(N__40038),
            .lcout(\c0.n10467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_15_13_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_15_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i28_LC_15_13_3  (
            .in0(N__50437),
            .in1(N__76997),
            .in2(_gnd_net_),
            .in3(N__48666),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1284_LC_15_13_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1284_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1284_LC_15_13_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1284_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__46349),
            .in2(_gnd_net_),
            .in3(N__46444),
            .lcout(\c0.n21441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__1__5476_LC_15_13_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__1__5476_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__1__5476_LC_15_13_5 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_frame_6__1__5476_LC_15_13_5  (
            .in0(N__48086),
            .in1(N__41276),
            .in2(N__41334),
            .in3(N__46094),
            .lcout(data_out_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__4__5449_LC_15_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__4__5449_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__4__5449_LC_15_13_6 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_frame_9__4__5449_LC_15_13_6  (
            .in0(N__46092),
            .in1(N__48087),
            .in2(N__45267),
            .in3(N__42923),
            .lcout(data_out_frame_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__2__5291_LC_15_13_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__2__5291_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__2__5291_LC_15_13_7 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_29__2__5291_LC_15_13_7  (
            .in0(N__48085),
            .in1(N__46093),
            .in2(N__41261),
            .in3(N__41865),
            .lcout(data_out_frame_29_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1300_LC_15_14_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1300_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1300_LC_15_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1300_LC_15_14_0  (
            .in0(N__41907),
            .in1(N__44864),
            .in2(N__45285),
            .in3(N__41241),
            .lcout(\c0.n24113 ),
            .ltout(\c0.n24113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2019_LC_15_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2019_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2019_LC_15_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2019_LC_15_14_1  (
            .in0(N__41181),
            .in1(N__44899),
            .in2(N__41235),
            .in3(N__50527),
            .lcout(\c0.n21349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1436_LC_15_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1436_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1436_LC_15_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1436_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__41231),
            .in2(_gnd_net_),
            .in3(N__46484),
            .lcout(\c0.n21358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2021_LC_15_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2021_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2021_LC_15_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2021_LC_15_14_3  (
            .in0(N__41180),
            .in1(N__44900),
            .in2(N__41115),
            .in3(N__41066),
            .lcout(\c0.n21311 ),
            .ltout(\c0.n21311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_2050_LC_15_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_2050_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_2050_LC_15_14_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_2050_LC_15_14_4  (
            .in0(N__46270),
            .in1(_gnd_net_),
            .in2(N__41670),
            .in3(N__46815),
            .lcout(),
            .ltout(\c0.n21273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__6__5295_LC_15_14_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__6__5295_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__6__5295_LC_15_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__6__5295_LC_15_14_5  (
            .in0(N__41667),
            .in1(N__41646),
            .in2(N__41625),
            .in3(N__46461),
            .lcout(\c0.data_out_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78663),
            .ce(N__45041),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_15_14_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_15_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_15_14_6  (
            .in0(N__43223),
            .in1(N__41622),
            .in2(_gnd_net_),
            .in3(N__41610),
            .lcout(\c0.n26_adj_4702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1797_LC_15_15_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1797_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1797_LC_15_15_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1797_LC_15_15_0  (
            .in0(N__41588),
            .in1(N__41454),
            .in2(N__46264),
            .in3(N__41922),
            .lcout(),
            .ltout(\c0.n18_adj_4684_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1798_LC_15_15_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1798_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1798_LC_15_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1798_LC_15_15_1  (
            .in0(N__41571),
            .in1(N__45098),
            .in2(N__41541),
            .in3(N__41538),
            .lcout(),
            .ltout(\c0.n20_adj_4685_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__7__5294_LC_15_15_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__7__5294_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__7__5294_LC_15_15_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__7__5294_LC_15_15_2  (
            .in0(N__41945),
            .in1(N__41517),
            .in2(N__41505),
            .in3(N__41502),
            .lcout(\c0.data_out_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78651),
            .ce(N__45055),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1743_LC_15_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1743_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1743_LC_15_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1743_LC_15_15_3  (
            .in0(N__46139),
            .in1(N__46498),
            .in2(_gnd_net_),
            .in3(N__46151),
            .lcout(\c0.n22461 ),
            .ltout(\c0.n22461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1440_LC_15_15_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1440_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1440_LC_15_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1440_LC_15_15_4  (
            .in0(N__41447),
            .in1(N__46716),
            .in2(N__41436),
            .in3(N__41921),
            .lcout(),
            .ltout(\c0.n14_adj_4478_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1470_LC_15_15_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1470_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1470_LC_15_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1470_LC_15_15_5  (
            .in0(N__41433),
            .in1(N__41944),
            .in2(N__41925),
            .in3(N__46539),
            .lcout(data_out_frame_29__2__N_1748),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1438_LC_15_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1438_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1438_LC_15_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1438_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__46533),
            .in2(_gnd_net_),
            .in3(N__46460),
            .lcout(\c0.n22193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1888_LC_15_16_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1888_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1888_LC_15_16_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1888_LC_15_16_0  (
            .in0(N__41913),
            .in1(N__46632),
            .in2(N__41877),
            .in3(N__41861),
            .lcout(\c0.n19_adj_4720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i96_LC_15_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i96_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i96_LC_15_16_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i96_LC_15_16_1  (
            .in0(N__73520),
            .in1(N__76625),
            .in2(N__76398),
            .in3(N__55611),
            .lcout(\c0.data_in_frame_11_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_15_16_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_15_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_15_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i10_LC_15_16_2  (
            .in0(N__50424),
            .in1(N__41837),
            .in2(_gnd_net_),
            .in3(N__43367),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_15_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_15_16_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i4_LC_15_16_3  (
            .in0(N__41700),
            .in1(N__50423),
            .in2(_gnd_net_),
            .in3(N__42123),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__3__5290_LC_15_16_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__3__5290_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__3__5290_LC_15_16_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_out_frame_29__3__5290_LC_15_16_5  (
            .in0(N__46078),
            .in1(N__48188),
            .in2(N__41801),
            .in3(N__46670),
            .lcout(data_out_frame_29_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__4__5425_LC_15_16_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__4__5425_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__4__5425_LC_15_16_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_12__4__5425_LC_15_16_6  (
            .in0(N__48187),
            .in1(N__46079),
            .in2(N__41781),
            .in3(N__41714),
            .lcout(data_out_frame_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_LC_15_16_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_LC_15_16_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i4_2_lut_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__41699),
            .in2(_gnd_net_),
            .in3(N__42064),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_15_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_15_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i29_LC_15_17_0  (
            .in0(N__71916),
            .in1(N__50427),
            .in2(_gnd_net_),
            .in3(N__42093),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i93_LC_15_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i93_LC_15_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i93_LC_15_17_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i93_LC_15_17_1  (
            .in0(N__76624),
            .in1(N__73522),
            .in2(N__70774),
            .in3(N__71917),
            .lcout(\c0.data_in_frame_11_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i23_LC_15_17_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i23_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i23_LC_15_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i23_LC_15_17_2  (
            .in0(N__47721),
            .in1(N__42078),
            .in2(_gnd_net_),
            .in3(N__42701),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i224_LC_15_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i224_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i224_LC_15_17_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i224_LC_15_17_3  (
            .in0(N__79464),
            .in1(N__76355),
            .in2(N__56560),
            .in3(N__76653),
            .lcout(\c0.data_in_frame_27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_15_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_15_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i9_LC_15_17_4  (
            .in0(N__50425),
            .in1(N__42065),
            .in2(_gnd_net_),
            .in3(N__42194),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i217_LC_15_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i217_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i217_LC_15_17_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i217_LC_15_17_5  (
            .in0(N__79463),
            .in1(N__80616),
            .in2(N__75678),
            .in3(N__76652),
            .lcout(\c0.data_in_frame_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i8_LC_15_17_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i8_LC_15_17_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i8_LC_15_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i8_LC_15_17_6  (
            .in0(N__47722),
            .in1(N__42042),
            .in2(_gnd_net_),
            .in3(N__42855),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_LC_15_17_7 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_LC_15_17_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.rx.i3_4_lut_LC_15_17_7  (
            .in0(N__42026),
            .in1(N__50034),
            .in2(N__50183),
            .in3(N__49940),
            .lcout(\c0.rx.n12909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i236_LC_15_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i236_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i236_LC_15_18_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i236_LC_15_18_0  (
            .in0(N__77045),
            .in1(N__56480),
            .in2(N__47408),
            .in3(N__75326),
            .lcout(\c0.data_in_frame_29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1363_LC_15_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1363_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1363_LC_15_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1363_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__43396),
            .in2(_gnd_net_),
            .in3(N__42559),
            .lcout(),
            .ltout(\c0.n22199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1383_LC_15_18_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1383_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1383_LC_15_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1383_LC_15_18_2  (
            .in0(N__42390),
            .in1(N__42845),
            .in2(N__42354),
            .in3(N__42207),
            .lcout(\c0.n22834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1360_LC_15_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1360_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1360_LC_15_18_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1360_LC_15_18_3  (
            .in0(N__42288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47456),
            .lcout(\c0.n13665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_15_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_15_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1752_LC_15_18_5  (
            .in0(N__47051),
            .in1(N__42688),
            .in2(_gnd_net_),
            .in3(N__42261),
            .lcout(\c0.n6_adj_4366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_15_18_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_15_18_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i17_LC_15_18_6  (
            .in0(N__42193),
            .in1(N__50404),
            .in2(_gnd_net_),
            .in3(N__49425),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14131_2_lut_3_lut_LC_15_18_7 .C_ON=1'b0;
    defparam \c0.i14131_2_lut_3_lut_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14131_2_lut_3_lut_LC_15_18_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i14131_2_lut_3_lut_LC_15_18_7  (
            .in0(N__50403),
            .in1(N__50208),
            .in2(_gnd_net_),
            .in3(N__53802),
            .lcout(\c0.n17734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i7_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i7_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i7_LC_15_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i7_LC_15_19_0  (
            .in0(N__42597),
            .in1(N__71133),
            .in2(_gnd_net_),
            .in3(N__47351),
            .lcout(control_mode_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1336_LC_15_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1336_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1336_LC_15_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1336_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__46949),
            .in2(_gnd_net_),
            .in3(N__45340),
            .lcout(),
            .ltout(\c0.n22256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1270_LC_15_19_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1270_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1270_LC_15_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1270_LC_15_19_2  (
            .in0(N__42170),
            .in1(N__42726),
            .in2(N__42150),
            .in3(N__47276),
            .lcout(\c0.n22772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_15_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_15_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i12_LC_15_19_3  (
            .in0(N__50483),
            .in1(N__42121),
            .in2(_gnd_net_),
            .in3(N__46920),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i4_LC_15_19_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i4_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i4_LC_15_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i4_LC_15_19_4  (
            .in0(N__43274),
            .in1(N__60573),
            .in2(_gnd_net_),
            .in3(N__47350),
            .lcout(control_mode_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21015_3_lut_LC_15_19_5 .C_ON=1'b0;
    defparam \c0.i21015_3_lut_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21015_3_lut_LC_15_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i21015_3_lut_LC_15_19_5  (
            .in0(N__43186),
            .in1(N__42924),
            .in2(_gnd_net_),
            .in3(N__42909),
            .lcout(\c0.n24782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i0_LC_15_19_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i0_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i0_LC_15_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i0_LC_15_19_6  (
            .in0(N__45158),
            .in1(N__61068),
            .in2(_gnd_net_),
            .in3(N__47349),
            .lcout(control_mode_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78652),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1321_LC_15_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1321_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1321_LC_15_19_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1321_LC_15_19_7  (
            .in0(N__42703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42856),
            .lcout(\c0.n22423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1268_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1268_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1268_LC_15_20_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1268_LC_15_20_0  (
            .in0(N__47053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42787),
            .lcout(\c0.n6_adj_4293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1382_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1382_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1382_LC_15_20_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1382_LC_15_20_1  (
            .in0(N__42702),
            .in1(N__47052),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n22385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1304_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1304_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1304_LC_15_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1304_LC_15_20_2  (
            .in0(N__42659),
            .in1(N__42601),
            .in2(N__42570),
            .in3(N__42560),
            .lcout(\c0.n20325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_15_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_15_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_15_20_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i14_LC_15_20_3  (
            .in0(N__42427),
            .in1(N__50464),
            .in2(_gnd_net_),
            .in3(N__42471),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i225_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i225_LC_15_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i225_LC_15_20_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i225_LC_15_20_4  (
            .in0(N__80605),
            .in1(N__80094),
            .in2(N__51800),
            .in3(N__79420),
            .lcout(\c0.data_in_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13969_2_lut_LC_15_20_5 .C_ON=1'b0;
    defparam \c0.rx.i13969_2_lut_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13969_2_lut_LC_15_20_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.rx.i13969_2_lut_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49730),
            .in3(N__49648),
            .lcout(n17571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_107_i4_2_lut_LC_15_20_6 .C_ON=1'b0;
    defparam \c0.rx.equal_107_i4_2_lut_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_107_i4_2_lut_LC_15_20_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.rx.equal_107_i4_2_lut_LC_15_20_6  (
            .in0(N__49649),
            .in1(N__49723),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n4_adj_4762),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i6_LC_15_20_7 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i6_LC_15_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i6_LC_15_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i6_LC_15_20_7  (
            .in0(N__43395),
            .in1(N__58056),
            .in2(_gnd_net_),
            .in3(N__47348),
            .lcout(control_mode_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i195_LC_15_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i195_LC_15_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i195_LC_15_21_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i195_LC_15_21_1  (
            .in0(N__67532),
            .in1(N__79084),
            .in2(N__72996),
            .in3(N__79366),
            .lcout(\c0.data_in_frame_24_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14114_2_lut_LC_15_21_2 .C_ON=1'b0;
    defparam \c0.i14114_2_lut_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14114_2_lut_LC_15_21_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i14114_2_lut_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__53894),
            .in2(_gnd_net_),
            .in3(N__49828),
            .lcout(\c0.n937 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_15_21_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i2_LC_15_21_3  (
            .in0(N__50458),
            .in1(N__43347),
            .in2(_gnd_net_),
            .in3(N__43371),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_15_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_15_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_15_21_4 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \c0.data_in_0___i27_LC_15_21_4  (
            .in0(N__79083),
            .in1(N__50459),
            .in2(N__43328),
            .in3(_gnd_net_),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19184_3_lut_LC_15_21_5 .C_ON=1'b0;
    defparam \c0.i19184_3_lut_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i19184_3_lut_LC_15_21_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.i19184_3_lut_LC_15_21_5  (
            .in0(N__44046),
            .in1(N__44158),
            .in2(_gnd_net_),
            .in3(N__44269),
            .lcout(\c0.n17856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i155_LC_15_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i155_LC_15_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i155_LC_15_21_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i155_LC_15_21_6  (
            .in0(N__76675),
            .in1(N__80428),
            .in2(N__79141),
            .in3(N__63328),
            .lcout(\c0.data_in_frame_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i173_LC_15_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i173_LC_15_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i173_LC_15_21_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0__i173_LC_15_21_7  (
            .in0(N__67640),
            .in1(_gnd_net_),
            .in2(N__71966),
            .in3(N__66746),
            .lcout(data_in_frame_21_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_LC_15_22_0 .C_ON=1'b0;
    defparam \c0.i13_2_lut_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_LC_15_22_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i13_2_lut_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__53448),
            .in2(_gnd_net_),
            .in3(N__52769),
            .lcout(\c0.n39_adj_4295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_7_i3_2_lut_LC_15_22_2 .C_ON=1'b0;
    defparam \c0.select_367_Select_7_i3_2_lut_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_7_i3_2_lut_LC_15_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_7_i3_2_lut_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__52632),
            .in2(_gnd_net_),
            .in3(N__71428),
            .lcout(\c0.n3_adj_4422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1280_LC_15_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1280_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1280_LC_15_22_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1280_LC_15_22_3  (
            .in0(N__66662),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56148),
            .lcout(\c0.n5_adj_4302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1374_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1374_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1374_LC_15_22_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1374_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__63961),
            .in2(_gnd_net_),
            .in3(N__63507),
            .lcout(\c0.n22577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1484_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1484_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1484_LC_15_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1484_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__47878),
            .in2(_gnd_net_),
            .in3(N__43604),
            .lcout(\c0.n74_adj_4525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i11_LC_15_22_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_15_22_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_15_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_15_22_6  (
            .in0(N__47879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49003),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78695),
            .ce(),
            .sr(N__47850));
    defparam \c0.i1_2_lut_3_lut_adj_1988_LC_15_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1988_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1988_LC_15_23_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1988_LC_15_23_1  (
            .in0(N__62253),
            .in1(N__74666),
            .in2(_gnd_net_),
            .in3(N__74470),
            .lcout(\c0.n4_adj_4266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1246_LC_15_23_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1246_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1246_LC_15_23_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \c0.i2_4_lut_adj_1246_LC_15_23_2  (
            .in0(N__74469),
            .in1(N__74382),
            .in2(N__74674),
            .in3(N__49552),
            .lcout(\c0.n23912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14109_2_lut_3_lut_LC_15_23_4 .C_ON=1'b0;
    defparam \c0.i14109_2_lut_3_lut_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14109_2_lut_3_lut_LC_15_23_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \c0.i14109_2_lut_3_lut_LC_15_23_4  (
            .in0(N__53909),
            .in1(N__80924),
            .in2(_gnd_net_),
            .in3(N__49553),
            .lcout(\c0.n3844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_2030_LC_15_23_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_2030_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_2030_LC_15_23_5 .LUT_INIT=16'b0000000011001101;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_2030_LC_15_23_5  (
            .in0(N__49554),
            .in1(N__53910),
            .in2(N__80951),
            .in3(N__44277),
            .lcout(),
            .ltout(\c0.n22098_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1286_LC_15_23_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1286_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1286_LC_15_23_6 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \c0.i1_4_lut_adj_1286_LC_15_23_6  (
            .in0(N__53911),
            .in1(N__49827),
            .in2(N__44238),
            .in3(N__48483),
            .lcout(),
            .ltout(\c0.n63_adj_4305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_15_23_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_15_23_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i0_LC_15_23_7 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_15_23_7  (
            .in0(N__44013),
            .in1(N__44235),
            .in2(N__44229),
            .in3(N__44194),
            .lcout(\c0.FRAME_MATCHER_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78707),
            .ce(),
            .sr(N__44995));
    defparam \c0.i1_2_lut_4_lut_adj_1996_LC_15_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1996_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1996_LC_15_24_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1996_LC_15_24_0  (
            .in0(N__44109),
            .in1(N__44057),
            .in2(N__44012),
            .in3(N__43530),
            .lcout(\c0.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1906_LC_15_24_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1906_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1906_LC_15_24_5 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \c0.i2_4_lut_adj_1906_LC_15_24_5  (
            .in0(N__43924),
            .in1(N__43869),
            .in2(N__49755),
            .in3(N__43837),
            .lcout(),
            .ltout(\c0.n24591_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_15_24_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_15_24_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i2_LC_15_24_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_15_24_6  (
            .in0(N__43710),
            .in1(N__43671),
            .in2(N__43638),
            .in3(N__43635),
            .lcout(\c0.FRAME_MATCHER_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78717),
            .ce(),
            .sr(N__45027));
    defparam \c0.FRAME_MATCHER_state_i15_LC_15_25_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_15_25_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_15_25_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(N__43598),
            .in2(_gnd_net_),
            .in3(N__48979),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78731),
            .ce(),
            .sr(N__43563));
    defparam \c0.FRAME_MATCHER_state_i1_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_15_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i1_LC_15_26_0 .LUT_INIT=16'b1101110111011100;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_15_26_0  (
            .in0(N__49786),
            .in1(N__43551),
            .in2(N__43545),
            .in3(N__43532),
            .lcout(\c0.FRAME_MATCHER_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78743),
            .ce(),
            .sr(N__45028));
    defparam \c0.FRAME_MATCHER_state_i20_LC_15_27_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_15_27_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_15_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_15_27_5  (
            .in0(_gnd_net_),
            .in1(N__44314),
            .in2(_gnd_net_),
            .in3(N__48999),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78756),
            .ce(),
            .sr(N__44292));
    defparam \c0.equal_88_i9_2_lut_3_lut_LC_16_6_0 .C_ON=1'b0;
    defparam \c0.equal_88_i9_2_lut_3_lut_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.equal_88_i9_2_lut_3_lut_LC_16_6_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.equal_88_i9_2_lut_3_lut_LC_16_6_0  (
            .in0(N__74344),
            .in1(N__74480),
            .in2(_gnd_net_),
            .in3(N__74636),
            .lcout(\c0.n9_adj_4273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i200_LC_16_8_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i200_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i200_LC_16_8_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i200_LC_16_8_0  (
            .in0(N__72860),
            .in1(N__76324),
            .in2(N__52071),
            .in3(N__79483),
            .lcout(\c0.data_in_frame_24_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i65_LC_16_8_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i65_LC_16_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i65_LC_16_8_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i65_LC_16_8_1  (
            .in0(N__80707),
            .in1(N__73596),
            .in2(N__61548),
            .in3(N__72861),
            .lcout(\c0.data_in_frame_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i215_LC_16_8_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i215_LC_16_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i215_LC_16_8_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i215_LC_16_8_2  (
            .in0(N__69166),
            .in1(N__73155),
            .in2(N__75989),
            .in3(N__79484),
            .lcout(\c0.data_in_frame_26_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i154_LC_16_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i154_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i154_LC_16_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i154_LC_16_8_5  (
            .in0(N__76623),
            .in1(N__80398),
            .in2(N__63412),
            .in3(N__75243),
            .lcout(\c0.data_in_frame_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i82_LC_16_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i82_LC_16_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i82_LC_16_8_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i82_LC_16_8_6  (
            .in0(N__73595),
            .in1(N__75244),
            .in2(N__69200),
            .in3(N__55070),
            .lcout(\c0.data_in_frame_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_16_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_16_8_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i9_LC_16_8_7  (
            .in0(N__70151),
            .in1(N__74069),
            .in2(N__80739),
            .in3(N__61035),
            .lcout(data_in_frame_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_16_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_16_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_16_9_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_16_9_0  (
            .in0(N__76622),
            .in1(N__70152),
            .in2(N__54950),
            .in3(N__75242),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1904_LC_16_9_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1904_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1904_LC_16_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1904_LC_16_9_1  (
            .in0(N__70299),
            .in1(N__51336),
            .in2(N__61176),
            .in3(N__71100),
            .lcout(\c0.n20_adj_4726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_16_9_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_16_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i7_LC_16_9_3  (
            .in0(N__50401),
            .in1(N__44565),
            .in2(_gnd_net_),
            .in3(N__44513),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_16_9_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_16_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i31_LC_16_9_6  (
            .in0(N__73153),
            .in1(N__50402),
            .in2(_gnd_net_),
            .in3(N__44466),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_16_9_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_16_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_16_9_7 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_16_9_7  (
            .in0(N__44588),
            .in1(N__73154),
            .in2(N__50864),
            .in3(N__49389),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1929_LC_16_10_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1929_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1929_LC_16_10_1 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \c0.i10_4_lut_adj_1929_LC_16_10_1  (
            .in0(N__48594),
            .in1(N__61142),
            .in2(N__44448),
            .in3(N__68217),
            .lcout(\c0.n27_adj_4735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_2_i3_2_lut_LC_16_10_3 .C_ON=1'b0;
    defparam \c0.select_367_Select_2_i3_2_lut_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_2_i3_2_lut_LC_16_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_2_i3_2_lut_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__74659),
            .in2(_gnd_net_),
            .in3(N__71542),
            .lcout(\c0.n3_adj_4432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_74_i9_2_lut_3_lut_LC_16_10_7 .C_ON=1'b0;
    defparam \c0.equal_74_i9_2_lut_3_lut_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.equal_74_i9_2_lut_3_lut_LC_16_10_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.equal_74_i9_2_lut_3_lut_LC_16_10_7  (
            .in0(N__74365),
            .in1(N__74498),
            .in2(_gnd_net_),
            .in3(N__74658),
            .lcout(\c0.n9_adj_4601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_2__I_0_2_lut_LC_16_11_0 .C_ON=1'b0;
    defparam \c0.control_mode_2__I_0_2_lut_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.control_mode_2__I_0_2_lut_LC_16_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.control_mode_2__I_0_2_lut_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__47294),
            .in2(_gnd_net_),
            .in3(N__47012),
            .lcout(\c0.data_out_frame_29__7__N_735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1362_LC_16_11_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1362_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1362_LC_16_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1362_LC_16_11_1  (
            .in0(N__47293),
            .in1(N__44830),
            .in2(N__45323),
            .in3(N__44405),
            .lcout(\c0.n22754 ),
            .ltout(\c0.n22754_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1318_LC_16_11_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1318_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1318_LC_16_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1318_LC_16_11_2  (
            .in0(N__44363),
            .in1(N__45627),
            .in2(N__44352),
            .in3(N__44808),
            .lcout(\c0.n22243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1298_LC_16_11_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1298_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1298_LC_16_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1298_LC_16_11_3  (
            .in0(N__47298),
            .in1(N__44910),
            .in2(N__44802),
            .in3(N__45262),
            .lcout(\c0.n10477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i18_LC_16_11_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i18_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i18_LC_16_11_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \quad_counter0.count_i0_i18_LC_16_11_4  (
            .in0(N__44880),
            .in1(_gnd_net_),
            .in2(N__44846),
            .in3(N__47720),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78718),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1759_LC_16_11_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1759_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1759_LC_16_11_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1759_LC_16_11_5  (
            .in0(N__47013),
            .in1(_gnd_net_),
            .in2(N__47305),
            .in3(N__44831),
            .lcout(\c0.n22641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1316_LC_16_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1316_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1316_LC_16_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1316_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__47011),
            .in2(_gnd_net_),
            .in3(N__45184),
            .lcout(\c0.n22583 ),
            .ltout(\c0.n22583_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1292_LC_16_11_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1292_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1292_LC_16_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1292_LC_16_11_7  (
            .in0(N__44798),
            .in1(N__44769),
            .in2(N__44718),
            .in3(N__44703),
            .lcout(\c0.n13872 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i20_LC_16_12_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i20_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i20_LC_16_12_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \quad_counter0.count_i0_i20_LC_16_12_2  (
            .in0(N__47612),
            .in1(_gnd_net_),
            .in2(N__44607),
            .in3(N__45322),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1720_LC_16_12_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1720_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1720_LC_16_12_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1720_LC_16_12_3  (
            .in0(N__61391),
            .in1(N__62244),
            .in2(_gnd_net_),
            .in3(N__75327),
            .lcout(n22101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_16_12_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_16_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_16_12_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_16_12_4  (
            .in0(N__44589),
            .in1(N__76154),
            .in2(N__50913),
            .in3(N__50718),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1315_LC_16_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1315_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1315_LC_16_12_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1315_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__45648),
            .in2(_gnd_net_),
            .in3(N__46954),
            .lcout(\c0.n22252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__3__5474_LC_16_12_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__3__5474_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__3__5474_LC_16_12_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_out_frame_6__3__5474_LC_16_12_6  (
            .in0(N__48077),
            .in1(N__46031),
            .in2(N__45615),
            .in3(N__45533),
            .lcout(data_out_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1405_LC_16_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1405_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1405_LC_16_13_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1405_LC_16_13_0  (
            .in0(N__45518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45444),
            .lcout(\c0.n22553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1763_LC_16_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1763_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1763_LC_16_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1763_LC_16_13_1  (
            .in0(N__45392),
            .in1(N__46955),
            .in2(_gnd_net_),
            .in3(N__45321),
            .lcout(\c0.n22689 ),
            .ltout(\c0.n22689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1338_LC_16_13_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1338_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1338_LC_16_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1338_LC_16_13_2  (
            .in0(N__45276),
            .in1(N__45260),
            .in2(N__45192),
            .in3(N__45185),
            .lcout(\c0.n10455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_16_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_16_14_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_LC_16_14_0  (
            .in0(N__46483),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46272),
            .lcout(\c0.n22522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2048_LC_16_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2048_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2048_LC_16_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2048_LC_16_14_1  (
            .in0(N__46271),
            .in1(N__46553),
            .in2(N__46827),
            .in3(N__46482),
            .lcout(\c0.n20312 ),
            .ltout(\c0.n20312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1749_LC_16_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1749_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1749_LC_16_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1749_LC_16_14_2  (
            .in0(N__46500),
            .in1(N__46879),
            .in2(N__45087),
            .in3(N__46822),
            .lcout(),
            .ltout(\c0.n6_adj_4674_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__4__5289_LC_16_14_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__4__5289_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__4__5289_LC_16_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_29__4__5289_LC_16_14_3  (
            .in0(N__45084),
            .in1(N__46704),
            .in2(N__45078),
            .in3(N__46743),
            .lcout(\c0.data_out_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78679),
            .ce(N__45037),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1275_LC_16_14_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1275_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1275_LC_16_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1275_LC_16_14_4  (
            .in0(N__46742),
            .in1(N__46631),
            .in2(_gnd_net_),
            .in3(N__46614),
            .lcout(\c0.n20786 ),
            .ltout(\c0.n20786_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1451_LC_16_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1451_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1451_LC_16_14_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_1451_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46542),
            .in3(N__46499),
            .lcout(\c0.n9_adj_4494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1344_LC_16_14_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1344_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1344_LC_16_14_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1344_LC_16_14_6  (
            .in0(N__46741),
            .in1(N__46184),
            .in2(N__46485),
            .in3(N__46532),
            .lcout(\c0.n21433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2023_LC_16_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2023_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2023_LC_16_14_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2023_LC_16_14_7  (
            .in0(N__46183),
            .in1(N__46478),
            .in2(N__46826),
            .in3(N__46740),
            .lcout(\c0.n12590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1655_LC_16_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1655_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1655_LC_16_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1655_LC_16_15_0  (
            .in0(N__46449),
            .in1(N__46378),
            .in2(N__46362),
            .in3(N__46254),
            .lcout(\c0.n10531 ),
            .ltout(\c0.n10531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2025_LC_16_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2025_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2025_LC_16_15_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2025_LC_16_15_1  (
            .in0(N__46823),
            .in1(N__46188),
            .in2(N__46158),
            .in3(N__46744),
            .lcout(\c0.n21451 ),
            .ltout(\c0.n21451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1346_LC_16_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1346_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1346_LC_16_15_2 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \c0.i1_2_lut_adj_1346_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__46133),
            .in2(N__46101),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_frame_29__3__N_1730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__6__5455_LC_16_15_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__6__5455_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__6__5455_LC_16_15_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_frame_8__6__5455_LC_16_15_3  (
            .in0(N__48186),
            .in1(N__46090),
            .in2(N__45692),
            .in3(N__47484),
            .lcout(data_out_frame_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__6__I_721_2_lut_LC_16_15_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__6__I_721_2_lut_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_frame_29__6__I_721_2_lut_LC_16_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_frame_29__6__I_721_2_lut_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__46878),
            .in2(_gnd_net_),
            .in3(N__46825),
            .lcout(\c0.data_out_frame_29__6__N_1538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1439_LC_16_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1439_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1439_LC_16_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1439_LC_16_15_5  (
            .in0(N__46824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46745),
            .lcout(\c0.n4_adj_4271 ),
            .ltout(\c0.n4_adj_4271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1251_LC_16_15_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1251_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1251_LC_16_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1251_LC_16_15_6  (
            .in0(N__46710),
            .in1(N__46703),
            .in2(N__46680),
            .in3(N__46677),
            .lcout(data_out_frame_29__3__N_1661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_16_15_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_16_15_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.i1_2_lut_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__47231),
            .in2(_gnd_net_),
            .in3(N__46652),
            .lcout(n12904),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2036_LC_16_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2036_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2036_LC_16_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_2036_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__48768),
            .in2(_gnd_net_),
            .in3(N__47841),
            .lcout(\c0.n21647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1544_LC_16_16_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1544_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1544_LC_16_16_1 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1544_LC_16_16_1  (
            .in0(N__61384),
            .in1(N__62309),
            .in2(_gnd_net_),
            .in3(N__61425),
            .lcout(\c0.n22112 ),
            .ltout(\c0.n22112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i86_LC_16_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i86_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i86_LC_16_16_2 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i86_LC_16_16_2  (
            .in0(N__61582),
            .in1(N__69161),
            .in2(N__46635),
            .in3(N__79791),
            .lcout(\c0.data_in_frame_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i166_LC_16_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i166_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i166_LC_16_16_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i166_LC_16_16_3  (
            .in0(N__80417),
            .in1(N__79984),
            .in2(N__79796),
            .in3(N__56143),
            .lcout(\c0.data_in_frame_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i151_LC_16_16_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i151_LC_16_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i151_LC_16_16_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i151_LC_16_16_4  (
            .in0(N__73214),
            .in1(N__80418),
            .in2(N__61897),
            .in3(N__69162),
            .lcout(\c0.data_in_frame_18_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i102_LC_16_16_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i102_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i102_LC_16_16_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i102_LC_16_16_5  (
            .in0(N__79787),
            .in1(N__73519),
            .in2(N__55742),
            .in3(N__79985),
            .lcout(\c0.data_in_frame_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i124_LC_16_16_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i124_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i124_LC_16_16_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i124_LC_16_16_6  (
            .in0(N__73518),
            .in1(N__80867),
            .in2(N__65426),
            .in3(N__77128),
            .lcout(\c0.data_in_frame_15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_16_16_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_16_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_16_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i20_LC_16_16_7  (
            .in0(N__50454),
            .in1(N__48680),
            .in2(_gnd_net_),
            .in3(N__46906),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_2011_LC_16_17_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_2011_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_2011_LC_16_17_0 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_2011_LC_16_17_0  (
            .in0(N__74673),
            .in1(N__74520),
            .in2(N__74386),
            .in3(N__61424),
            .lcout(\c0.n22099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1783_LC_16_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1783_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1783_LC_16_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1783_LC_16_17_1  (
            .in0(N__66099),
            .in1(N__66569),
            .in2(_gnd_net_),
            .in3(N__65406),
            .lcout(),
            .ltout(\c0.n82_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i61_4_lut_LC_16_17_2 .C_ON=1'b0;
    defparam \c0.i61_4_lut_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i61_4_lut_LC_16_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i61_4_lut_LC_16_17_2  (
            .in0(N__56056),
            .in1(N__66637),
            .in2(N__46887),
            .in3(N__72049),
            .lcout(\c0.n142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i146_LC_16_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i146_LC_16_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i146_LC_16_17_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i146_LC_16_17_3  (
            .in0(N__72050),
            .in1(N__75110),
            .in2(N__69199),
            .in3(N__80420),
            .lcout(\c0.data_in_frame_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i118_LC_16_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i118_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i118_LC_16_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i118_LC_16_17_4  (
            .in0(N__62396),
            .in1(N__59190),
            .in2(_gnd_net_),
            .in3(N__79776),
            .lcout(data_in_frame_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i150_LC_16_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i150_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i150_LC_16_17_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i150_LC_16_17_5  (
            .in0(N__79777),
            .in1(N__80419),
            .in2(N__56072),
            .in3(N__69157),
            .lcout(\c0.data_in_frame_18_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i122_LC_16_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i122_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i122_LC_16_17_7 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i122_LC_16_17_7  (
            .in0(N__80899),
            .in1(N__73521),
            .in2(N__62459),
            .in3(N__75111),
            .lcout(\c0.data_in_frame_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1925_LC_16_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1925_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1925_LC_16_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1925_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__49196),
            .in2(_gnd_net_),
            .in3(N__47837),
            .lcout(\c0.n21629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_1166_LC_16_18_1 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_1166_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_1166_LC_16_18_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_3_lut_adj_1166_LC_16_18_1  (
            .in0(N__47234),
            .in1(N__49718),
            .in2(_gnd_net_),
            .in3(N__49657),
            .lcout(),
            .ltout(\c0.rx.n17834_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i11373_3_lut_LC_16_18_2 .C_ON=1'b0;
    defparam \c0.rx.i11373_3_lut_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i11373_3_lut_LC_16_18_2 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \c0.rx.i11373_3_lut_LC_16_18_2  (
            .in0(N__50153),
            .in1(_gnd_net_),
            .in2(N__47154),
            .in3(N__47151),
            .lcout(n14988),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1445_LC_16_18_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1445_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1445_LC_16_18_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_adj_1445_LC_16_18_3  (
            .in0(N__67884),
            .in1(N__64133),
            .in2(_gnd_net_),
            .in3(N__56632),
            .lcout(\c0.n17_adj_4483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1867_LC_16_18_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1867_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1867_LC_16_18_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1867_LC_16_18_6  (
            .in0(N__56223),
            .in1(N__62296),
            .in2(_gnd_net_),
            .in3(N__75301),
            .lcout(n22103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i5_LC_16_19_0 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i5_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i5_LC_16_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i5_LC_16_19_0  (
            .in0(N__47057),
            .in1(N__60438),
            .in2(_gnd_net_),
            .in3(N__47347),
            .lcout(control_mode_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1520_LC_16_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1520_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1520_LC_16_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1520_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__62397),
            .in2(_gnd_net_),
            .in3(N__62458),
            .lcout(\c0.n4_adj_4352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i1_LC_16_19_2 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i1_LC_16_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i1_LC_16_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i1_LC_16_19_2  (
            .in0(N__47007),
            .in1(N__51237),
            .in2(_gnd_net_),
            .in3(N__47343),
            .lcout(control_mode_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i3_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i3_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i3_LC_16_19_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.control_mode_i0_i3_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__46953),
            .in2(N__47352),
            .in3(N__51480),
            .lcout(control_mode_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i134_LC_16_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i134_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i134_LC_16_19_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i134_LC_16_19_4  (
            .in0(N__79785),
            .in1(N__80421),
            .in2(N__62526),
            .in3(N__72990),
            .lcout(\c0.data_in_frame_16_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78666),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i14_LC_16_19_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i14_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i14_LC_16_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i14_LC_16_19_5  (
            .in0(N__47723),
            .in1(N__47520),
            .in2(_gnd_net_),
            .in3(N__47468),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_16_19_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_16_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_16_19_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_16_19_7  (
            .in0(N__47430),
            .in1(N__78979),
            .in2(N__50912),
            .in3(N__49369),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1442_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1442_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1442_LC_16_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i10_4_lut_adj_1442_LC_16_20_0  (
            .in0(N__51944),
            .in1(N__63942),
            .in2(N__47409),
            .in3(N__51887),
            .lcout(),
            .ltout(\c0.n26_adj_4480_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1447_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1447_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1447_LC_16_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_1447_LC_16_20_1  (
            .in0(N__47739),
            .in1(N__47388),
            .in2(N__47376),
            .in3(N__76710),
            .lcout(\c0.n24539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1507_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1507_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1507_LC_16_20_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i16_4_lut_adj_1507_LC_16_20_2  (
            .in0(N__47373),
            .in1(N__67680),
            .in2(N__56925),
            .in3(N__49533),
            .lcout(),
            .ltout(\c0.n34_adj_4546_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1522_LC_16_20_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1522_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1522_LC_16_20_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i17_4_lut_adj_1522_LC_16_20_3  (
            .in0(N__47241),
            .in1(N__56946),
            .in2(N__47355),
            .in3(N__60000),
            .lcout(n24622),
            .ltout(n24622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i2_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i2_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i2_LC_16_20_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.control_mode_i0_i2_LC_16_20_4  (
            .in0(N__57270),
            .in1(_gnd_net_),
            .in2(N__47319),
            .in3(N__47277),
            .lcout(control_mode_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20968_4_lut_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.i20968_4_lut_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20968_4_lut_LC_16_20_5 .LUT_INIT=16'b0110100100000000;
    LogicCell40 \c0.i20968_4_lut_LC_16_20_5  (
            .in0(N__51888),
            .in1(N__49431),
            .in2(N__59670),
            .in3(N__47247),
            .lcout(\c0.n24733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i157_LC_16_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i157_LC_16_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i157_LC_16_21_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i157_LC_16_21_0  (
            .in0(N__80422),
            .in1(N__76682),
            .in2(N__71967),
            .in3(N__56185),
            .lcout(\c0.data_in_frame_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i238_LC_16_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i238_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i238_LC_16_21_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i238_LC_16_21_1  (
            .in0(N__49446),
            .in1(N__56487),
            .in2(N__79800),
            .in3(N__75337),
            .lcout(\c0.data_in_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1739_LC_16_21_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1739_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1739_LC_16_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1739_LC_16_21_3  (
            .in0(N__75611),
            .in1(N__76749),
            .in2(N__75576),
            .in3(N__63609),
            .lcout(\c0.n18_adj_4485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i199_LC_16_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i199_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i199_LC_16_21_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i199_LC_16_21_4  (
            .in0(N__73207),
            .in1(N__72981),
            .in2(N__67150),
            .in3(N__79361),
            .lcout(\c0.data_in_frame_24_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i207_LC_16_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i207_LC_16_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i207_LC_16_21_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i207_LC_16_21_5  (
            .in0(N__79359),
            .in1(N__74220),
            .in2(N__59629),
            .in3(N__73209),
            .lcout(\c0.data_in_frame_25_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i193_LC_16_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i193_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i193_LC_16_21_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i193_LC_16_21_6  (
            .in0(N__80738),
            .in1(N__72980),
            .in2(N__78017),
            .in3(N__79360),
            .lcout(\c0.data_in_frame_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i135_LC_16_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i135_LC_16_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i135_LC_16_21_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i135_LC_16_21_7  (
            .in0(N__72979),
            .in1(N__80423),
            .in2(N__58930),
            .in3(N__73208),
            .lcout(\c0.data_in_frame_16_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1443_LC_16_22_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1443_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1443_LC_16_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1443_LC_16_22_0  (
            .in0(N__56814),
            .in1(N__59578),
            .in2(N__63877),
            .in3(N__67248),
            .lcout(\c0.n24384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i196_LC_16_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i196_LC_16_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i196_LC_16_22_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i196_LC_16_22_1  (
            .in0(N__76912),
            .in1(N__72942),
            .in2(N__59587),
            .in3(N__79356),
            .lcout(\c0.data_in_frame_24_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1660_LC_16_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1660_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1660_LC_16_22_2 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1660_LC_16_22_2  (
            .in0(N__56241),
            .in1(N__62319),
            .in2(_gnd_net_),
            .in3(N__61433),
            .lcout(\c0.n22134 ),
            .ltout(\c0.n22134_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i222_LC_16_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i222_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i222_LC_16_22_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i222_LC_16_22_3  (
            .in0(N__76694),
            .in1(N__79792),
            .in2(N__47898),
            .in3(N__56886),
            .lcout(\c0.data_in_frame_27_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i214_LC_16_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i214_LC_16_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i214_LC_16_22_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i214_LC_16_22_4  (
            .in0(N__79355),
            .in1(N__79647),
            .in2(N__63878),
            .in3(N__69227),
            .lcout(\c0.data_in_frame_26_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i209_LC_16_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i209_LC_16_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i209_LC_16_22_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i209_LC_16_22_5  (
            .in0(N__69226),
            .in1(N__56588),
            .in2(N__80671),
            .in3(N__79357),
            .lcout(\c0.data_in_frame_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i197_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i197_LC_16_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i197_LC_16_22_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i197_LC_16_22_6  (
            .in0(N__79354),
            .in1(N__71939),
            .in2(N__72977),
            .in3(N__67249),
            .lcout(\c0.data_in_frame_24_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i223_LC_16_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i223_LC_16_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i223_LC_16_22_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i223_LC_16_22_7  (
            .in0(N__76695),
            .in1(N__73210),
            .in2(N__56853),
            .in3(N__79358),
            .lcout(\c0.data_in_frame_27_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1949_LC_16_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1949_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1949_LC_16_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1949_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__47883),
            .in2(_gnd_net_),
            .in3(N__47829),
            .lcout(\c0.n21633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i232_LC_16_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i232_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i232_LC_16_23_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i232_LC_16_23_1  (
            .in0(N__80093),
            .in1(N__76317),
            .in2(N__52241),
            .in3(N__79365),
            .lcout(\c0.data_in_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78719),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1198_LC_16_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1198_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1198_LC_16_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1198_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(N__48416),
            .in2(_gnd_net_),
            .in3(N__47828),
            .lcout(\c0.n21651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i218_LC_16_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i218_LC_16_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i218_LC_16_23_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i218_LC_16_23_3  (
            .in0(N__76687),
            .in1(N__75185),
            .in2(N__64139),
            .in3(N__79364),
            .lcout(\c0.data_in_frame_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78719),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19136_4_lut_LC_16_23_4 .C_ON=1'b0;
    defparam \c0.i19136_4_lut_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19136_4_lut_LC_16_23_4 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \c0.i19136_4_lut_LC_16_23_4  (
            .in0(N__49845),
            .in1(N__52408),
            .in2(N__48528),
            .in3(N__53915),
            .lcout(\c0.n5024 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1543_LC_16_24_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1543_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1543_LC_16_24_3 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i1_4_lut_adj_1543_LC_16_24_3  (
            .in0(N__48482),
            .in1(N__48450),
            .in2(N__48432),
            .in3(N__53803),
            .lcout(\c0.n2119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i31_LC_16_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_16_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_16_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__48412),
            .in2(_gnd_net_),
            .in3(N__48980),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78744),
            .ce(),
            .sr(N__48390));
    defparam \c0.select_367_Select_4_i3_2_lut_LC_17_5_1 .C_ON=1'b0;
    defparam \c0.select_367_Select_4_i3_2_lut_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_4_i3_2_lut_LC_17_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_4_i3_2_lut_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(N__52374),
            .in2(_gnd_net_),
            .in3(N__71553),
            .lcout(\c0.n3_adj_4428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_adj_1941_LC_17_6_6 .C_ON=1'b0;
    defparam \c0.i23_3_lut_adj_1941_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_adj_1941_LC_17_6_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i23_3_lut_adj_1941_LC_17_6_6  (
            .in0(N__60714),
            .in1(N__60588),
            .in2(_gnd_net_),
            .in3(N__49863),
            .lcout(FRAME_MATCHER_state_31_N_2975_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1654_LC_17_7_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1654_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1654_LC_17_7_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1654_LC_17_7_0  (
            .in0(N__48710),
            .in1(N__47904),
            .in2(N__64458),
            .in3(N__48534),
            .lcout(),
            .ltout(\c0.n22_adj_4643_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1674_LC_17_7_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1674_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1674_LC_17_7_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1674_LC_17_7_1  (
            .in0(N__55184),
            .in1(N__55508),
            .in2(N__47910),
            .in3(N__60548),
            .lcout(\c0.n24433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1644_LC_17_7_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1644_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1644_LC_17_7_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1644_LC_17_7_2  (
            .in0(N__55021),
            .in1(N__50984),
            .in2(N__61541),
            .in3(N__50971),
            .lcout(),
            .ltout(\c0.n10_adj_4639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1649_LC_17_7_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1649_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1649_LC_17_7_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1649_LC_17_7_3  (
            .in0(N__55069),
            .in1(N__48744),
            .in2(N__47907),
            .in3(N__50945),
            .lcout(\c0.n13_adj_4640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_1677_LC_17_7_4 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_1677_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_1677_LC_17_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_1677_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(N__57942),
            .in2(_gnd_net_),
            .in3(N__61031),
            .lcout(\c0.n12_adj_4657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1607_LC_17_7_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1607_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1607_LC_17_7_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1607_LC_17_7_5  (
            .in0(N__50972),
            .in1(N__55020),
            .in2(N__50988),
            .in3(N__50944),
            .lcout(\c0.n23666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_adj_1875_LC_17_7_7 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_adj_1875_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_adj_1875_LC_17_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_adj_1875_LC_17_7_7  (
            .in0(N__55220),
            .in1(N__51085),
            .in2(N__57376),
            .in3(N__64764),
            .lcout(\c0.n20_adj_4642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_17_8_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_17_8_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i10_LC_17_8_0  (
            .in0(N__74066),
            .in1(N__70172),
            .in2(N__75254),
            .in3(N__51207),
            .lcout(data_in_frame_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_17_8_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_17_8_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i11_LC_17_8_1  (
            .in0(N__70170),
            .in1(N__74067),
            .in2(N__57244),
            .in3(N__79189),
            .lcout(data_in_frame_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i47_3_lut_4_lut_LC_17_8_2 .C_ON=1'b0;
    defparam \c0.i47_3_lut_4_lut_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i47_3_lut_4_lut_LC_17_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i47_3_lut_4_lut_LC_17_8_2  (
            .in0(N__64614),
            .in1(N__55664),
            .in2(N__55746),
            .in3(N__69903),
            .lcout(\c0.n128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1735_LC_17_8_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1735_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1735_LC_17_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1735_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__50969),
            .in2(_gnd_net_),
            .in3(N__50943),
            .lcout(\c0.n5_adj_4268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_17_8_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_17_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i46_LC_17_8_4  (
            .in0(N__50970),
            .in1(N__79628),
            .in2(_gnd_net_),
            .in3(N__69437),
            .lcout(data_in_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_17_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_17_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i29_LC_17_8_5  (
            .in0(N__70171),
            .in1(N__76550),
            .in2(N__50949),
            .in3(N__71957),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1831_LC_17_8_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1831_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1831_LC_17_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1831_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__51206),
            .in2(_gnd_net_),
            .in3(N__51418),
            .lcout(\c0.n22626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_1603_LC_17_8_7 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_1603_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_1603_LC_17_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_1603_LC_17_8_7  (
            .in0(N__57228),
            .in1(N__51564),
            .in2(_gnd_net_),
            .in3(N__50942),
            .lcout(\c0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_17_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_17_9_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i30_LC_17_9_0  (
            .in0(N__76548),
            .in1(N__70153),
            .in2(N__79677),
            .in3(N__51573),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78758),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1645_LC_17_9_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1645_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1645_LC_17_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1645_LC_17_9_1  (
            .in0(N__54936),
            .in1(N__51211),
            .in2(_gnd_net_),
            .in3(N__57484),
            .lcout(\c0.n23305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_1594_LC_17_9_2 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_1594_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_1594_LC_17_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_1594_LC_17_9_2  (
            .in0(N__71099),
            .in1(N__61030),
            .in2(N__60409),
            .in3(N__58012),
            .lcout(),
            .ltout(\c0.n14_adj_4607_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1832_LC_17_9_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1832_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1832_LC_17_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1832_LC_17_9_3  (
            .in0(N__48542),
            .in1(N__60305),
            .in2(N__48558),
            .in3(N__48554),
            .lcout(\c0.data_out_frame_0__7__N_2626 ),
            .ltout(\c0.data_out_frame_0__7__N_2626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_4_lut_LC_17_9_4 .C_ON=1'b0;
    defparam \c0.i32_4_lut_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i32_4_lut_LC_17_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i32_4_lut_LC_17_9_4  (
            .in0(N__48555),
            .in1(N__51335),
            .in2(N__48546),
            .in3(N__57564),
            .lcout(\c0.n88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_1830_LC_17_9_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_1830_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_1830_LC_17_9_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_1830_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__57232),
            .in2(_gnd_net_),
            .in3(N__60490),
            .lcout(\c0.n30_adj_4585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_4_lut_LC_17_9_6 .C_ON=1'b0;
    defparam \c0.i8_2_lut_4_lut_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_4_lut_LC_17_9_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_2_lut_4_lut_LC_17_9_6  (
            .in0(N__57233),
            .in1(N__60386),
            .in2(N__60533),
            .in3(N__58013),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_3_lut_4_lut_LC_17_9_7 .C_ON=1'b0;
    defparam \c0.i15_2_lut_3_lut_4_lut_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_3_lut_4_lut_LC_17_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_2_lut_3_lut_4_lut_LC_17_9_7  (
            .in0(N__48543),
            .in1(N__51212),
            .in2(N__51465),
            .in3(N__55331),
            .lcout(\c0.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_17_10_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_17_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i49_LC_17_10_0  (
            .in0(N__57593),
            .in1(N__80655),
            .in2(_gnd_net_),
            .in3(N__68442),
            .lcout(data_in_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1243_LC_17_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1243_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1243_LC_17_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1243_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__51562),
            .in2(_gnd_net_),
            .in3(N__57592),
            .lcout(),
            .ltout(\c0.n6_adj_4254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1244_LC_17_10_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1244_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1244_LC_17_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1244_LC_17_10_2  (
            .in0(N__60835),
            .in1(N__60378),
            .in2(N__48573),
            .in3(N__51439),
            .lcout(\c0.n13223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1918_LC_17_10_3 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1918_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1918_LC_17_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i11_4_lut_adj_1918_LC_17_10_3  (
            .in0(N__64346),
            .in1(N__61194),
            .in2(N__51099),
            .in3(N__61860),
            .lcout(\c0.n28_adj_4731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_17_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_17_10_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i31_LC_17_10_4  (
            .in0(N__76549),
            .in1(N__60850),
            .in2(N__70186),
            .in3(N__73156),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_17_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_17_10_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i14_LC_17_10_5  (
            .in0(N__79587),
            .in1(N__74104),
            .in2(N__60408),
            .in3(N__70178),
            .lcout(data_in_frame_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1860_LC_17_10_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1860_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1860_LC_17_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1860_LC_17_10_6  (
            .in0(N__60834),
            .in1(N__60377),
            .in2(N__57488),
            .in3(N__51223),
            .lcout(\c0.n15_adj_4710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_17_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_17_10_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i27_LC_17_10_7  (
            .in0(N__79190),
            .in1(N__70174),
            .in2(N__76599),
            .in3(N__57483),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_17_11_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_17_11_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i24_LC_17_11_0  (
            .in0(N__76148),
            .in1(N__70149),
            .in2(N__64755),
            .in3(N__69117),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_17_11_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_17_11_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i56_LC_17_11_1  (
            .in0(N__68422),
            .in1(N__76149),
            .in2(_gnd_net_),
            .in3(N__64873),
            .lcout(data_in_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_17_11_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_17_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i48_LC_17_11_2  (
            .in0(N__57638),
            .in1(N__76153),
            .in2(_gnd_net_),
            .in3(N__69411),
            .lcout(data_in_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i80_LC_17_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i80_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i80_LC_17_11_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i80_LC_17_11_3  (
            .in0(N__76152),
            .in1(N__73658),
            .in2(N__55023),
            .in3(N__74021),
            .lcout(\c0.data_in_frame_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1218_LC_17_11_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1218_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1218_LC_17_11_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i6_4_lut_adj_1218_LC_17_11_4  (
            .in0(N__49238),
            .in1(N__49303),
            .in2(N__48684),
            .in3(N__48636),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1843_LC_17_11_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1843_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1843_LC_17_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1843_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__57637),
            .in2(_gnd_net_),
            .in3(N__48743),
            .lcout(\c0.n6_adj_4704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1914_LC_17_11_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1914_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1914_LC_17_11_7 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \c0.i3_4_lut_adj_1914_LC_17_11_7  (
            .in0(N__51159),
            .in1(N__57782),
            .in2(N__51015),
            .in3(N__64377),
            .lcout(\c0.n20_adj_4729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_17_12_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_17_12_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i47_LC_17_12_0  (
            .in0(N__48739),
            .in1(N__69410),
            .in2(_gnd_net_),
            .in3(N__73201),
            .lcout(data_in_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78720),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1844_LC_17_12_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1844_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1844_LC_17_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1844_LC_17_12_1  (
            .in0(N__51574),
            .in1(N__58199),
            .in2(N__48588),
            .in3(N__60535),
            .lcout(\c0.n14016 ),
            .ltout(\c0.n14016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_1640_LC_17_12_2 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_1640_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_1640_LC_17_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i3_3_lut_adj_1640_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__61552),
            .in2(N__48579),
            .in3(N__55455),
            .lcout(\c0.n13329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_1826_LC_17_12_4 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_1826_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_1826_LC_17_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i6_2_lut_adj_1826_LC_17_12_4  (
            .in0(N__60534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48731),
            .lcout(\c0.n20 ),
            .ltout(\c0.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1347_LC_17_12_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1347_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1347_LC_17_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1347_LC_17_12_5  (
            .in0(N__55512),
            .in1(N__57636),
            .in2(N__48576),
            .in3(N__48697),
            .lcout(\c0.n4_adj_4333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_LC_17_12_6 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_17_12_6 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_17_12_6  (
            .in0(N__60536),
            .in1(N__48732),
            .in2(N__71187),
            .in3(N__55513),
            .lcout(\c0.n23_adj_4590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i114_LC_17_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i114_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i114_LC_17_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i114_LC_17_12_7  (
            .in0(N__75255),
            .in1(N__59207),
            .in2(_gnd_net_),
            .in3(N__55429),
            .lcout(data_in_frame_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78720),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i62_LC_17_13_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i62_LC_17_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i62_LC_17_13_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i62_LC_17_13_0  (
            .in0(N__79626),
            .in1(N__70147),
            .in2(N__64450),
            .in3(N__80920),
            .lcout(\c0.data_in_frame_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1717_LC_17_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1717_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1717_LC_17_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1717_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__65184),
            .in2(_gnd_net_),
            .in3(N__65073),
            .lcout(\c0.n5_adj_4443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i55_3_lut_4_lut_LC_17_13_2 .C_ON=1'b0;
    defparam \c0.i55_3_lut_4_lut_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i55_3_lut_4_lut_LC_17_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i55_3_lut_4_lut_LC_17_13_2  (
            .in0(N__62614),
            .in1(N__59259),
            .in2(N__61987),
            .in3(N__51275),
            .lcout(\c0.n136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i128_LC_17_13_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i128_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i128_LC_17_13_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i128_LC_17_13_3  (
            .in0(N__80919),
            .in1(N__73669),
            .in2(N__61991),
            .in3(N__76151),
            .lcout(\c0.data_in_frame_15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i101_LC_17_13_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i101_LC_17_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i101_LC_17_13_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i101_LC_17_13_4  (
            .in0(N__73668),
            .in1(N__59010),
            .in2(N__80099),
            .in3(N__71762),
            .lcout(\c0.data_in_frame_12_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i113_LC_17_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i113_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i113_LC_17_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i113_LC_17_13_5  (
            .in0(N__80575),
            .in1(N__59206),
            .in2(_gnd_net_),
            .in3(N__58614),
            .lcout(data_in_frame_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i64_LC_17_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i64_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i64_LC_17_13_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i64_LC_17_13_6  (
            .in0(N__76150),
            .in1(N__70148),
            .in2(N__48711),
            .in3(N__80921),
            .lcout(\c0.data_in_frame_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_17_13_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_17_13_7 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_17_13_7  (
            .in0(N__71761),
            .in1(N__49572),
            .in2(N__50904),
            .in3(N__49385),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i7_LC_17_14_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_17_14_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_17_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__49186),
            .in2(_gnd_net_),
            .in3(N__49007),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78697),
            .ce(),
            .sr(N__49170));
    defparam \c0.i6_4_lut_adj_1597_LC_17_14_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1597_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1597_LC_17_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1597_LC_17_14_2  (
            .in0(N__57663),
            .in1(N__61553),
            .in2(N__59011),
            .in3(N__58892),
            .lcout(\c0.n16_adj_4608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1202_LC_17_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1202_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1202_LC_17_14_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1202_LC_17_14_3  (
            .in0(N__55727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59001),
            .lcout(\c0.n13186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1901_LC_17_14_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1901_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1901_LC_17_14_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i8_4_lut_adj_1901_LC_17_14_4  (
            .in0(N__64884),
            .in1(N__57816),
            .in2(N__57671),
            .in3(N__64638),
            .lcout(\c0.n25_adj_4723 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_LC_17_14_5 .C_ON=1'b0;
    defparam \c0.i8_2_lut_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_LC_17_14_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i8_2_lut_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__64883),
            .in2(_gnd_net_),
            .in3(N__68127),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1900_LC_17_14_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1900_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1900_LC_17_14_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_adj_1900_LC_17_14_7  (
            .in0(N__64834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64737),
            .lcout(\c0.n7_adj_4337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1973_LC_17_15_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1973_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1973_LC_17_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1973_LC_17_15_0  (
            .in0(N__49143),
            .in1(N__49107),
            .in2(N__49083),
            .in3(N__48766),
            .lcout(\c0.n22049 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i27_LC_17_15_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_17_15_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_17_15_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_17_15_1  (
            .in0(N__48767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49011),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78681),
            .ce(),
            .sr(N__48753));
    defparam \c0.i42_4_lut_LC_17_15_7 .C_ON=1'b0;
    defparam \c0.i42_4_lut_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i42_4_lut_LC_17_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i42_4_lut_LC_17_15_7  (
            .in0(N__72689),
            .in1(N__72154),
            .in2(N__58937),
            .in3(N__59105),
            .lcout(\c0.n123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_9_i3_2_lut_LC_17_16_0 .C_ON=1'b0;
    defparam \c0.select_367_Select_9_i3_2_lut_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_9_i3_2_lut_LC_17_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_9_i3_2_lut_LC_17_16_0  (
            .in0(N__71519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52776),
            .lcout(\c0.n3_adj_4418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1348_LC_17_16_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1348_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1348_LC_17_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1348_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__62445),
            .in2(_gnd_net_),
            .in3(N__65405),
            .lcout(\c0.n22463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_17_16_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_17_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i3_LC_17_16_4  (
            .in0(N__50480),
            .in1(N__49272),
            .in2(_gnd_net_),
            .in3(N__49237),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78667),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_1701_LC_17_16_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_1701_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_1701_LC_17_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_1701_LC_17_16_5  (
            .in0(N__62379),
            .in1(N__59018),
            .in2(_gnd_net_),
            .in3(N__58775),
            .lcout(\c0.n15_adj_4301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1919_LC_17_16_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1919_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1919_LC_17_16_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1919_LC_17_16_6  (
            .in0(N__51291),
            .in1(N__58618),
            .in2(N__70482),
            .in3(N__62854),
            .lcout(\c0.n10_adj_4732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1231_LC_17_16_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1231_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1231_LC_17_16_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1231_LC_17_16_7  (
            .in0(N__49320),
            .in1(N__65460),
            .in2(N__69669),
            .in3(N__51279),
            .lcout(\c0.n21491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1920_LC_17_17_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1920_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1920_LC_17_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1920_LC_17_17_1  (
            .in0(N__62931),
            .in1(N__64662),
            .in2(N__49215),
            .in3(N__68556),
            .lcout(),
            .ltout(\c0.n26_adj_4733_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1989_LC_17_17_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1989_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1989_LC_17_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1989_LC_17_17_2  (
            .in0(N__68883),
            .in1(N__65538),
            .in2(N__49206),
            .in3(N__68593),
            .lcout(\c0.n20409 ),
            .ltout(\c0.n20409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1232_LC_17_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1232_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1232_LC_17_17_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1232_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49203),
            .in3(N__63542),
            .lcout(\c0.n22716 ),
            .ltout(\c0.n22716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_2042_LC_17_17_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_2042_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_2042_LC_17_17_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_2042_LC_17_17_4  (
            .in0(N__51773),
            .in1(N__56139),
            .in2(N__49323),
            .in3(N__59742),
            .lcout(\c0.n21389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1542_LC_17_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1542_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1542_LC_17_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1542_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__56193),
            .in2(_gnd_net_),
            .in3(N__58833),
            .lcout(\c0.n6_adj_4577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_17_17_7 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_17_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_17_17_7  (
            .in0(N__58619),
            .in1(N__66228),
            .in2(_gnd_net_),
            .in3(N__60063),
            .lcout(\c0.n8_adj_4248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_17_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_17_18_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i26_LC_17_18_0  (
            .in0(N__75028),
            .in1(N__50473),
            .in2(_gnd_net_),
            .in3(N__49302),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i171_LC_17_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i171_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i171_LC_17_18_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i171_LC_17_18_1  (
            .in0(N__78978),
            .in1(N__67620),
            .in2(_gnd_net_),
            .in3(N__51729),
            .lcout(data_in_frame_21_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1952_LC_17_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1952_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1952_LC_17_18_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1952_LC_17_18_2  (
            .in0(N__52480),
            .in1(N__52410),
            .in2(_gnd_net_),
            .in3(N__52568),
            .lcout(\c0.n12989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i148_LC_17_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i148_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i148_LC_17_18_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i148_LC_17_18_3  (
            .in0(N__80318),
            .in1(N__77102),
            .in2(N__69225),
            .in3(N__66650),
            .lcout(\c0.data_in_frame_18_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i172_LC_17_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i172_LC_17_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i172_LC_17_18_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i172_LC_17_18_4  (
            .in0(N__67621),
            .in1(N__77101),
            .in2(_gnd_net_),
            .in3(N__65884),
            .lcout(data_in_frame_21_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_14_i3_2_lut_LC_17_18_5 .C_ON=1'b0;
    defparam \c0.select_367_Select_14_i3_2_lut_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_14_i3_2_lut_LC_17_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_14_i3_2_lut_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__52955),
            .in2(_gnd_net_),
            .in3(N__71482),
            .lcout(\c0.n3_adj_4408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i168_LC_17_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i168_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i168_LC_17_18_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i168_LC_17_18_6  (
            .in0(N__80096),
            .in1(N__76389),
            .in2(N__56370),
            .in3(N__80319),
            .lcout(\c0.data_in_frame_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78668),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_16_i3_2_lut_LC_17_18_7 .C_ON=1'b0;
    defparam \c0.select_367_Select_16_i3_2_lut_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_16_i3_2_lut_LC_17_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_16_i3_2_lut_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__53054),
            .in2(_gnd_net_),
            .in3(N__71483),
            .lcout(\c0.n3_adj_4404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1642_LC_17_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1642_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1642_LC_17_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1642_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__72219),
            .in2(_gnd_net_),
            .in3(N__72161),
            .lcout(\c0.n13756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1478_LC_17_19_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1478_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1478_LC_17_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1478_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__59876),
            .in2(_gnd_net_),
            .in3(N__56515),
            .lcout(\c0.n15_adj_4508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_17_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_17_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i25_LC_17_19_2  (
            .in0(N__50484),
            .in1(N__80508),
            .in2(_gnd_net_),
            .in3(N__49422),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78682),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1536_LC_17_19_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1536_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1536_LC_17_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1536_LC_17_19_3  (
            .in0(N__58689),
            .in1(N__66579),
            .in2(N__61962),
            .in3(N__66369),
            .lcout(\c0.n23718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1365_LC_17_19_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1365_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1365_LC_17_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i2_2_lut_adj_1365_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__56354),
            .in2(_gnd_net_),
            .in3(N__63560),
            .lcout(\c0.n15_adj_4344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1390_LC_17_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1390_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1390_LC_17_19_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1390_LC_17_19_5  (
            .in0(N__56815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77273),
            .lcout(\c0.n5_adj_4370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_17_19_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_17_19_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_17_19_6  (
            .in0(N__49349),
            .in1(N__80509),
            .in2(N__50911),
            .in3(N__49378),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78682),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_17_19_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_17_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_17_19_7 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_17_19_7  (
            .in0(N__75027),
            .in1(N__49350),
            .in2(N__50910),
            .in3(N__50719),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78682),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1401_LC_17_20_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1401_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1401_LC_17_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1401_LC_17_20_0  (
            .in0(N__49332),
            .in1(N__66654),
            .in2(N__62982),
            .in3(N__56736),
            .lcout(\c0.n20_adj_4441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1541_LC_17_20_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1541_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1541_LC_17_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1541_LC_17_20_2  (
            .in0(N__51810),
            .in1(N__49473),
            .in2(N__52097),
            .in3(N__56738),
            .lcout(\c0.n14_adj_4576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1369_LC_17_20_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1369_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1369_LC_17_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1369_LC_17_20_3  (
            .in0(N__51777),
            .in1(N__59493),
            .in2(N__49494),
            .in3(N__61934),
            .lcout(),
            .ltout(\c0.n12_adj_4348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1486_LC_17_20_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1486_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1486_LC_17_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1486_LC_17_20_4  (
            .in0(N__66897),
            .in1(N__63306),
            .in2(N__49476),
            .in3(N__66710),
            .lcout(\c0.n8_adj_4526 ),
            .ltout(\c0.n8_adj_4526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1489_LC_17_20_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1489_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1489_LC_17_20_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1489_LC_17_20_5  (
            .in0(N__56737),
            .in1(N__52205),
            .in2(N__49467),
            .in3(N__51809),
            .lcout(\c0.n14_adj_4528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1496_LC_17_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1496_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1496_LC_17_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1496_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__76828),
            .in2(_gnd_net_),
            .in3(N__63241),
            .lcout(\c0.n9_adj_4536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1498_LC_17_21_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1498_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1498_LC_17_21_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1498_LC_17_21_0  (
            .in0(N__56276),
            .in1(N__49464),
            .in2(N__59875),
            .in3(N__49458),
            .lcout(\c0.n24547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1550_LC_17_21_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1550_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1550_LC_17_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1550_LC_17_21_1  (
            .in0(N__51870),
            .in1(N__51945),
            .in2(N__56649),
            .in3(N__49452),
            .lcout(\c0.n24098 ),
            .ltout(\c0.n24098_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1446_LC_17_21_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1446_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1446_LC_17_21_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1446_LC_17_21_2  (
            .in0(N__49445),
            .in1(N__52035),
            .in2(N__49434),
            .in3(N__51897),
            .lcout(\c0.n10_adj_4484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_adj_1736_LC_17_21_4 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_adj_1736_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_adj_1736_LC_17_21_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_3_lut_4_lut_adj_1736_LC_17_21_4  (
            .in0(N__77291),
            .in1(N__76833),
            .in2(N__59628),
            .in3(N__56752),
            .lcout(\c0.n20_adj_4512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i170_LC_17_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i170_LC_17_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i170_LC_17_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i170_LC_17_21_6  (
            .in0(N__66426),
            .in1(N__75113),
            .in2(_gnd_net_),
            .in3(N__67644),
            .lcout(data_in_frame_21_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78711),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1370_LC_17_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1370_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1370_LC_17_21_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1370_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__66425),
            .in2(_gnd_net_),
            .in3(N__51778),
            .lcout(\c0.n5_adj_4349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1435_LC_17_22_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1435_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1435_LC_17_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1435_LC_17_22_0  (
            .in0(N__56670),
            .in1(N__49500),
            .in2(N__49523),
            .in3(N__59524),
            .lcout(),
            .ltout(\c0.n52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_adj_1500_LC_17_22_1 .C_ON=1'b0;
    defparam \c0.i30_4_lut_adj_1500_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_adj_1500_LC_17_22_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i30_4_lut_adj_1500_LC_17_22_1  (
            .in0(N__59557),
            .in1(N__72371),
            .in2(N__49539),
            .in3(N__67038),
            .lcout(\c0.n64_adj_4539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_1513_LC_17_22_2 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_1513_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_1513_LC_17_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_1513_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__59556),
            .in2(_gnd_net_),
            .in3(N__59525),
            .lcout(),
            .ltout(\c0.n47_adj_4537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1497_LC_17_22_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1497_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1497_LC_17_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1497_LC_17_22_3  (
            .in0(N__57076),
            .in1(N__49508),
            .in2(N__49536),
            .in3(N__56893),
            .lcout(\c0.n24581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i234_LC_17_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i234_LC_17_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i234_LC_17_22_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i234_LC_17_22_4  (
            .in0(N__75112),
            .in1(N__56461),
            .in2(N__49524),
            .in3(N__75407),
            .lcout(\c0.data_in_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i239_LC_17_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i239_LC_17_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i239_LC_17_22_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i239_LC_17_22_5  (
            .in0(N__75406),
            .in1(N__73346),
            .in2(N__56479),
            .in3(N__49509),
            .lcout(\c0.data_in_frame_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1704_LC_17_22_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1704_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1704_LC_17_22_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1704_LC_17_22_6  (
            .in0(N__67121),
            .in1(N__52028),
            .in2(N__57021),
            .in3(N__51998),
            .lcout(\c0.n20793 ),
            .ltout(\c0.n20793_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_LC_17_22_7 .C_ON=1'b0;
    defparam \c0.i28_4_lut_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_LC_17_22_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i28_4_lut_LC_17_22_7  (
            .in0(N__63018),
            .in1(N__59912),
            .in2(N__49557),
            .in3(N__72370),
            .lcout(\c0.n70_adj_4514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_4_lut_LC_17_23_0 .C_ON=1'b0;
    defparam \c0.i4_2_lut_4_lut_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_4_lut_LC_17_23_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_2_lut_4_lut_LC_17_23_0  (
            .in0(N__66430),
            .in1(N__56369),
            .in2(N__56411),
            .in3(N__51779),
            .lcout(\c0.n14_adj_4529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i216_LC_17_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i216_LC_17_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i216_LC_17_23_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i216_LC_17_23_2  (
            .in0(N__79362),
            .in1(N__69224),
            .in2(N__76365),
            .in3(N__67296),
            .lcout(\c0.data_in_frame_26_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i167_LC_17_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i167_LC_17_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i167_LC_17_23_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i167_LC_17_23_4  (
            .in0(N__73298),
            .in1(N__56406),
            .in2(N__80100),
            .in3(N__80424),
            .lcout(\c0.data_in_frame_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1277_LC_17_23_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1277_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1277_LC_17_23_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1277_LC_17_23_5  (
            .in0(N__62316),
            .in1(N__52407),
            .in2(_gnd_net_),
            .in3(N__49844),
            .lcout(\c0.n12927 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i211_LC_17_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i211_LC_17_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i211_LC_17_23_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i211_LC_17_23_7  (
            .in0(N__69223),
            .in1(N__79173),
            .in2(N__66807),
            .in3(N__79363),
            .lcout(\c0.data_in_frame_26_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_15_i3_2_lut_LC_17_24_0 .C_ON=1'b0;
    defparam \c0.select_367_Select_15_i3_2_lut_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_15_i3_2_lut_LC_17_24_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_15_i3_2_lut_LC_17_24_0  (
            .in0(N__71348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53006),
            .lcout(\c0.n3_adj_4406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_11_i3_2_lut_LC_17_24_1 .C_ON=1'b0;
    defparam \c0.select_367_Select_11_i3_2_lut_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_11_i3_2_lut_LC_17_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_11_i3_2_lut_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__52836),
            .in2(_gnd_net_),
            .in3(N__71347),
            .lcout(\c0.n3_adj_4414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_6_i3_2_lut_LC_17_24_2 .C_ON=1'b0;
    defparam \c0.select_367_Select_6_i3_2_lut_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_6_i3_2_lut_LC_17_24_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_6_i3_2_lut_LC_17_24_2  (
            .in0(N__71351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52575),
            .lcout(\c0.n3_adj_4424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i204_LC_17_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i204_LC_17_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i204_LC_17_24_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i204_LC_17_24_3  (
            .in0(N__74216),
            .in1(N__76945),
            .in2(N__52204),
            .in3(N__79421),
            .lcout(\c0.data_in_frame_25_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_23_i3_2_lut_LC_17_24_4 .C_ON=1'b0;
    defparam \c0.select_367_Select_23_i3_2_lut_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_23_i3_2_lut_LC_17_24_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_23_i3_2_lut_LC_17_24_4  (
            .in0(N__71350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53309),
            .lcout(\c0.n3_adj_4390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_22_i3_2_lut_LC_17_24_7 .C_ON=1'b0;
    defparam \c0.select_367_Select_22_i3_2_lut_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_22_i3_2_lut_LC_17_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_22_i3_2_lut_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__53271),
            .in2(_gnd_net_),
            .in3(N__71349),
            .lcout(\c0.n3_adj_4392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_24_i3_2_lut_LC_17_25_0 .C_ON=1'b0;
    defparam \c0.select_367_Select_24_i3_2_lut_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_24_i3_2_lut_LC_17_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_24_i3_2_lut_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__53346),
            .in2(_gnd_net_),
            .in3(N__71372),
            .lcout(\c0.n3_adj_4388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1953_LC_17_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1953_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1953_LC_17_25_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1953_LC_17_25_1  (
            .in0(N__52409),
            .in1(N__52485),
            .in2(_gnd_net_),
            .in3(N__52561),
            .lcout(\c0.n12973 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_1276_LC_17_25_7 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_1276_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_1276_LC_17_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i25_4_lut_adj_1276_LC_17_25_7  (
            .in0(N__49857),
            .in1(N__52140),
            .in2(N__52215),
            .in3(N__52257),
            .lcout(\c0.n13043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1267_LC_17_26_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1267_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1267_LC_17_26_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_1267_LC_17_26_1  (
            .in0(N__53409),
            .in1(N__52835),
            .in2(N__53058),
            .in3(N__53270),
            .lcout(\c0.n41_adj_4292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19124_2_lut_3_lut_LC_17_27_6 .C_ON=1'b0;
    defparam \c0.i19124_2_lut_3_lut_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i19124_2_lut_3_lut_LC_17_27_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.i19124_2_lut_3_lut_LC_17_27_6  (
            .in0(N__53908),
            .in1(N__49830),
            .in2(_gnd_net_),
            .in3(N__49787),
            .lcout(\c0.n22885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_31_i3_2_lut_LC_17_32_4 .C_ON=1'b0;
    defparam \c0.select_367_Select_31_i3_2_lut_LC_17_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_31_i3_2_lut_LC_17_32_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_31_i3_2_lut_LC_17_32_4  (
            .in0(_gnd_net_),
            .in1(N__53881),
            .in2(_gnd_net_),
            .in3(N__71536),
            .lcout(\c0.n3_adj_4373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_102_i4_2_lut_LC_18_1_0 .C_ON=1'b0;
    defparam \c0.rx.equal_102_i4_2_lut_LC_18_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_102_i4_2_lut_LC_18_1_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.equal_102_i4_2_lut_LC_18_1_0  (
            .in0(_gnd_net_),
            .in1(N__49740),
            .in2(_gnd_net_),
            .in3(N__49662),
            .lcout(n4),
            .ltout(n4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_18_1_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_18_1_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_18_1_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_18_1_1  (
            .in0(N__79542),
            .in1(N__50909),
            .in2(N__50736),
            .in3(N__50733),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78822),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_18_1_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_18_1_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_18_1_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_18_1_2  (
            .in0(N__50234),
            .in1(N__49943),
            .in2(N__50184),
            .in3(N__50679),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78822),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_LC_18_1_3 .C_ON=1'b0;
    defparam \c0.i14_2_lut_LC_18_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_LC_18_1_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i14_2_lut_LC_18_1_3  (
            .in0(_gnd_net_),
            .in1(N__50198),
            .in2(_gnd_net_),
            .in3(N__50233),
            .lcout(\c0.n161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1887_LC_18_1_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1887_LC_18_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1887_LC_18_1_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1887_LC_18_1_4  (
            .in0(N__50664),
            .in1(N__50634),
            .in2(N__50598),
            .in3(N__50541),
            .lcout(\c0.n21_adj_4719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_18_1_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_18_1_5 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_18_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_18_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50235),
            .lcout(\c0.FRAME_MATCHER_rx_data_ready_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78822),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21281_2_lut_3_lut_LC_18_1_6 .C_ON=1'b0;
    defparam \c0.rx.i21281_2_lut_3_lut_LC_18_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21281_2_lut_3_lut_LC_18_1_6 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.rx.i21281_2_lut_3_lut_LC_18_1_6  (
            .in0(N__50179),
            .in1(N__50055),
            .in2(_gnd_net_),
            .in3(N__49942),
            .lcout(\c0.rx.n22094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_1940_LC_18_6_0 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_1940_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_1940_LC_18_6_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.i22_4_lut_adj_1940_LC_18_6_0  (
            .in0(N__50994),
            .in1(N__51000),
            .in2(N__59949),
            .in3(N__60327),
            .lcout(\c0.n46_adj_4739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_99_i9_2_lut_3_lut_LC_18_6_2 .C_ON=1'b0;
    defparam \c0.equal_99_i9_2_lut_3_lut_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.equal_99_i9_2_lut_3_lut_LC_18_6_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.equal_99_i9_2_lut_3_lut_LC_18_6_2  (
            .in0(N__74625),
            .in1(N__74288),
            .in2(_gnd_net_),
            .in3(N__74499),
            .lcout(\c0.n9_adj_4563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_5_i3_2_lut_LC_18_6_7 .C_ON=1'b0;
    defparam \c0.select_367_Select_5_i3_2_lut_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_5_i3_2_lut_LC_18_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_5_i3_2_lut_LC_18_6_7  (
            .in0(_gnd_net_),
            .in1(N__52455),
            .in2(_gnd_net_),
            .in3(N__71545),
            .lcout(\c0.n3_adj_4426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i59_LC_18_7_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i59_LC_18_7_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i59_LC_18_7_1 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i59_LC_18_7_1  (
            .in0(N__80871),
            .in1(N__70173),
            .in2(N__70741),
            .in3(N__79107),
            .lcout(\c0.data_in_frame_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78786),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1933_LC_18_7_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1933_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1933_LC_18_7_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.i15_4_lut_adj_1933_LC_18_7_3  (
            .in0(N__64272),
            .in1(N__71032),
            .in2(N__68555),
            .in3(N__51219),
            .lcout(\c0.n39_adj_4737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1932_LC_18_7_4 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1932_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1932_LC_18_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14_4_lut_adj_1932_LC_18_7_4  (
            .in0(N__57243),
            .in1(N__51460),
            .in2(N__61064),
            .in3(N__58043),
            .lcout(\c0.n38_adj_4736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1663_LC_18_8_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1663_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1663_LC_18_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1663_LC_18_8_0  (
            .in0(N__60229),
            .in1(N__51424),
            .in2(_gnd_net_),
            .in3(N__51216),
            .lcout(\c0.n4_adj_4267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_LC_18_8_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_LC_18_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_LC_18_8_1  (
            .in0(N__51217),
            .in1(N__57930),
            .in2(N__51447),
            .in3(N__60230),
            .lcout(\c0.n23562 ),
            .ltout(\c0.n23562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_LC_18_8_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_LC_18_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_LC_18_8_2  (
            .in0(N__50941),
            .in1(_gnd_net_),
            .in2(N__50976),
            .in3(N__50973),
            .lcout(\c0.n13280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_adj_1837_LC_18_8_3 .C_ON=1'b0;
    defparam \c0.i13_2_lut_adj_1837_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_adj_1837_LC_18_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i13_2_lut_adj_1837_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(N__55322),
            .in2(_gnd_net_),
            .in3(N__57235),
            .lcout(\c0.n22_adj_4647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_18_8_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_18_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_18_8_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i28_LC_18_8_4  (
            .in0(N__77065),
            .in1(N__76595),
            .in2(N__57949),
            .in3(N__70169),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1851_LC_18_8_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1851_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1851_LC_18_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1851_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__50940),
            .in2(_gnd_net_),
            .in3(N__57234),
            .lcout(\c0.n22511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1722_LC_18_8_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1722_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1722_LC_18_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1722_LC_18_8_6  (
            .in0(N__57236),
            .in1(N__57507),
            .in2(N__60239),
            .in3(N__51021),
            .lcout(\c0.n13141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_18_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_18_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_18_8_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i16_LC_18_8_7  (
            .in0(N__70168),
            .in1(N__74145),
            .in2(N__71078),
            .in3(N__76285),
            .lcout(data_in_frame_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_4_lut_LC_18_9_0 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_4_lut_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_4_lut_LC_18_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_2_lut_3_lut_4_lut_LC_18_9_0  (
            .in0(N__55332),
            .in1(N__51420),
            .in2(N__57535),
            .in3(N__51218),
            .lcout(\c0.n18_adj_4228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_3_lut_4_lut_LC_18_9_1 .C_ON=1'b0;
    defparam \c0.i10_3_lut_4_lut_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_3_lut_4_lut_LC_18_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_3_lut_4_lut_LC_18_9_1  (
            .in0(N__71031),
            .in1(N__56013),
            .in2(N__60545),
            .in3(N__51136),
            .lcout(\c0.n23_adj_4648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_3_lut_4_lut_LC_18_9_2 .C_ON=1'b0;
    defparam \c0.i27_3_lut_4_lut_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i27_3_lut_4_lut_LC_18_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_3_lut_4_lut_LC_18_9_2  (
            .in0(N__60387),
            .in1(N__71030),
            .in2(N__72414),
            .in3(N__58014),
            .lcout(\c0.n63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_1593_LC_18_9_3 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_1593_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_1593_LC_18_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_1593_LC_18_9_3  (
            .in0(N__55124),
            .in1(N__51613),
            .in2(_gnd_net_),
            .in3(N__55980),
            .lcout(\c0.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1853_LC_18_9_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1853_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1853_LC_18_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1853_LC_18_9_4  (
            .in0(N__51563),
            .in1(N__60507),
            .in2(_gnd_net_),
            .in3(N__51419),
            .lcout(\c0.n22160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_18_9_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_18_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_18_9_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i12_LC_18_9_7  (
            .in0(N__77129),
            .in1(N__74179),
            .in2(N__51446),
            .in3(N__70179),
            .lcout(data_in_frame_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78771),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_LC_18_10_0 .C_ON=1'b0;
    defparam \c0.i9_2_lut_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_LC_18_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i9_2_lut_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__60511),
            .in2(_gnd_net_),
            .in3(N__60385),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_18_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_18_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_18_10_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i15_LC_18_10_2  (
            .in0(N__70138),
            .in1(N__74068),
            .in2(N__58055),
            .in3(N__73349),
            .lcout(data_in_frame_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_18_10_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_18_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_18_10_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i13_LC_18_10_3  (
            .in0(N__71915),
            .in1(N__74051),
            .in2(N__60546),
            .in3(N__70140),
            .lcout(data_in_frame_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_1993_LC_18_10_4 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_1993_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_1993_LC_18_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_1993_LC_18_10_4  (
            .in0(N__69728),
            .in1(N__61263),
            .in2(N__71220),
            .in3(N__71077),
            .lcout(\c0.n44_adj_4744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i63_LC_18_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i63_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i63_LC_18_10_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i63_LC_18_10_5  (
            .in0(N__73348),
            .in1(N__70139),
            .in2(N__57308),
            .in3(N__80888),
            .lcout(\c0.data_in_frame_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1666_LC_18_10_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1666_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1666_LC_18_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1666_LC_18_10_6  (
            .in0(N__68545),
            .in1(N__68126),
            .in2(N__67944),
            .in3(N__51044),
            .lcout(\c0.n13_adj_4584 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i117_LC_18_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i117_LC_18_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i117_LC_18_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i117_LC_18_10_7  (
            .in0(N__71914),
            .in1(N__59208),
            .in2(_gnd_net_),
            .in3(N__55919),
            .lcout(data_in_frame_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1263_LC_18_11_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1263_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1263_LC_18_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1263_LC_18_11_0  (
            .in0(N__51150),
            .in1(N__51117),
            .in2(N__55383),
            .in3(N__61302),
            .lcout(),
            .ltout(\c0.n38_adj_4285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_18_11_1 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_18_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_LC_18_11_1  (
            .in0(N__51030),
            .in1(N__51054),
            .in2(N__51057),
            .in3(N__70233),
            .lcout(\c0.n24527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_2_lut_3_lut_4_lut_adj_2029_LC_18_11_2 .C_ON=1'b0;
    defparam \c0.i11_2_lut_3_lut_4_lut_adj_2029_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_2_lut_3_lut_4_lut_adj_2029_LC_18_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_2_lut_3_lut_4_lut_adj_2029_LC_18_11_2  (
            .in0(N__51233),
            .in1(N__57563),
            .in2(N__51464),
            .in3(N__51138),
            .lcout(\c0.n26_adj_4289 ),
            .ltout(\c0.n26_adj_4289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_3_lut_4_lut_adj_1622_LC_18_11_3 .C_ON=1'b0;
    defparam \c0.i13_3_lut_4_lut_adj_1622_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_3_lut_4_lut_adj_1622_LC_18_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_3_lut_4_lut_adj_1622_LC_18_11_3  (
            .in0(N__51029),
            .in1(N__57721),
            .in2(N__51048),
            .in3(N__58169),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_2_lut_3_lut_LC_18_11_4 .C_ON=1'b0;
    defparam \c0.i11_2_lut_3_lut_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_2_lut_3_lut_LC_18_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i11_2_lut_3_lut_LC_18_11_4  (
            .in0(N__64839),
            .in1(N__64724),
            .in2(_gnd_net_),
            .in3(N__51045),
            .lcout(\c0.n20_adj_4290 ),
            .ltout(\c0.n20_adj_4290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_2_lut_3_lut_4_lut_adj_2026_LC_18_11_5 .C_ON=1'b0;
    defparam \c0.i21_2_lut_3_lut_4_lut_adj_2026_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21_2_lut_3_lut_4_lut_adj_2026_LC_18_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_2_lut_3_lut_4_lut_adj_2026_LC_18_11_5  (
            .in0(N__57562),
            .in1(N__51448),
            .in2(N__51240),
            .in3(N__51232),
            .lcout(\c0.n51 ),
            .ltout(\c0.n51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_3_lut_LC_18_11_6 .C_ON=1'b0;
    defparam \c0.i26_3_lut_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i26_3_lut_LC_18_11_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i26_3_lut_LC_18_11_6  (
            .in0(N__51149),
            .in1(_gnd_net_),
            .in2(N__51141),
            .in3(N__51137),
            .lcout(\c0.n56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_2_lut_3_lut_4_lut_LC_18_12_0 .C_ON=1'b0;
    defparam \c0.i21_2_lut_3_lut_4_lut_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21_2_lut_3_lut_4_lut_LC_18_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_2_lut_3_lut_4_lut_LC_18_12_0  (
            .in0(N__57381),
            .in1(N__55221),
            .in2(N__51108),
            .in3(N__64677),
            .lcout(\c0.n102 ),
            .ltout(\c0.n102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_adj_1261_LC_18_12_1 .C_ON=1'b0;
    defparam \c0.i12_3_lut_adj_1261_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_adj_1261_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i12_3_lut_adj_1261_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__55430),
            .in2(N__51120),
            .in3(N__64988),
            .lcout(\c0.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_LC_18_12_2 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_LC_18_12_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i4_2_lut_3_lut_LC_18_12_2  (
            .in0(N__70551),
            .in1(N__58751),
            .in2(_gnd_net_),
            .in3(N__58967),
            .lcout(\c0.n16_adj_4256 ),
            .ltout(\c0.n16_adj_4256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i45_4_lut_LC_18_12_3 .C_ON=1'b0;
    defparam \c0.i45_4_lut_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i45_4_lut_LC_18_12_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i45_4_lut_LC_18_12_3  (
            .in0(N__51063),
            .in1(N__54984),
            .in2(N__51111),
            .in3(N__69800),
            .lcout(\c0.n126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_1646_LC_18_12_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_1646_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_1646_LC_18_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3_2_lut_adj_1646_LC_18_12_4  (
            .in0(N__55185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64733),
            .lcout(\c0.n9_adj_4279 ),
            .ltout(\c0.n9_adj_4279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_18_12_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_18_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_18_12_5  (
            .in0(N__51092),
            .in1(N__55242),
            .in2(N__51069),
            .in3(N__64440),
            .lcout(\c0.n23574 ),
            .ltout(\c0.n23574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_LC_18_12_6 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_LC_18_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_3_lut_4_lut_LC_18_12_6  (
            .in0(N__55186),
            .in1(N__70352),
            .in2(N__51066),
            .in3(N__64606),
            .lcout(\c0.n11_adj_4257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1995_LC_18_13_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1995_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1995_LC_18_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1995_LC_18_13_0  (
            .in0(N__69898),
            .in1(N__60159),
            .in2(N__64239),
            .in3(N__64017),
            .lcout(\c0.n41_adj_4745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_adj_2045_LC_18_13_1 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_adj_2045_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_adj_2045_LC_18_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_3_lut_4_lut_adj_2045_LC_18_13_1  (
            .in0(N__70353),
            .in1(N__51328),
            .in2(N__69902),
            .in3(N__57537),
            .lcout(\c0.n38_adj_4573 ),
            .ltout(\c0.n38_adj_4573_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_3_lut_4_lut_LC_18_13_2 .C_ON=1'b0;
    defparam \c0.i19_3_lut_4_lut_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i19_3_lut_4_lut_LC_18_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_3_lut_4_lut_LC_18_13_2  (
            .in0(N__58419),
            .in1(N__64347),
            .in2(N__51312),
            .in3(N__70298),
            .lcout(),
            .ltout(\c0.n43_adj_4574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_adj_2009_LC_18_13_3 .C_ON=1'b0;
    defparam \c0.i23_4_lut_adj_2009_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_adj_2009_LC_18_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_adj_2009_LC_18_13_3  (
            .in0(N__51309),
            .in1(N__67998),
            .in2(N__51300),
            .in3(N__51297),
            .lcout(\c0.n24048 ),
            .ltout(\c0.n24048_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_3_lut_LC_18_13_4 .C_ON=1'b0;
    defparam \c0.i28_3_lut_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i28_3_lut_LC_18_13_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i28_3_lut_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__65964),
            .in2(N__51282),
            .in3(N__56043),
            .lcout(\c0.n109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_18_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_18_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_18_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i53_LC_18_13_5  (
            .in0(N__71816),
            .in1(N__68441),
            .in2(_gnd_net_),
            .in3(N__65193),
            .lcout(data_in_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1923_LC_18_14_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1923_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1923_LC_18_14_0 .LUT_INIT=16'b1111011111111101;
    LogicCell40 \c0.i12_4_lut_adj_1923_LC_18_14_0  (
            .in0(N__64613),
            .in1(N__57579),
            .in2(N__51264),
            .in3(N__58373),
            .lcout(\c0.n29_adj_4734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1829_LC_18_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1829_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1829_LC_18_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1829_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__55125),
            .in2(_gnd_net_),
            .in3(N__55976),
            .lcout(\c0.n7_adj_4221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i35_LC_18_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i35_LC_18_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i35_LC_18_14_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i35_LC_18_14_2  (
            .in0(N__79203),
            .in1(N__70078),
            .in2(N__80098),
            .in3(N__65069),
            .lcout(\c0.data_in_frame_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1653_LC_18_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1653_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1653_LC_18_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1653_LC_18_14_3  (
            .in0(N__58137),
            .in1(N__64409),
            .in2(_gnd_net_),
            .in3(N__58080),
            .lcout(\c0.n16_adj_4641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_18_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_18_14_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i32_LC_18_14_4  (
            .in0(N__76315),
            .in1(N__76612),
            .in2(N__58090),
            .in3(N__70079),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1651_LC_18_14_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1651_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1651_LC_18_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1651_LC_18_14_5  (
            .in0(N__65068),
            .in1(N__58079),
            .in2(_gnd_net_),
            .in3(N__55798),
            .lcout(\c0.n23313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i34_LC_18_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i34_LC_18_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i34_LC_18_14_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i34_LC_18_14_6  (
            .in0(N__55800),
            .in1(N__75256),
            .in2(N__80097),
            .in3(N__70080),
            .lcout(\c0.data_in_frame_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1854_LC_18_14_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1854_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1854_LC_18_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1854_LC_18_14_7  (
            .in0(N__54951),
            .in1(N__58078),
            .in2(_gnd_net_),
            .in3(N__55799),
            .lcout(\c0.n14_adj_4707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1195_LC_18_15_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1195_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1195_LC_18_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1195_LC_18_15_0  (
            .in0(N__51467),
            .in1(N__51354),
            .in2(N__55905),
            .in3(N__51521),
            .lcout(\c0.n20_adj_4222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_2_lut_3_lut_4_lut_LC_18_15_1 .C_ON=1'b0;
    defparam \c0.i22_2_lut_3_lut_4_lut_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i22_2_lut_3_lut_4_lut_LC_18_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_2_lut_3_lut_4_lut_LC_18_15_1  (
            .in0(N__60906),
            .in1(N__55901),
            .in2(N__51522),
            .in3(N__57731),
            .lcout(\c0.n58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1813_LC_18_15_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1813_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1813_LC_18_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1813_LC_18_15_2  (
            .in0(N__58372),
            .in1(N__57900),
            .in2(N__60562),
            .in3(N__51345),
            .lcout(\c0.n23116 ),
            .ltout(\c0.n23116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1827_LC_18_15_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1827_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1827_LC_18_15_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_1827_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51339),
            .in3(N__55899),
            .lcout(\c0.n11_adj_4614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i48_4_lut_LC_18_15_4 .C_ON=1'b0;
    defparam \c0.i48_4_lut_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i48_4_lut_LC_18_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i48_4_lut_LC_18_15_4  (
            .in0(N__55900),
            .in1(N__51517),
            .in2(N__58173),
            .in3(N__66173),
            .lcout(),
            .ltout(\c0.n129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i73_4_lut_LC_18_15_5 .C_ON=1'b0;
    defparam \c0.i73_4_lut_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i73_4_lut_LC_18_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i73_4_lut_LC_18_15_5  (
            .in0(N__51507),
            .in1(N__55644),
            .in2(N__51492),
            .in3(N__58242),
            .lcout(\c0.n154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1611_LC_18_15_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1611_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1611_LC_18_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1611_LC_18_15_6  (
            .in0(N__51581),
            .in1(N__60552),
            .in2(N__55682),
            .in3(N__62084),
            .lcout(),
            .ltout(\c0.n16_adj_4613_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1612_LC_18_15_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1612_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1612_LC_18_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1612_LC_18_15_7  (
            .in0(N__60905),
            .in1(N__51489),
            .in2(N__51483),
            .in3(N__51466),
            .lcout(\c0.n23390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_18_16_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_18_16_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_LC_18_16_0  (
            .in0(N__56085),
            .in1(N__55566),
            .in2(N__73861),
            .in3(N__65835),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1585_LC_18_16_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1585_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1585_LC_18_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1585_LC_18_16_1  (
            .in0(N__58544),
            .in1(N__58776),
            .in2(N__59243),
            .in3(N__56084),
            .lcout(\c0.n21_adj_4605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1584_LC_18_16_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1584_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1584_LC_18_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1584_LC_18_16_2  (
            .in0(N__61616),
            .in1(N__61658),
            .in2(N__72693),
            .in3(N__58890),
            .lcout(\c0.n19_adj_4604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i116_LC_18_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i116_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i116_LC_18_16_3 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \c0.data_in_frame_0__i116_LC_18_16_3  (
            .in0(N__76954),
            .in1(N__59197),
            .in2(N__55823),
            .in3(_gnd_net_),
            .lcout(data_in_frame_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78683),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i63_4_lut_LC_18_16_4 .C_ON=1'b0;
    defparam \c0.i63_4_lut_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i63_4_lut_LC_18_16_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i63_4_lut_LC_18_16_4  (
            .in0(N__51372),
            .in1(N__58891),
            .in2(N__51675),
            .in3(N__66160),
            .lcout(),
            .ltout(\c0.n144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i77_4_lut_LC_18_16_5 .C_ON=1'b0;
    defparam \c0.i77_4_lut_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i77_4_lut_LC_18_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i77_4_lut_LC_18_16_5  (
            .in0(N__62151),
            .in1(N__51363),
            .in2(N__51357),
            .in3(N__51681),
            .lcout(\c0.n158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i119_LC_18_16_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i119_LC_18_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i119_LC_18_16_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_frame_0__i119_LC_18_16_7  (
            .in0(N__59231),
            .in1(_gnd_net_),
            .in2(N__73356),
            .in3(N__59198),
            .lcout(data_in_frame_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78683),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1586_LC_18_17_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1586_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1586_LC_18_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1586_LC_18_17_0  (
            .in0(N__51671),
            .in1(N__51657),
            .in2(N__51651),
            .in3(N__51642),
            .lcout(\c0.n21344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1196_LC_18_17_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1196_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1196_LC_18_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1196_LC_18_17_1  (
            .in0(N__59300),
            .in1(N__51633),
            .in2(N__55275),
            .in3(N__55523),
            .lcout(),
            .ltout(\c0.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_18_17_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_18_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_18_17_2  (
            .in0(N__51626),
            .in1(N__55741),
            .in2(N__51597),
            .in3(N__51594),
            .lcout(),
            .ltout(\c0.n22_adj_4223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_18_17_3 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_18_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_18_17_3  (
            .in0(N__58263),
            .in1(N__51585),
            .in2(N__51531),
            .in3(N__60553),
            .lcout(\c0.n21_adj_4225 ),
            .ltout(\c0.n21_adj_4225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1257_LC_18_17_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1257_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1257_LC_18_17_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_1257_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51528),
            .in3(N__77654),
            .lcout(),
            .ltout(\c0.n10_adj_4277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1258_LC_18_17_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1258_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1258_LC_18_17_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1258_LC_18_17_5  (
            .in0(N__56163),
            .in1(N__66309),
            .in2(N__51525),
            .in3(N__77583),
            .lcout(\c0.n13_adj_4281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1587_LC_18_18_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1587_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1587_LC_18_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1587_LC_18_18_0  (
            .in0(N__61901),
            .in1(N__66570),
            .in2(N__63441),
            .in3(N__58871),
            .lcout(\c0.n10_adj_4591 ),
            .ltout(\c0.n10_adj_4591_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1565_LC_18_18_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1565_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1565_LC_18_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_1565_LC_18_18_1  (
            .in0(N__51727),
            .in1(N__73854),
            .in2(N__51738),
            .in3(N__62711),
            .lcout(\c0.n41_adj_4592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1589_LC_18_18_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1589_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1589_LC_18_18_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1589_LC_18_18_2  (
            .in0(N__62712),
            .in1(N__51735),
            .in2(N__73862),
            .in3(N__65846),
            .lcout(),
            .ltout(\c0.n12_adj_4606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1590_LC_18_18_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1590_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1590_LC_18_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1590_LC_18_18_3  (
            .in0(N__51728),
            .in1(N__59479),
            .in2(N__51714),
            .in3(N__63471),
            .lcout(\c0.n21325 ),
            .ltout(\c0.n21325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1559_LC_18_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1559_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1559_LC_18_18_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1559_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51711),
            .in3(N__76832),
            .lcout(\c0.n4_adj_4464 ),
            .ltout(\c0.n4_adj_4464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1460_LC_18_18_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1460_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1460_LC_18_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1460_LC_18_18_5  (
            .in0(N__51708),
            .in1(N__56268),
            .in2(N__51693),
            .in3(N__74733),
            .lcout(\c0.n12_adj_4506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i189_LC_18_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i189_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i189_LC_18_18_6 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.data_in_frame_0__i189_LC_18_18_6  (
            .in0(N__59480),
            .in1(N__71913),
            .in2(N__80982),
            .in3(N__80324),
            .lcout(\c0.data_in_frame_23_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1569_LC_18_19_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1569_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1569_LC_18_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1569_LC_18_19_0  (
            .in0(N__51687),
            .in1(N__51864),
            .in2(N__63089),
            .in3(N__59440),
            .lcout(\c0.n23863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1570_LC_18_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1570_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1570_LC_18_19_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1570_LC_18_19_1  (
            .in0(N__65853),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63381),
            .lcout(\c0.n21428 ),
            .ltout(\c0.n21428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1566_LC_18_19_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1566_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1566_LC_18_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_4_lut_adj_1566_LC_18_19_2  (
            .in0(N__51834),
            .in1(N__58527),
            .in2(N__51690),
            .in3(N__56323),
            .lcout(\c0.n24_adj_4593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_LC_18_19_3 .C_ON=1'b0;
    defparam \c0.i8_3_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_LC_18_19_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i8_3_lut_LC_18_19_3  (
            .in0(N__65854),
            .in1(N__66431),
            .in2(_gnd_net_),
            .in3(N__51843),
            .lcout(\c0.n23_adj_4598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1372_LC_18_19_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1372_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1372_LC_18_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1372_LC_18_19_4  (
            .in0(N__77688),
            .in1(N__58482),
            .in2(N__51858),
            .in3(N__58794),
            .lcout(\c0.n23_adj_4353 ),
            .ltout(\c0.n23_adj_4353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1393_LC_18_19_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1393_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1393_LC_18_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1393_LC_18_19_5  (
            .in0(N__72360),
            .in1(N__56427),
            .in2(N__51837),
            .in3(N__51833),
            .lcout(\c0.n16_adj_4437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1394_LC_18_19_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1394_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1394_LC_18_19_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_adj_1394_LC_18_19_6  (
            .in0(N__58523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56322),
            .lcout(),
            .ltout(\c0.n11_adj_4438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1395_LC_18_19_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1395_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1395_LC_18_19_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1395_LC_18_19_7  (
            .in0(N__59286),
            .in1(N__51825),
            .in2(N__51819),
            .in3(N__51816),
            .lcout(\c0.n21280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_18_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_18_20_0  (
            .in0(N__66987),
            .in1(N__57887),
            .in2(N__66900),
            .in3(N__59442),
            .lcout(\c0.n22420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1463_LC_18_20_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1463_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1463_LC_18_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i11_4_lut_adj_1463_LC_18_20_1  (
            .in0(N__67706),
            .in1(N__56272),
            .in2(N__51801),
            .in3(N__51903),
            .lcout(\c0.n24_adj_4509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_adj_1397_LC_18_20_2 .C_ON=1'b0;
    defparam \c0.i7_2_lut_adj_1397_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_adj_1397_LC_18_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i7_2_lut_adj_1397_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__57886),
            .in2(_gnd_net_),
            .in3(N__59441),
            .lcout(),
            .ltout(\c0.n23187_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1399_LC_18_20_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1399_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1399_LC_18_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1399_LC_18_20_3  (
            .in0(N__51780),
            .in1(N__67194),
            .in2(N__51741),
            .in3(N__66986),
            .lcout(),
            .ltout(\c0.n10_adj_4439_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1402_LC_18_20_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1402_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1402_LC_18_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1402_LC_18_20_4  (
            .in0(N__59738),
            .in1(N__66893),
            .in2(N__51960),
            .in3(N__66929),
            .lcout(),
            .ltout(\c0.n13_adj_4442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1403_LC_18_20_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1403_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1403_LC_18_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1403_LC_18_20_5  (
            .in0(N__51957),
            .in1(N__63276),
            .in2(N__51951),
            .in3(N__61935),
            .lcout(\c0.n24528 ),
            .ltout(\c0.n24528_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1551_LC_18_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1551_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1551_LC_18_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1551_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__73772),
            .in2(N__51948),
            .in3(N__51943),
            .lcout(\c0.n23533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1477_LC_18_21_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1477_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1477_LC_18_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1477_LC_18_21_0  (
            .in0(N__62549),
            .in1(N__63792),
            .in2(N__52101),
            .in3(N__51924),
            .lcout(\c0.n10_adj_4513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1466_LC_18_21_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1466_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1466_LC_18_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1466_LC_18_21_1  (
            .in0(N__63243),
            .in1(N__51915),
            .in2(N__62980),
            .in3(N__51909),
            .lcout(\c0.n24559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1462_LC_18_21_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1462_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1462_LC_18_21_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_4_lut_adj_1462_LC_18_21_3  (
            .in0(N__56854),
            .in1(N__52133),
            .in2(N__56574),
            .in3(N__67505),
            .lcout(\c0.n22_adj_4507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1481_LC_18_21_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1481_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1481_LC_18_21_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1481_LC_18_21_4  (
            .in0(N__52132),
            .in1(N__51969),
            .in2(N__77292),
            .in3(N__56751),
            .lcout(\c0.n23627 ),
            .ltout(\c0.n23627_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1733_LC_18_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1733_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1733_LC_18_21_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1733_LC_18_21_5  (
            .in0(N__52167),
            .in1(N__52206),
            .in2(N__51891),
            .in3(N__51881),
            .lcout(\c0.n21353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1540_LC_18_21_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1540_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1540_LC_18_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1540_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__52166),
            .in2(_gnd_net_),
            .in3(N__63242),
            .lcout(\c0.n10_adj_4575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i205_LC_18_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i205_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i205_LC_18_22_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i205_LC_18_22_1  (
            .in0(N__74135),
            .in1(N__59868),
            .in2(N__71921),
            .in3(N__79397),
            .lcout(\c0.data_in_frame_25_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1519_LC_18_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1519_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1519_LC_18_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1519_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__67140),
            .in2(_gnd_net_),
            .in3(N__52090),
            .lcout(\c0.n22505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i221_LC_18_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i221_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i221_LC_18_22_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i221_LC_18_22_3  (
            .in0(N__76655),
            .in1(N__71866),
            .in2(N__57081),
            .in3(N__79398),
            .lcout(\c0.data_in_frame_27_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i220_LC_18_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i220_LC_18_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i220_LC_18_22_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i220_LC_18_22_4  (
            .in0(N__79396),
            .in1(N__76944),
            .in2(N__57112),
            .in3(N__76656),
            .lcout(\c0.data_in_frame_27_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_345_2_lut_LC_18_22_5 .C_ON=1'b0;
    defparam \c0.i1_rep_345_2_lut_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_345_2_lut_LC_18_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_rep_345_2_lut_LC_18_22_5  (
            .in0(_gnd_net_),
            .in1(N__57102),
            .in2(_gnd_net_),
            .in3(N__57072),
            .lcout(\c0.n25467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1504_LC_18_22_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1504_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1504_LC_18_22_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1504_LC_18_22_6  (
            .in0(N__67883),
            .in1(N__52029),
            .in2(N__52017),
            .in3(N__51999),
            .lcout(\c0.n10_adj_4544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1487_LC_18_22_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1487_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1487_LC_18_22_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1487_LC_18_22_7  (
            .in0(N__52110),
            .in1(N__59867),
            .in2(N__51984),
            .in3(N__56753),
            .lcout(\c0.n10874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_17_i3_2_lut_LC_18_23_0 .C_ON=1'b0;
    defparam \c0.select_367_Select_17_i3_2_lut_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_17_i3_2_lut_LC_18_23_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_17_i3_2_lut_LC_18_23_0  (
            .in0(N__53099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71471),
            .lcout(\c0.n3_adj_4402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_19_i3_2_lut_LC_18_23_1 .C_ON=1'b0;
    defparam \c0.select_367_Select_19_i3_2_lut_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_19_i3_2_lut_LC_18_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_19_i3_2_lut_LC_18_23_1  (
            .in0(N__71472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53180),
            .lcout(\c0.n3_adj_4398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_1755_LC_18_23_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_1755_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_1755_LC_18_23_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_1755_LC_18_23_2  (
            .in0(N__56372),
            .in1(_gnd_net_),
            .in2(N__56407),
            .in3(N__63240),
            .lcout(\c0.n10_adj_4371 ),
            .ltout(\c0.n10_adj_4371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1391_LC_18_23_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1391_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1391_LC_18_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1391_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__52134),
            .in2(N__52113),
            .in3(N__56522),
            .lcout(\c0.n12_adj_4372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_20_i3_2_lut_LC_18_23_4 .C_ON=1'b0;
    defparam \c0.select_367_Select_20_i3_2_lut_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_20_i3_2_lut_LC_18_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_20_i3_2_lut_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__53136),
            .in2(_gnd_net_),
            .in3(N__71473),
            .lcout(\c0.n3_adj_4396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1724_LC_18_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1724_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1724_LC_18_23_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_1724_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__56239),
            .in2(_gnd_net_),
            .in3(N__62317),
            .lcout(\c0.n12_adj_4671 ),
            .ltout(\c0.n12_adj_4671_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i235_LC_18_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i235_LC_18_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i235_LC_18_23_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i235_LC_18_23_6  (
            .in0(N__79125),
            .in1(N__56705),
            .in2(N__52104),
            .in3(N__75393),
            .lcout(\c0.data_in_frame_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3725_2_lut_LC_18_23_7 .C_ON=1'b0;
    defparam \c0.i3725_2_lut_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3725_2_lut_LC_18_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3725_2_lut_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__56396),
            .in2(_gnd_net_),
            .in3(N__56371),
            .lcout(\c0.n6404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_LC_18_24_0 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_LC_18_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_LC_18_24_0  (
            .in0(N__63906),
            .in1(N__56797),
            .in2(N__57001),
            .in3(N__74874),
            .lcout(\c0.n23_adj_4551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_21_i3_2_lut_LC_18_24_1 .C_ON=1'b0;
    defparam \c0.select_367_Select_21_i3_2_lut_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_21_i3_2_lut_LC_18_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_21_i3_2_lut_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(N__53220),
            .in2(_gnd_net_),
            .in3(N__71394),
            .lcout(\c0.n3_adj_4394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1503_LC_18_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1503_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1503_LC_18_24_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1503_LC_18_24_2  (
            .in0(N__63907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56798),
            .lcout(\c0.n22227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i208_LC_18_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i208_LC_18_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i208_LC_18_24_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i208_LC_18_24_3  (
            .in0(N__74203),
            .in1(N__76354),
            .in2(N__63917),
            .in3(N__79440),
            .lcout(\c0.data_in_frame_25_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1453_LC_18_24_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1453_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1453_LC_18_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1453_LC_18_24_4  (
            .in0(N__74837),
            .in1(N__75969),
            .in2(N__52245),
            .in3(N__59901),
            .lcout(\c0.n22_adj_4498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i201_LC_18_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i201_LC_18_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i201_LC_18_24_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i201_LC_18_24_5  (
            .in0(N__74202),
            .in1(N__80703),
            .in2(N__79477),
            .in3(N__56994),
            .lcout(\c0.data_in_frame_25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i206_LC_18_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i206_LC_18_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i206_LC_18_24_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i206_LC_18_24_6  (
            .in0(N__79439),
            .in1(N__74204),
            .in2(N__56816),
            .in3(N__79627),
            .lcout(\c0.data_in_frame_25_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1273_LC_18_24_7 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1273_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1273_LC_18_24_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_adj_1273_LC_18_24_7  (
            .in0(N__52481),
            .in1(N__53376),
            .in2(N__53181),
            .in3(N__52694),
            .lcout(\c0.n45_adj_4298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1482_LC_18_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1482_LC_18_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1482_LC_18_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1482_LC_18_25_2  (
            .in0(_gnd_net_),
            .in1(N__52155),
            .in2(_gnd_net_),
            .in3(N__52191),
            .lcout(\c0.n22334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1250_LC_18_25_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1250_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1250_LC_18_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_adj_1250_LC_18_25_3  (
            .in0(N__53341),
            .in1(N__53219),
            .in2(N__53103),
            .in3(N__53514),
            .lcout(\c0.n44_adj_4270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i203_LC_18_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i203_LC_18_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i203_LC_18_25_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i203_LC_18_25_5  (
            .in0(N__79441),
            .in1(N__79172),
            .in2(N__52165),
            .in3(N__74209),
            .lcout(\c0.data_in_frame_25_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_12_i3_2_lut_LC_18_25_6 .C_ON=1'b0;
    defparam \c0.select_367_Select_12_i3_2_lut_LC_18_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_12_i3_2_lut_LC_18_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_12_i3_2_lut_LC_18_25_6  (
            .in0(_gnd_net_),
            .in1(N__52905),
            .in2(_gnd_net_),
            .in3(N__71454),
            .lcout(\c0.n3_adj_4412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1269_LC_18_26_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1269_LC_18_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1269_LC_18_26_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_1269_LC_18_26_0  (
            .in0(N__53007),
            .in1(N__52721),
            .in2(N__53487),
            .in3(N__70400),
            .lcout(\c0.n40_adj_4294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_10_i3_2_lut_LC_18_26_2 .C_ON=1'b0;
    defparam \c0.select_367_Select_10_i3_2_lut_LC_18_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_10_i3_2_lut_LC_18_26_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_10_i3_2_lut_LC_18_26_2  (
            .in0(_gnd_net_),
            .in1(N__52722),
            .in2(_gnd_net_),
            .in3(N__71455),
            .lcout(\c0.n3_adj_4416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_25_i3_2_lut_LC_18_26_4 .C_ON=1'b0;
    defparam \c0.select_367_Select_25_i3_2_lut_LC_18_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_25_i3_2_lut_LC_18_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_25_i3_2_lut_LC_18_26_4  (
            .in0(_gnd_net_),
            .in1(N__53375),
            .in2(_gnd_net_),
            .in3(N__71456),
            .lcout(\c0.n3_adj_4386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_18_26_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_18_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_18_26_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_LC_18_26_5  (
            .in0(N__52552),
            .in1(N__71588),
            .in2(N__53313),
            .in3(N__53547),
            .lcout(),
            .ltout(\c0.n42_adj_4272_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_1271_LC_18_26_6 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_1271_LC_18_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_1271_LC_18_26_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i24_4_lut_adj_1271_LC_18_26_6  (
            .in0(N__52251),
            .in1(N__52272),
            .in2(N__52266),
            .in3(N__52263),
            .lcout(\c0.n50_adj_4296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_18_27_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_18_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_18_27_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_LC_18_27_1  (
            .in0(N__52628),
            .in1(N__53132),
            .in2(N__52959),
            .in3(N__52904),
            .lcout(\c0.n43_adj_4275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_26_i3_2_lut_LC_18_27_5 .C_ON=1'b0;
    defparam \c0.select_367_Select_26_i3_2_lut_LC_18_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_26_i3_2_lut_LC_18_27_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_26_i3_2_lut_LC_18_27_5  (
            .in0(N__71457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53408),
            .lcout(\c0.n3_adj_4384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_27_i3_2_lut_LC_18_28_0 .C_ON=1'b0;
    defparam \c0.select_367_Select_27_i3_2_lut_LC_18_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_27_i3_2_lut_LC_18_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_27_i3_2_lut_LC_18_28_0  (
            .in0(_gnd_net_),
            .in1(N__53441),
            .in2(_gnd_net_),
            .in3(N__71458),
            .lcout(\c0.n3_adj_4382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_28_i3_2_lut_LC_18_29_1 .C_ON=1'b0;
    defparam \c0.select_367_Select_28_i3_2_lut_LC_18_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_28_i3_2_lut_LC_18_29_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_367_Select_28_i3_2_lut_LC_18_29_1  (
            .in0(N__71504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53480),
            .lcout(\c0.n3_adj_4380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_29_i3_2_lut_LC_18_30_4 .C_ON=1'b0;
    defparam \c0.select_367_Select_29_i3_2_lut_LC_18_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_29_i3_2_lut_LC_18_30_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_29_i3_2_lut_LC_18_30_4  (
            .in0(_gnd_net_),
            .in1(N__53543),
            .in2(_gnd_net_),
            .in3(N__71505),
            .lcout(\c0.n3_adj_4378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_30_i3_2_lut_LC_18_31_0 .C_ON=1'b0;
    defparam \c0.select_367_Select_30_i3_2_lut_LC_18_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_30_i3_2_lut_LC_18_31_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_30_i3_2_lut_LC_18_31_0  (
            .in0(_gnd_net_),
            .in1(N__53510),
            .in2(_gnd_net_),
            .in3(N__71506),
            .lcout(\c0.n3_adj_4376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i0_LC_19_1_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i0_LC_19_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i0_LC_19_1_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_19_1_0  (
            .in0(_gnd_net_),
            .in1(N__74238),
            .in2(N__52284),
            .in3(N__53765),
            .lcout(\c0.FRAME_MATCHER_i_0 ),
            .ltout(),
            .carryin(bfn_19_1_0_),
            .carryout(\c0.n19625 ),
            .clk(N__78825),
            .ce(),
            .sr(N__54903));
    defparam \c0.add_49_2_THRU_CRY_0_LC_19_1_1 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_0_LC_19_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_0_LC_19_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_0_LC_19_1_1  (
            .in0(_gnd_net_),
            .in1(N__54581),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625 ),
            .carryout(\c0.n19625_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_1_LC_19_1_2 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_1_LC_19_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_1_LC_19_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_1_LC_19_1_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54630),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19625_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_2_LC_19_1_3 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_2_LC_19_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_2_LC_19_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_2_LC_19_1_3  (
            .in0(_gnd_net_),
            .in1(N__54585),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19625_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_3_LC_19_1_4 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_3_LC_19_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_3_LC_19_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_3_LC_19_1_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54631),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19625_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_4_LC_19_1_5 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_4_LC_19_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_4_LC_19_1_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_4_LC_19_1_5  (
            .in0(_gnd_net_),
            .in1(N__54589),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19625_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_5_LC_19_1_6 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_5_LC_19_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_5_LC_19_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_5_LC_19_1_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19625_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_6_LC_19_1_7 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_6_LC_19_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_6_LC_19_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_6_LC_19_1_7  (
            .in0(_gnd_net_),
            .in1(N__54593),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19625_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19625_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i1_LC_19_2_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i1_LC_19_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_19_2_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_19_2_0  (
            .in0(N__53764),
            .in1(N__74406),
            .in2(_gnd_net_),
            .in3(N__52275),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(bfn_19_2_0_),
            .carryout(\c0.n19626 ),
            .clk(N__78823),
            .ce(),
            .sr(N__52317));
    defparam \c0.add_49_3_THRU_CRY_0_LC_19_2_1 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_0_LC_19_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_0_LC_19_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_0_LC_19_2_1  (
            .in0(_gnd_net_),
            .in1(N__54462),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626 ),
            .carryout(\c0.n19626_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_1_LC_19_2_2 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_1_LC_19_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_1_LC_19_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_1_LC_19_2_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54578),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19626_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_2_LC_19_2_3 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_2_LC_19_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_2_LC_19_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_2_LC_19_2_3  (
            .in0(_gnd_net_),
            .in1(N__54466),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19626_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_3_LC_19_2_4 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_3_LC_19_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_3_LC_19_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_3_LC_19_2_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19626_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_4_LC_19_2_5 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_4_LC_19_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_4_LC_19_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_4_LC_19_2_5  (
            .in0(_gnd_net_),
            .in1(N__54470),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19626_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_5_LC_19_2_6 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_5_LC_19_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_5_LC_19_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_5_LC_19_2_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19626_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_6_LC_19_2_7 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_6_LC_19_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_6_LC_19_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_6_LC_19_2_7  (
            .in0(_gnd_net_),
            .in1(N__54474),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19626_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19626_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_19_3_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i2_LC_19_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_19_3_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_19_3_0  (
            .in0(N__53769),
            .in1(N__74562),
            .in2(_gnd_net_),
            .in3(N__52302),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(bfn_19_3_0_),
            .carryout(\c0.n19627 ),
            .clk(N__78821),
            .ce(),
            .sr(N__52299));
    defparam \c0.add_49_4_THRU_CRY_0_LC_19_3_1 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_0_LC_19_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_0_LC_19_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_0_LC_19_3_1  (
            .in0(_gnd_net_),
            .in1(N__54449),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627 ),
            .carryout(\c0.n19627_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_1_LC_19_3_2 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_1_LC_19_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_1_LC_19_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_1_LC_19_3_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19627_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_2_LC_19_3_3 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_2_LC_19_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_2_LC_19_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_2_LC_19_3_3  (
            .in0(_gnd_net_),
            .in1(N__54453),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19627_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_3_LC_19_3_4 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_3_LC_19_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_3_LC_19_3_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_3_LC_19_3_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54576),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19627_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_4_LC_19_3_5 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_4_LC_19_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_4_LC_19_3_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_4_LC_19_3_5  (
            .in0(_gnd_net_),
            .in1(N__54457),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19627_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_5_LC_19_3_6 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_5_LC_19_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_5_LC_19_3_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_5_LC_19_3_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54577),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19627_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_6_LC_19_3_7 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_6_LC_19_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_6_LC_19_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_6_LC_19_3_7  (
            .in0(_gnd_net_),
            .in1(N__54461),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19627_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19627_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i3_LC_19_4_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i3_LC_19_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_19_4_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_19_4_0  (
            .in0(N__53760),
            .in1(N__62197),
            .in2(_gnd_net_),
            .in3(N__52320),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(bfn_19_4_0_),
            .carryout(\c0.n19628 ),
            .clk(N__78817),
            .ce(),
            .sr(N__62166));
    defparam \c0.add_49_5_THRU_CRY_0_LC_19_4_1 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_0_LC_19_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_0_LC_19_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_0_LC_19_4_1  (
            .in0(_gnd_net_),
            .in1(N__54436),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628 ),
            .carryout(\c0.n19628_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_1_LC_19_4_2 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_1_LC_19_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_1_LC_19_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_1_LC_19_4_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54572),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19628_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_2_LC_19_4_3 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_2_LC_19_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_2_LC_19_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_2_LC_19_4_3  (
            .in0(_gnd_net_),
            .in1(N__54440),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19628_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_3_LC_19_4_4 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_3_LC_19_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_3_LC_19_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_3_LC_19_4_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19628_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_4_LC_19_4_5 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_4_LC_19_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_4_LC_19_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_4_LC_19_4_5  (
            .in0(_gnd_net_),
            .in1(N__54444),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19628_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_5_LC_19_4_6 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_5_LC_19_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_5_LC_19_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_5_LC_19_4_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54574),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19628_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_6_LC_19_4_7 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_6_LC_19_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_6_LC_19_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_6_LC_19_4_7  (
            .in0(_gnd_net_),
            .in1(N__54448),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19628_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19628_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i4_LC_19_5_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i4_LC_19_5_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_19_5_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_19_5_0  (
            .in0(N__53759),
            .in1(N__52362),
            .in2(_gnd_net_),
            .in3(N__52335),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(bfn_19_5_0_),
            .carryout(\c0.n19629 ),
            .clk(N__78813),
            .ce(),
            .sr(N__52332));
    defparam \c0.add_49_6_THRU_CRY_0_LC_19_5_1 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_0_LC_19_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_0_LC_19_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_0_LC_19_5_1  (
            .in0(_gnd_net_),
            .in1(N__54423),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629 ),
            .carryout(\c0.n19629_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_1_LC_19_5_2 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_1_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_1_LC_19_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_1_LC_19_5_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54569),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19629_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_2_LC_19_5_3 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_2_LC_19_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_2_LC_19_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_2_LC_19_5_3  (
            .in0(_gnd_net_),
            .in1(N__54427),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19629_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_3_LC_19_5_4 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_3_LC_19_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_3_LC_19_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_3_LC_19_5_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54570),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19629_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_4_LC_19_5_5 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_4_LC_19_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_4_LC_19_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_4_LC_19_5_5  (
            .in0(_gnd_net_),
            .in1(N__54431),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19629_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_5_LC_19_5_6 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_5_LC_19_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_5_LC_19_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_5_LC_19_5_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19629_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_6_LC_19_5_7 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_6_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_6_LC_19_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_6_LC_19_5_7  (
            .in0(_gnd_net_),
            .in1(N__54435),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19629_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19629_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_19_6_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i5_LC_19_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_19_6_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_19_6_0  (
            .in0(N__53748),
            .in1(N__52454),
            .in2(_gnd_net_),
            .in3(N__52425),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(bfn_19_6_0_),
            .carryout(\c0.n19630 ),
            .clk(N__78804),
            .ce(),
            .sr(N__52422));
    defparam \c0.add_49_7_THRU_CRY_0_LC_19_6_1 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_0_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_0_LC_19_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_0_LC_19_6_1  (
            .in0(_gnd_net_),
            .in1(N__54231),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630 ),
            .carryout(\c0.n19630_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_1_LC_19_6_2 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_1_LC_19_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_1_LC_19_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_1_LC_19_6_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54420),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19630_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_2_LC_19_6_3 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_2_LC_19_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_2_LC_19_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_2_LC_19_6_3  (
            .in0(_gnd_net_),
            .in1(N__54235),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19630_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_3_LC_19_6_4 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_3_LC_19_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_3_LC_19_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_3_LC_19_6_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54421),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19630_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_4_LC_19_6_5 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_4_LC_19_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_4_LC_19_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_4_LC_19_6_5  (
            .in0(_gnd_net_),
            .in1(N__54239),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19630_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_5_LC_19_6_6 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_5_LC_19_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_5_LC_19_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_5_LC_19_6_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54422),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19630_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_6_LC_19_6_7 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_6_LC_19_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_6_LC_19_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_6_LC_19_6_7  (
            .in0(_gnd_net_),
            .in1(N__54243),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19630_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19630_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i6_LC_19_7_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i6_LC_19_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_19_7_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_19_7_0  (
            .in0(N__53747),
            .in1(N__52525),
            .in2(_gnd_net_),
            .in3(N__52509),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\c0.n19631 ),
            .clk(N__78795),
            .ce(),
            .sr(N__52506));
    defparam \c0.add_49_8_THRU_CRY_0_LC_19_7_1 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_0_LC_19_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_0_LC_19_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_0_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(N__54218),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631 ),
            .carryout(\c0.n19631_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_1_LC_19_7_2 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_1_LC_19_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_1_LC_19_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_1_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19631_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_2_LC_19_7_3 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_2_LC_19_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_2_LC_19_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_2_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__54222),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19631_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_3_LC_19_7_4 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_3_LC_19_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_3_LC_19_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_3_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54418),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19631_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_4_LC_19_7_5 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_4_LC_19_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_4_LC_19_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_4_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(N__54226),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19631_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_5_LC_19_7_6 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_5_LC_19_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_5_LC_19_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_5_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54419),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19631_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_6_LC_19_7_7 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_6_LC_19_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_6_LC_19_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_6_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(N__54230),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19631_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19631_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i7_LC_19_8_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i7_LC_19_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_19_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_19_8_0  (
            .in0(N__53746),
            .in1(N__52615),
            .in2(_gnd_net_),
            .in3(N__52599),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(bfn_19_8_0_),
            .carryout(\c0.n19632 ),
            .clk(N__78788),
            .ce(),
            .sr(N__52596));
    defparam \c0.add_49_9_THRU_CRY_0_LC_19_8_1 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_0_LC_19_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_0_LC_19_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_0_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(N__54138),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632 ),
            .carryout(\c0.n19632_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_1_LC_19_8_2 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_1_LC_19_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_1_LC_19_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_1_LC_19_8_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54314),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19632_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_2_LC_19_8_3 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_2_LC_19_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_2_LC_19_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_2_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(N__54142),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19632_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_3_LC_19_8_4 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_3_LC_19_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_3_LC_19_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_3_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54315),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19632_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_4_LC_19_8_5 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_4_LC_19_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_4_LC_19_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_4_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(N__54146),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19632_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_5_LC_19_8_6 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_5_LC_19_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_5_LC_19_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_5_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19632_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_6_LC_19_8_7 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_6_LC_19_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_6_LC_19_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_6_LC_19_8_7  (
            .in0(_gnd_net_),
            .in1(N__54150),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19632_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19632_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i8_LC_19_9_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i8_LC_19_9_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_19_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_19_9_0  (
            .in0(N__53745),
            .in1(N__52669),
            .in2(_gnd_net_),
            .in3(N__52653),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(bfn_19_9_0_),
            .carryout(\c0.n19633 ),
            .clk(N__78782),
            .ce(),
            .sr(N__52650));
    defparam \c0.add_49_10_THRU_CRY_0_LC_19_9_1 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_0_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_0_LC_19_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_0_LC_19_9_1  (
            .in0(_gnd_net_),
            .in1(N__53995),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633 ),
            .carryout(\c0.n19633_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_1_LC_19_9_2 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_1_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_1_LC_19_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_1_LC_19_9_2  (
            .in0(_gnd_net_),
            .in1(N__53999),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19633_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_2_LC_19_9_3 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_2_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_2_LC_19_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_2_LC_19_9_3  (
            .in0(_gnd_net_),
            .in1(N__53996),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19633_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_3_LC_19_9_4 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_3_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_3_LC_19_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_3_LC_19_9_4  (
            .in0(_gnd_net_),
            .in1(N__54000),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19633_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_4_LC_19_9_5 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_4_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_4_LC_19_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_4_LC_19_9_5  (
            .in0(_gnd_net_),
            .in1(N__53997),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19633_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_5_LC_19_9_6 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_5_LC_19_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_5_LC_19_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_5_LC_19_9_6  (
            .in0(_gnd_net_),
            .in1(N__54001),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19633_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_6_LC_19_9_7 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_6_LC_19_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_6_LC_19_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_6_LC_19_9_7  (
            .in0(_gnd_net_),
            .in1(N__53998),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19633_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19633_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i9_LC_19_10_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i9_LC_19_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_19_10_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_19_10_0  (
            .in0(N__53744),
            .in1(N__52756),
            .in2(_gnd_net_),
            .in3(N__52740),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(bfn_19_10_0_),
            .carryout(\c0.n19634 ),
            .clk(N__78772),
            .ce(),
            .sr(N__52737));
    defparam \c0.add_49_11_THRU_CRY_0_LC_19_10_1 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_0_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_0_LC_19_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_0_LC_19_10_1  (
            .in0(_gnd_net_),
            .in1(N__54307),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634 ),
            .carryout(\c0.n19634_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_1_LC_19_10_2 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_1_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_1_LC_19_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_1_LC_19_10_2  (
            .in0(_gnd_net_),
            .in1(N__54311),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19634_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_2_LC_19_10_3 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_2_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_2_LC_19_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_2_LC_19_10_3  (
            .in0(_gnd_net_),
            .in1(N__54308),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19634_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_3_LC_19_10_4 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_3_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_3_LC_19_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_3_LC_19_10_4  (
            .in0(_gnd_net_),
            .in1(N__54312),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19634_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_4_LC_19_10_5 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_4_LC_19_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_4_LC_19_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_4_LC_19_10_5  (
            .in0(_gnd_net_),
            .in1(N__54309),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19634_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_5_LC_19_10_6 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_5_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_5_LC_19_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_5_LC_19_10_6  (
            .in0(_gnd_net_),
            .in1(N__54313),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19634_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_6_LC_19_10_7 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_6_LC_19_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_6_LC_19_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_6_LC_19_10_7  (
            .in0(_gnd_net_),
            .in1(N__54310),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19634_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19634_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i10_LC_19_11_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i10_LC_19_11_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_19_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_19_11_0  (
            .in0(N__53743),
            .in1(N__52712),
            .in2(_gnd_net_),
            .in3(N__52698),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(bfn_19_11_0_),
            .carryout(\c0.n19635 ),
            .clk(N__78761),
            .ce(),
            .sr(N__52854));
    defparam \c0.add_49_12_THRU_CRY_0_LC_19_11_1 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_0_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_0_LC_19_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_0_LC_19_11_1  (
            .in0(_gnd_net_),
            .in1(N__54317),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635 ),
            .carryout(\c0.n19635_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_1_LC_19_11_2 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_1_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_1_LC_19_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_1_LC_19_11_2  (
            .in0(_gnd_net_),
            .in1(N__54321),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19635_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_2_LC_19_11_3 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_2_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_2_LC_19_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_2_LC_19_11_3  (
            .in0(_gnd_net_),
            .in1(N__54318),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19635_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_3_LC_19_11_4 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_3_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_3_LC_19_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_3_LC_19_11_4  (
            .in0(_gnd_net_),
            .in1(N__54322),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19635_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_4_LC_19_11_5 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_4_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_4_LC_19_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_4_LC_19_11_5  (
            .in0(_gnd_net_),
            .in1(N__54319),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19635_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_5_LC_19_11_6 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_5_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_5_LC_19_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_5_LC_19_11_6  (
            .in0(_gnd_net_),
            .in1(N__54323),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19635_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_6_LC_19_11_7 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_6_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_6_LC_19_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_6_LC_19_11_7  (
            .in0(_gnd_net_),
            .in1(N__54320),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19635_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19635_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i11_LC_19_12_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i11_LC_19_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_19_12_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_19_12_0  (
            .in0(N__53742),
            .in1(N__52816),
            .in2(_gnd_net_),
            .in3(N__52800),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(bfn_19_12_0_),
            .carryout(\c0.n19636 ),
            .clk(N__78749),
            .ce(),
            .sr(N__52797));
    defparam \c0.add_49_13_THRU_CRY_0_LC_19_12_1 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_0_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_0_LC_19_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_0_LC_19_12_1  (
            .in0(_gnd_net_),
            .in1(N__54324),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636 ),
            .carryout(\c0.n19636_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_1_LC_19_12_2 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_1_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_1_LC_19_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_1_LC_19_12_2  (
            .in0(_gnd_net_),
            .in1(N__54328),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19636_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_2_LC_19_12_3 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_2_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_2_LC_19_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_2_LC_19_12_3  (
            .in0(_gnd_net_),
            .in1(N__54325),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19636_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_3_LC_19_12_4 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_3_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_3_LC_19_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_3_LC_19_12_4  (
            .in0(_gnd_net_),
            .in1(N__54329),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19636_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_4_LC_19_12_5 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_4_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_4_LC_19_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_4_LC_19_12_5  (
            .in0(_gnd_net_),
            .in1(N__54326),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19636_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_5_LC_19_12_6 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_5_LC_19_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_5_LC_19_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_5_LC_19_12_6  (
            .in0(_gnd_net_),
            .in1(N__54330),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19636_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_6_LC_19_12_7 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_6_LC_19_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_6_LC_19_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_6_LC_19_12_7  (
            .in0(_gnd_net_),
            .in1(N__54327),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19636_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19636_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_19_13_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i12_LC_19_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_19_13_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_19_13_0  (
            .in0(N__53741),
            .in1(N__52891),
            .in2(_gnd_net_),
            .in3(N__52875),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(bfn_19_13_0_),
            .carryout(\c0.n19637 ),
            .clk(N__78736),
            .ce(),
            .sr(N__52872));
    defparam \c0.add_49_14_THRU_CRY_0_LC_19_13_1 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_0_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_0_LC_19_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_0_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(N__54331),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637 ),
            .carryout(\c0.n19637_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_1_LC_19_13_2 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_1_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_1_LC_19_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_1_LC_19_13_2  (
            .in0(_gnd_net_),
            .in1(N__54335),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19637_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_2_LC_19_13_3 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_2_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_2_LC_19_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_2_LC_19_13_3  (
            .in0(_gnd_net_),
            .in1(N__54332),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19637_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_3_LC_19_13_4 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_3_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_3_LC_19_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_3_LC_19_13_4  (
            .in0(_gnd_net_),
            .in1(N__54336),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19637_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_4_LC_19_13_5 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_4_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_4_LC_19_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_4_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(N__54333),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19637_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_5_LC_19_13_6 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_5_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_5_LC_19_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_5_LC_19_13_6  (
            .in0(_gnd_net_),
            .in1(N__54337),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19637_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_6_LC_19_13_7 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_6_LC_19_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_6_LC_19_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_6_LC_19_13_7  (
            .in0(_gnd_net_),
            .in1(N__54334),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19637_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19637_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i13_LC_19_14_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i13_LC_19_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_19_14_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_19_14_0  (
            .in0(N__53740),
            .in1(N__70387),
            .in2(_gnd_net_),
            .in3(N__52908),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(bfn_19_14_0_),
            .carryout(\c0.n19638 ),
            .clk(N__78723),
            .ce(),
            .sr(N__70368));
    defparam \c0.add_49_15_THRU_CRY_0_LC_19_14_1 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_0_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_0_LC_19_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_0_LC_19_14_1  (
            .in0(_gnd_net_),
            .in1(N__54490),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638 ),
            .carryout(\c0.n19638_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_1_LC_19_14_2 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_1_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_1_LC_19_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_1_LC_19_14_2  (
            .in0(_gnd_net_),
            .in1(N__54494),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19638_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_2_LC_19_14_3 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_2_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_2_LC_19_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_2_LC_19_14_3  (
            .in0(_gnd_net_),
            .in1(N__54491),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19638_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_3_LC_19_14_4 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_3_LC_19_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_3_LC_19_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_3_LC_19_14_4  (
            .in0(_gnd_net_),
            .in1(N__54495),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19638_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_4_LC_19_14_5 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_4_LC_19_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_4_LC_19_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_4_LC_19_14_5  (
            .in0(_gnd_net_),
            .in1(N__54492),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19638_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_5_LC_19_14_6 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_5_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_5_LC_19_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_5_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(N__54496),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19638_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_6_LC_19_14_7 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_6_LC_19_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_6_LC_19_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_6_LC_19_14_7  (
            .in0(_gnd_net_),
            .in1(N__54493),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19638_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19638_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i14_LC_19_15_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i14_LC_19_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_19_15_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_19_15_0  (
            .in0(N__53768),
            .in1(N__52942),
            .in2(_gnd_net_),
            .in3(N__52923),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(bfn_19_15_0_),
            .carryout(\c0.n19639 ),
            .clk(N__78713),
            .ce(),
            .sr(N__52920));
    defparam \c0.add_49_16_THRU_CRY_0_LC_19_15_1 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_0_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_0_LC_19_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_0_LC_19_15_1  (
            .in0(_gnd_net_),
            .in1(N__54497),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639 ),
            .carryout(\c0.n19639_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_1_LC_19_15_2 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_1_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_1_LC_19_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_1_LC_19_15_2  (
            .in0(_gnd_net_),
            .in1(N__54501),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19639_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_2_LC_19_15_3 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_2_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_2_LC_19_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_2_LC_19_15_3  (
            .in0(_gnd_net_),
            .in1(N__54498),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19639_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_3_LC_19_15_4 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_3_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_3_LC_19_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_3_LC_19_15_4  (
            .in0(_gnd_net_),
            .in1(N__54502),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19639_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_4_LC_19_15_5 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_4_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_4_LC_19_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_4_LC_19_15_5  (
            .in0(_gnd_net_),
            .in1(N__54499),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19639_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_5_LC_19_15_6 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_5_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_5_LC_19_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_5_LC_19_15_6  (
            .in0(_gnd_net_),
            .in1(N__54503),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19639_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_6_LC_19_15_7 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_6_LC_19_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_6_LC_19_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_6_LC_19_15_7  (
            .in0(_gnd_net_),
            .in1(N__54500),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19639_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19639_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i15_LC_19_16_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i15_LC_19_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_19_16_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_19_16_0  (
            .in0(N__53767),
            .in1(N__52996),
            .in2(_gnd_net_),
            .in3(N__52977),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(bfn_19_16_0_),
            .carryout(\c0.n19640 ),
            .clk(N__78698),
            .ce(),
            .sr(N__52974));
    defparam \c0.add_49_17_THRU_CRY_0_LC_19_16_1 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_0_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_0_LC_19_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_0_LC_19_16_1  (
            .in0(_gnd_net_),
            .in1(N__54504),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640 ),
            .carryout(\c0.n19640_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_1_LC_19_16_2 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_1_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_1_LC_19_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_1_LC_19_16_2  (
            .in0(_gnd_net_),
            .in1(N__54508),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19640_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_2_LC_19_16_3 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_2_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_2_LC_19_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_2_LC_19_16_3  (
            .in0(_gnd_net_),
            .in1(N__54505),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19640_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_3_LC_19_16_4 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_3_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_3_LC_19_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_3_LC_19_16_4  (
            .in0(_gnd_net_),
            .in1(N__54509),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19640_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_4_LC_19_16_5 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_4_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_4_LC_19_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_4_LC_19_16_5  (
            .in0(_gnd_net_),
            .in1(N__54506),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19640_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_5_LC_19_16_6 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_5_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_5_LC_19_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_5_LC_19_16_6  (
            .in0(_gnd_net_),
            .in1(N__54510),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19640_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_6_LC_19_16_7 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_6_LC_19_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_6_LC_19_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_6_LC_19_16_7  (
            .in0(_gnd_net_),
            .in1(N__54507),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19640_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19640_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_19_17_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i16_LC_19_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_19_17_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_19_17_0  (
            .in0(N__53766),
            .in1(N__53038),
            .in2(_gnd_net_),
            .in3(N__53022),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(bfn_19_17_0_),
            .carryout(\c0.n19641 ),
            .clk(N__78670),
            .ce(),
            .sr(N__53019));
    defparam \c0.add_49_18_THRU_CRY_0_LC_19_17_1 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_0_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_0_LC_19_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_0_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__54511),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641 ),
            .carryout(\c0.n19641_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_1_LC_19_17_2 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_1_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_1_LC_19_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_1_LC_19_17_2  (
            .in0(_gnd_net_),
            .in1(N__54515),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19641_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_2_LC_19_17_3 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_2_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_2_LC_19_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_2_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__54512),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19641_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_3_LC_19_17_4 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_3_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_3_LC_19_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_3_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(N__54516),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19641_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_4_LC_19_17_5 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_4_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_4_LC_19_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_4_LC_19_17_5  (
            .in0(_gnd_net_),
            .in1(N__54513),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19641_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_5_LC_19_17_6 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_5_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_5_LC_19_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_5_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__54517),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19641_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_6_LC_19_17_7 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_6_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_6_LC_19_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_6_LC_19_17_7  (
            .in0(_gnd_net_),
            .in1(N__54514),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19641_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19641_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i17_LC_19_18_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i17_LC_19_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_19_18_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_19_18_0  (
            .in0(N__53724),
            .in1(N__53089),
            .in2(_gnd_net_),
            .in3(N__53073),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(bfn_19_18_0_),
            .carryout(\c0.n19642 ),
            .clk(N__78699),
            .ce(),
            .sr(N__53070));
    defparam \c0.add_49_19_THRU_CRY_0_LC_19_18_1 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_0_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_0_LC_19_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_0_LC_19_18_1  (
            .in0(_gnd_net_),
            .in1(N__54020),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642 ),
            .carryout(\c0.n19642_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_1_LC_19_18_2 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_1_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_1_LC_19_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_1_LC_19_18_2  (
            .in0(_gnd_net_),
            .in1(N__54024),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19642_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_2_LC_19_18_3 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_2_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_2_LC_19_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_2_LC_19_18_3  (
            .in0(_gnd_net_),
            .in1(N__54021),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19642_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_3_LC_19_18_4 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_3_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_3_LC_19_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_3_LC_19_18_4  (
            .in0(_gnd_net_),
            .in1(N__54025),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19642_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_4_LC_19_18_5 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_4_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_4_LC_19_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_4_LC_19_18_5  (
            .in0(_gnd_net_),
            .in1(N__54022),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19642_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_5_LC_19_18_6 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_5_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_5_LC_19_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_5_LC_19_18_6  (
            .in0(_gnd_net_),
            .in1(N__54026),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19642_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_6_LC_19_18_7 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_6_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_6_LC_19_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_6_LC_19_18_7  (
            .in0(_gnd_net_),
            .in1(N__54023),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19642_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19642_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_19_19_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i18_LC_19_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_19_19_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_19_19_0  (
            .in0(N__53749),
            .in1(N__71572),
            .in2(_gnd_net_),
            .in3(N__53106),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(bfn_19_19_0_),
            .carryout(\c0.n19643 ),
            .clk(N__78714),
            .ce(),
            .sr(N__71295));
    defparam \c0.add_49_20_THRU_CRY_0_LC_19_19_1 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_0_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_0_LC_19_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_0_LC_19_19_1  (
            .in0(_gnd_net_),
            .in1(N__54594),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643 ),
            .carryout(\c0.n19643_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_1_LC_19_19_2 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_1_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_1_LC_19_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_1_LC_19_19_2  (
            .in0(_gnd_net_),
            .in1(N__54598),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19643_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_2_LC_19_19_3 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_2_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_2_LC_19_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_2_LC_19_19_3  (
            .in0(_gnd_net_),
            .in1(N__54595),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19643_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_3_LC_19_19_4 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_3_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_3_LC_19_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_3_LC_19_19_4  (
            .in0(_gnd_net_),
            .in1(N__54599),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19643_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_4_LC_19_19_5 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_4_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_4_LC_19_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_4_LC_19_19_5  (
            .in0(_gnd_net_),
            .in1(N__54596),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19643_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_5_LC_19_19_6 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_5_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_5_LC_19_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_5_LC_19_19_6  (
            .in0(_gnd_net_),
            .in1(N__54600),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19643_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_6_LC_19_19_7 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_6_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_6_LC_19_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_6_LC_19_19_7  (
            .in0(_gnd_net_),
            .in1(N__54597),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19643_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19643_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i19_LC_19_20_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i19_LC_19_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_19_20_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_19_20_0  (
            .in0(N__53713),
            .in1(N__53170),
            .in2(_gnd_net_),
            .in3(N__53154),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(bfn_19_20_0_),
            .carryout(\c0.n19644 ),
            .clk(N__78724),
            .ce(),
            .sr(N__53151));
    defparam \c0.add_49_21_THRU_CRY_0_LC_19_20_1 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_0_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_0_LC_19_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_0_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(N__54601),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644 ),
            .carryout(\c0.n19644_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_1_LC_19_20_2 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_1_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_1_LC_19_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_1_LC_19_20_2  (
            .in0(_gnd_net_),
            .in1(N__54605),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19644_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_2_LC_19_20_3 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_2_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_2_LC_19_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_2_LC_19_20_3  (
            .in0(_gnd_net_),
            .in1(N__54602),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19644_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_3_LC_19_20_4 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_3_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_3_LC_19_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_3_LC_19_20_4  (
            .in0(_gnd_net_),
            .in1(N__54606),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19644_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_4_LC_19_20_5 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_4_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_4_LC_19_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_4_LC_19_20_5  (
            .in0(_gnd_net_),
            .in1(N__54603),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19644_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_5_LC_19_20_6 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_5_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_5_LC_19_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_5_LC_19_20_6  (
            .in0(_gnd_net_),
            .in1(N__54607),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19644_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_6_LC_19_20_7 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_6_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_6_LC_19_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_6_LC_19_20_7  (
            .in0(_gnd_net_),
            .in1(N__54604),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19644_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19644_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i20_LC_19_21_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i20_LC_19_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_19_21_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_19_21_0  (
            .in0(N__53712),
            .in1(N__53125),
            .in2(_gnd_net_),
            .in3(N__53109),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(bfn_19_21_0_),
            .carryout(\c0.n19645 ),
            .clk(N__78737),
            .ce(),
            .sr(N__53232));
    defparam \c0.add_49_22_THRU_CRY_0_LC_19_21_1 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_0_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_0_LC_19_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_0_LC_19_21_1  (
            .in0(_gnd_net_),
            .in1(N__54608),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645 ),
            .carryout(\c0.n19645_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_1_LC_19_21_2 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_1_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_1_LC_19_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_1_LC_19_21_2  (
            .in0(_gnd_net_),
            .in1(N__54612),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19645_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_2_LC_19_21_3 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_2_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_2_LC_19_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_2_LC_19_21_3  (
            .in0(_gnd_net_),
            .in1(N__54609),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19645_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_3_LC_19_21_4 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_3_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_3_LC_19_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_3_LC_19_21_4  (
            .in0(_gnd_net_),
            .in1(N__54613),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19645_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_4_LC_19_21_5 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_4_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_4_LC_19_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_4_LC_19_21_5  (
            .in0(_gnd_net_),
            .in1(N__54610),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19645_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_5_LC_19_21_6 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_5_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_5_LC_19_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_5_LC_19_21_6  (
            .in0(_gnd_net_),
            .in1(N__54614),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19645_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_6_LC_19_21_7 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_6_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_6_LC_19_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_6_LC_19_21_7  (
            .in0(_gnd_net_),
            .in1(N__54611),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19645_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19645_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i21_LC_19_22_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i21_LC_19_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_19_22_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_19_22_0  (
            .in0(N__53698),
            .in1(N__53212),
            .in2(_gnd_net_),
            .in3(N__53196),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(bfn_19_22_0_),
            .carryout(\c0.n19646 ),
            .clk(N__78750),
            .ce(),
            .sr(N__53193));
    defparam \c0.add_49_23_THRU_CRY_0_LC_19_22_1 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_0_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_0_LC_19_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_0_LC_19_22_1  (
            .in0(_gnd_net_),
            .in1(N__54714),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646 ),
            .carryout(\c0.n19646_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_1_LC_19_22_2 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_1_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_1_LC_19_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_1_LC_19_22_2  (
            .in0(_gnd_net_),
            .in1(N__54718),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19646_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_2_LC_19_22_3 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_2_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_2_LC_19_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_2_LC_19_22_3  (
            .in0(_gnd_net_),
            .in1(N__54715),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19646_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_3_LC_19_22_4 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_3_LC_19_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_3_LC_19_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_3_LC_19_22_4  (
            .in0(_gnd_net_),
            .in1(N__54719),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19646_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_4_LC_19_22_5 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_4_LC_19_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_4_LC_19_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_4_LC_19_22_5  (
            .in0(_gnd_net_),
            .in1(N__54716),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19646_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_5_LC_19_22_6 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_5_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_5_LC_19_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_5_LC_19_22_6  (
            .in0(_gnd_net_),
            .in1(N__54720),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19646_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_6_LC_19_22_7 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_6_LC_19_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_6_LC_19_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_6_LC_19_22_7  (
            .in0(_gnd_net_),
            .in1(N__54717),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19646_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19646_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i22_LC_19_23_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i22_LC_19_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_19_23_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_19_23_0  (
            .in0(N__53697),
            .in1(N__53263),
            .in2(_gnd_net_),
            .in3(N__53247),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(bfn_19_23_0_),
            .carryout(\c0.n19647 ),
            .clk(N__78762),
            .ce(),
            .sr(N__53244));
    defparam \c0.add_49_24_THRU_CRY_0_LC_19_23_1 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_0_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_0_LC_19_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_0_LC_19_23_1  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54827),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647 ),
            .carryout(\c0.n19647_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_1_LC_19_23_2 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_1_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_1_LC_19_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_1_LC_19_23_2  (
            .in0(_gnd_net_),
            .in1(N__54724),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19647_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_2_LC_19_23_3 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_2_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_2_LC_19_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_2_LC_19_23_3  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54828),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19647_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_3_LC_19_23_4 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_3_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_3_LC_19_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_3_LC_19_23_4  (
            .in0(_gnd_net_),
            .in1(N__54728),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19647_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_4_LC_19_23_5 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_4_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_4_LC_19_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_4_LC_19_23_5  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54829),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19647_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_5_LC_19_23_6 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_5_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_5_LC_19_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_5_LC_19_23_6  (
            .in0(_gnd_net_),
            .in1(N__54732),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19647_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_6_LC_19_23_7 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_6_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_6_LC_19_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_6_LC_19_23_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54830),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19647_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19647_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i23_LC_19_24_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i23_LC_19_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_19_24_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_19_24_0  (
            .in0(N__53696),
            .in1(N__53302),
            .in2(_gnd_net_),
            .in3(N__53283),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(bfn_19_24_0_),
            .carryout(\c0.n19648 ),
            .clk(N__78773),
            .ce(),
            .sr(N__53280));
    defparam \c0.add_49_25_THRU_CRY_0_LC_19_24_1 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_0_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_0_LC_19_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_0_LC_19_24_1  (
            .in0(_gnd_net_),
            .in1(N__54736),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648 ),
            .carryout(\c0.n19648_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_1_LC_19_24_2 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_1_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_1_LC_19_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_1_LC_19_24_2  (
            .in0(_gnd_net_),
            .in1(N__54740),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19648_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_2_LC_19_24_3 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_2_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_2_LC_19_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_2_LC_19_24_3  (
            .in0(_gnd_net_),
            .in1(N__54737),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19648_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_3_LC_19_24_4 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_3_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_3_LC_19_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_3_LC_19_24_4  (
            .in0(_gnd_net_),
            .in1(N__54741),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19648_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_4_LC_19_24_5 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_4_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_4_LC_19_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_4_LC_19_24_5  (
            .in0(_gnd_net_),
            .in1(N__54738),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19648_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_5_LC_19_24_6 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_5_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_5_LC_19_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_5_LC_19_24_6  (
            .in0(_gnd_net_),
            .in1(N__54742),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19648_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_6_LC_19_24_7 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_6_LC_19_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_6_LC_19_24_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_6_LC_19_24_7  (
            .in0(_gnd_net_),
            .in1(N__54739),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19648_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19648_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i24_LC_19_25_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i24_LC_19_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_19_25_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_19_25_0  (
            .in0(N__53695),
            .in1(N__53342),
            .in2(_gnd_net_),
            .in3(N__53325),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(bfn_19_25_0_),
            .carryout(\c0.n19649 ),
            .clk(N__78781),
            .ce(),
            .sr(N__53322));
    defparam \c0.add_49_26_THRU_CRY_0_LC_19_25_1 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_0_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_0_LC_19_25_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_0_LC_19_25_1  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54831),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649 ),
            .carryout(\c0.n19649_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_1_LC_19_25_2 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_1_LC_19_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_1_LC_19_25_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_1_LC_19_25_2  (
            .in0(_gnd_net_),
            .in1(N__54746),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19649_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_2_LC_19_25_3 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_2_LC_19_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_2_LC_19_25_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_2_LC_19_25_3  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54832),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19649_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_3_LC_19_25_4 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_3_LC_19_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_3_LC_19_25_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_3_LC_19_25_4  (
            .in0(_gnd_net_),
            .in1(N__54750),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19649_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_4_LC_19_25_5 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_4_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_4_LC_19_25_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_4_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54833),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19649_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_5_LC_19_25_6 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_5_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_5_LC_19_25_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_5_LC_19_25_6  (
            .in0(_gnd_net_),
            .in1(N__54754),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19649_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_6_LC_19_25_7 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_6_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_6_LC_19_25_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_6_LC_19_25_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__54834),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19649_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19649_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_19_26_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i25_LC_19_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_19_26_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_19_26_0  (
            .in0(N__53694),
            .in1(N__53374),
            .in2(_gnd_net_),
            .in3(N__53355),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(bfn_19_26_0_),
            .carryout(\c0.n19650 ),
            .clk(N__78787),
            .ce(),
            .sr(N__53352));
    defparam \c0.add_49_27_THRU_CRY_0_LC_19_26_1 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_0_LC_19_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_0_LC_19_26_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_0_LC_19_26_1  (
            .in0(_gnd_net_),
            .in1(N__54835),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650 ),
            .carryout(\c0.n19650_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_1_LC_19_26_2 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_1_LC_19_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_1_LC_19_26_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_1_LC_19_26_2  (
            .in0(_gnd_net_),
            .in1(N__54839),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19650_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_2_LC_19_26_3 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_2_LC_19_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_2_LC_19_26_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_2_LC_19_26_3  (
            .in0(_gnd_net_),
            .in1(N__54836),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19650_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_3_LC_19_26_4 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_3_LC_19_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_3_LC_19_26_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_3_LC_19_26_4  (
            .in0(_gnd_net_),
            .in1(N__54840),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19650_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_4_LC_19_26_5 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_4_LC_19_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_4_LC_19_26_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_4_LC_19_26_5  (
            .in0(_gnd_net_),
            .in1(N__54837),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19650_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_5_LC_19_26_6 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_5_LC_19_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_5_LC_19_26_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_5_LC_19_26_6  (
            .in0(_gnd_net_),
            .in1(N__54841),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19650_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_6_LC_19_26_7 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_6_LC_19_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_6_LC_19_26_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_6_LC_19_26_7  (
            .in0(_gnd_net_),
            .in1(N__54838),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19650_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19650_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i26_LC_19_27_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i26_LC_19_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_19_27_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_19_27_0  (
            .in0(N__53693),
            .in1(N__53404),
            .in2(_gnd_net_),
            .in3(N__53385),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(bfn_19_27_0_),
            .carryout(\c0.n19651 ),
            .clk(N__78794),
            .ce(),
            .sr(N__53382));
    defparam \c0.add_49_28_THRU_CRY_0_LC_19_27_1 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_0_LC_19_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_0_LC_19_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_0_LC_19_27_1  (
            .in0(_gnd_net_),
            .in1(N__54842),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651 ),
            .carryout(\c0.n19651_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_1_LC_19_27_2 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_1_LC_19_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_1_LC_19_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_1_LC_19_27_2  (
            .in0(_gnd_net_),
            .in1(N__54846),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19651_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_2_LC_19_27_3 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_2_LC_19_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_2_LC_19_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_2_LC_19_27_3  (
            .in0(_gnd_net_),
            .in1(N__54843),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19651_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_3_LC_19_27_4 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_3_LC_19_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_3_LC_19_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_3_LC_19_27_4  (
            .in0(_gnd_net_),
            .in1(N__54847),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19651_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_4_LC_19_27_5 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_4_LC_19_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_4_LC_19_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_4_LC_19_27_5  (
            .in0(_gnd_net_),
            .in1(N__54844),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19651_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_5_LC_19_27_6 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_5_LC_19_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_5_LC_19_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_5_LC_19_27_6  (
            .in0(_gnd_net_),
            .in1(N__54848),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19651_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_6_LC_19_27_7 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_6_LC_19_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_6_LC_19_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_6_LC_19_27_7  (
            .in0(_gnd_net_),
            .in1(N__54845),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19651_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19651_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i27_LC_19_28_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i27_LC_19_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_19_28_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_19_28_0  (
            .in0(N__53692),
            .in1(N__53440),
            .in2(_gnd_net_),
            .in3(N__53421),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(bfn_19_28_0_),
            .carryout(\c0.n19652 ),
            .clk(N__78803),
            .ce(),
            .sr(N__53418));
    defparam \c0.add_49_29_THRU_CRY_0_LC_19_28_1 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_0_LC_19_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_0_LC_19_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_0_LC_19_28_1  (
            .in0(_gnd_net_),
            .in1(N__54849),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652 ),
            .carryout(\c0.n19652_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_1_LC_19_28_2 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_1_LC_19_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_1_LC_19_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_1_LC_19_28_2  (
            .in0(_gnd_net_),
            .in1(N__54853),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19652_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_2_LC_19_28_3 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_2_LC_19_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_2_LC_19_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_2_LC_19_28_3  (
            .in0(_gnd_net_),
            .in1(N__54850),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19652_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_3_LC_19_28_4 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_3_LC_19_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_3_LC_19_28_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_3_LC_19_28_4  (
            .in0(_gnd_net_),
            .in1(N__54854),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19652_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_4_LC_19_28_5 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_4_LC_19_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_4_LC_19_28_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_4_LC_19_28_5  (
            .in0(_gnd_net_),
            .in1(N__54851),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19652_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_5_LC_19_28_6 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_5_LC_19_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_5_LC_19_28_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_5_LC_19_28_6  (
            .in0(_gnd_net_),
            .in1(N__54855),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19652_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_6_LC_19_28_7 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_6_LC_19_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_6_LC_19_28_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_6_LC_19_28_7  (
            .in0(_gnd_net_),
            .in1(N__54852),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19652_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19652_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i28_LC_19_29_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i28_LC_19_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_19_29_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_19_29_0  (
            .in0(N__53699),
            .in1(N__53479),
            .in2(_gnd_net_),
            .in3(N__53460),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(bfn_19_29_0_),
            .carryout(\c0.n19653 ),
            .clk(N__78812),
            .ce(),
            .sr(N__53457));
    defparam \c0.add_49_30_THRU_CRY_0_LC_19_29_1 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_0_LC_19_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_0_LC_19_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_0_LC_19_29_1  (
            .in0(_gnd_net_),
            .in1(N__54856),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653 ),
            .carryout(\c0.n19653_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_1_LC_19_29_2 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_1_LC_19_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_1_LC_19_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_1_LC_19_29_2  (
            .in0(_gnd_net_),
            .in1(N__54860),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19653_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_2_LC_19_29_3 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_2_LC_19_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_2_LC_19_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_2_LC_19_29_3  (
            .in0(_gnd_net_),
            .in1(N__54857),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19653_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_3_LC_19_29_4 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_3_LC_19_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_3_LC_19_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_3_LC_19_29_4  (
            .in0(_gnd_net_),
            .in1(N__54861),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19653_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_4_LC_19_29_5 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_4_LC_19_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_4_LC_19_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_4_LC_19_29_5  (
            .in0(_gnd_net_),
            .in1(N__54858),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19653_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_5_LC_19_29_6 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_5_LC_19_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_5_LC_19_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_5_LC_19_29_6  (
            .in0(_gnd_net_),
            .in1(N__54862),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19653_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_6_LC_19_29_7 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_6_LC_19_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_6_LC_19_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_6_LC_19_29_7  (
            .in0(_gnd_net_),
            .in1(N__54859),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19653_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19653_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i29_LC_19_30_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i29_LC_19_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_19_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_19_30_0  (
            .in0(N__53665),
            .in1(N__53542),
            .in2(_gnd_net_),
            .in3(N__53523),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(bfn_19_30_0_),
            .carryout(\c0.n19654 ),
            .clk(N__78816),
            .ce(),
            .sr(N__53520));
    defparam \c0.add_49_31_THRU_CRY_0_LC_19_30_1 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_0_LC_19_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_0_LC_19_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_0_LC_19_30_1  (
            .in0(_gnd_net_),
            .in1(N__54131),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654 ),
            .carryout(\c0.n19654_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_1_LC_19_30_2 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_1_LC_19_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_1_LC_19_30_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_1_LC_19_30_2  (
            .in0(_gnd_net_),
            .in1(N__54135),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19654_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_2_LC_19_30_3 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_2_LC_19_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_2_LC_19_30_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_2_LC_19_30_3  (
            .in0(_gnd_net_),
            .in1(N__54132),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19654_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_3_LC_19_30_4 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_3_LC_19_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_3_LC_19_30_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_3_LC_19_30_4  (
            .in0(_gnd_net_),
            .in1(N__54136),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19654_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_4_LC_19_30_5 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_4_LC_19_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_4_LC_19_30_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_4_LC_19_30_5  (
            .in0(_gnd_net_),
            .in1(N__54133),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19654_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_5_LC_19_30_6 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_5_LC_19_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_5_LC_19_30_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_5_LC_19_30_6  (
            .in0(_gnd_net_),
            .in1(N__54137),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19654_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_6_LC_19_30_7 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_6_LC_19_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_6_LC_19_30_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_6_LC_19_30_7  (
            .in0(_gnd_net_),
            .in1(N__54134),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19654_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19654_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i30_LC_19_31_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i30_LC_19_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_19_31_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_19_31_0  (
            .in0(N__53640),
            .in1(N__53509),
            .in2(_gnd_net_),
            .in3(N__53490),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(bfn_19_31_0_),
            .carryout(\c0.n19655 ),
            .clk(N__78820),
            .ce(),
            .sr(N__54894));
    defparam \c0.add_49_32_THRU_CRY_0_LC_19_31_1 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_0_LC_19_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_0_LC_19_31_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_0_LC_19_31_1  (
            .in0(_gnd_net_),
            .in1(N__54879),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655 ),
            .carryout(\c0.n19655_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_1_LC_19_31_2 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_1_LC_19_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_1_LC_19_31_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_1_LC_19_31_2  (
            .in0(_gnd_net_),
            .in1(N__54883),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n19655_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_2_LC_19_31_3 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_2_LC_19_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_2_LC_19_31_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_2_LC_19_31_3  (
            .in0(_gnd_net_),
            .in1(N__54880),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n19655_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_3_LC_19_31_4 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_3_LC_19_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_3_LC_19_31_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_3_LC_19_31_4  (
            .in0(_gnd_net_),
            .in1(N__54884),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n19655_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_4_LC_19_31_5 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_4_LC_19_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_4_LC_19_31_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_4_LC_19_31_5  (
            .in0(_gnd_net_),
            .in1(N__54881),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n19655_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_5_LC_19_31_6 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_5_LC_19_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_5_LC_19_31_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_5_LC_19_31_6  (
            .in0(_gnd_net_),
            .in1(N__54885),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n19655_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_6_LC_19_31_7 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_6_LC_19_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_6_LC_19_31_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_6_LC_19_31_7  (
            .in0(_gnd_net_),
            .in1(N__54882),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n19655_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n19655_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i31_LC_19_32_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_19_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_19_32_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_19_32_0  (
            .in0(N__53641),
            .in1(N__53877),
            .in2(_gnd_net_),
            .in3(N__53919),
            .lcout(\c0.FRAME_MATCHER_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78824),
            .ce(),
            .sr(N__53823));
    defparam \c0.i14251_1_lut_LC_19_32_1 .C_ON=1'b0;
    defparam \c0.i14251_1_lut_LC_19_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14251_1_lut_LC_19_32_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.i14251_1_lut_LC_19_32_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53814),
            .lcout(\c0.n1306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_0_i3_2_lut_LC_20_3_2 .C_ON=1'b0;
    defparam \c0.select_367_Select_0_i3_2_lut_LC_20_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_0_i3_2_lut_LC_20_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_0_i3_2_lut_LC_20_3_2  (
            .in0(_gnd_net_),
            .in1(N__74302),
            .in2(_gnd_net_),
            .in3(N__71552),
            .lcout(\c0.n3_adj_4436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1610_LC_20_7_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1610_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1610_LC_20_7_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1610_LC_20_7_0  (
            .in0(N__60131),
            .in1(N__60686),
            .in2(N__58403),
            .in3(N__60116),
            .lcout(\c0.n23677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i81_LC_20_7_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i81_LC_20_7_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i81_LC_20_7_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i81_LC_20_7_1  (
            .in0(N__73709),
            .in1(N__69183),
            .in2(N__80736),
            .in3(N__58399),
            .lcout(\c0.data_in_frame_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78805),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i41_4_lut_LC_20_7_2 .C_ON=1'b0;
    defparam \c0.i41_4_lut_LC_20_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i41_4_lut_LC_20_7_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i41_4_lut_LC_20_7_2  (
            .in0(N__55100),
            .in1(N__58395),
            .in2(N__69362),
            .in3(N__64529),
            .lcout(\c0.n97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i75_LC_20_7_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i75_LC_20_7_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i75_LC_20_7_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i75_LC_20_7_3  (
            .in0(N__64530),
            .in1(N__79108),
            .in2(N__73719),
            .in3(N__74115),
            .lcout(\c0.data_in_frame_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78805),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i74_LC_20_7_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i74_LC_20_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i74_LC_20_7_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i74_LC_20_7_4  (
            .in0(N__75249),
            .in1(N__74111),
            .in2(N__69363),
            .in3(N__73715),
            .lcout(\c0.data_in_frame_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78805),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13936_4_lut_LC_20_7_5 .C_ON=1'b0;
    defparam \c0.i13936_4_lut_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13936_4_lut_LC_20_7_5 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \c0.i13936_4_lut_LC_20_7_5  (
            .in0(N__57030),
            .in1(N__68757),
            .in2(N__60312),
            .in3(N__59931),
            .lcout(\c0.n17537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i66_LC_20_7_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i66_LC_20_7_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i66_LC_20_7_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i66_LC_20_7_6  (
            .in0(N__75248),
            .in1(N__72880),
            .in2(N__55113),
            .in3(N__73714),
            .lcout(\c0.data_in_frame_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78805),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i83_LC_20_7_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i83_LC_20_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i83_LC_20_7_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i83_LC_20_7_7  (
            .in0(N__73710),
            .in1(N__69184),
            .in2(N__55045),
            .in3(N__79109),
            .lcout(\c0.data_in_frame_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78805),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1613_LC_20_8_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1613_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1613_LC_20_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1613_LC_20_8_0  (
            .in0(N__57322),
            .in1(N__54909),
            .in2(N__55329),
            .in3(N__60295),
            .lcout(\c0.n10_adj_4615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1836_LC_20_8_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1836_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1836_LC_20_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1836_LC_20_8_1  (
            .in0(N__60631),
            .in1(N__54968),
            .in2(_gnd_net_),
            .in3(N__61036),
            .lcout(\c0.n22196 ),
            .ltout(\c0.n22196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_20_8_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_20_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_20_8_2  (
            .in0(N__57323),
            .in1(N__60296),
            .in2(N__54987),
            .in3(N__60741),
            .lcout(\c0.n12_adj_4299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1878_LC_20_8_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1878_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1878_LC_20_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1878_LC_20_8_3  (
            .in0(N__64581),
            .in1(N__70348),
            .in2(_gnd_net_),
            .in3(N__57399),
            .lcout(\c0.n10_adj_4283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1648_LC_20_8_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1648_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1648_LC_20_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1648_LC_20_8_4  (
            .in0(_gnd_net_),
            .in1(N__57355),
            .in2(_gnd_net_),
            .in3(N__55206),
            .lcout(\c0.n11_adj_4280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_20_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_20_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_20_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i8_LC_20_8_5  (
            .in0(N__70155),
            .in1(N__72862),
            .in2(N__60243),
            .in3(N__76316),
            .lcout(\c0.data_in_frame_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1874_LC_20_8_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1874_LC_20_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1874_LC_20_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1874_LC_20_8_6  (
            .in0(N__57365),
            .in1(N__55207),
            .in2(N__57409),
            .in3(N__64768),
            .lcout(\c0.n12_adj_4258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_20_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_20_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_20_8_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i25_LC_20_8_7  (
            .in0(N__70154),
            .in1(N__54969),
            .in2(N__76630),
            .in3(N__80711),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1620_LC_20_9_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1620_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1620_LC_20_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1620_LC_20_9_1  (
            .in0(_gnd_net_),
            .in1(N__68510),
            .in2(N__54960),
            .in3(N__60742),
            .lcout(\c0.n13523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1549_LC_20_9_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1549_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1549_LC_20_9_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_adj_1549_LC_20_9_2  (
            .in0(N__54943),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60186),
            .lcout(\c0.n7_adj_4300 ),
            .ltout(\c0.n7_adj_4300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1278_LC_20_9_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1278_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1278_LC_20_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1278_LC_20_9_3  (
            .in0(N__70742),
            .in1(N__55251),
            .in2(N__55245),
            .in3(N__68511),
            .lcout(\c0.n22316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1694_LC_20_9_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1694_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1694_LC_20_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1694_LC_20_9_4  (
            .in0(N__55134),
            .in1(N__55188),
            .in2(N__55241),
            .in3(N__64773),
            .lcout(\c0.n23655 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1643_LC_20_9_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1643_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1643_LC_20_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1643_LC_20_9_5  (
            .in0(N__60187),
            .in1(N__60635),
            .in2(_gnd_net_),
            .in3(N__60297),
            .lcout(\c0.n23251 ),
            .ltout(\c0.n23251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_4_lut_adj_1664_LC_20_9_6 .C_ON=1'b0;
    defparam \c0.i3_2_lut_4_lut_adj_1664_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_4_lut_adj_1664_LC_20_9_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_4_lut_adj_1664_LC_20_9_6  (
            .in0(N__57377),
            .in1(N__55187),
            .in2(N__55152),
            .in3(N__64772),
            .lcout(\c0.n7_adj_4282 ),
            .ltout(\c0.n7_adj_4282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1260_LC_20_9_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1260_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1260_LC_20_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1260_LC_20_9_7  (
            .in0(N__55630),
            .in1(N__55149),
            .in2(N__55137),
            .in3(N__55133),
            .lcout(\c0.n22472 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1686_LC_20_10_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1686_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1686_LC_20_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1686_LC_20_10_0  (
            .in0(N__55338),
            .in1(N__60235),
            .in2(N__57263),
            .in3(N__57298),
            .lcout(),
            .ltout(\c0.n13_adj_4638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1639_LC_20_10_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1639_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1639_LC_20_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1639_LC_20_10_1  (
            .in0(N__55049),
            .in1(N__55114),
            .in2(N__55080),
            .in3(N__57435),
            .lcout(\c0.n13_adj_4610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_LC_20_10_2 .C_ON=1'b0;
    defparam \c0.i12_2_lut_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_LC_20_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i12_2_lut_LC_20_10_2  (
            .in0(_gnd_net_),
            .in1(N__57297),
            .in2(_gnd_net_),
            .in3(N__60234),
            .lcout(\c0.n68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i42_4_lut_adj_1409_LC_20_10_3 .C_ON=1'b0;
    defparam \c0.i42_4_lut_adj_1409_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i42_4_lut_adj_1409_LC_20_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i42_4_lut_adj_1409_LC_20_10_3  (
            .in0(N__57416),
            .in1(N__55077),
            .in2(N__55050),
            .in3(N__55022),
            .lcout(\c0.n98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1249_LC_20_10_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1249_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1249_LC_20_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1249_LC_20_10_4  (
            .in0(N__57958),
            .in1(N__55362),
            .in2(N__55564),
            .in3(N__55350),
            .lcout(\c0.n4_adj_4269 ),
            .ltout(\c0.n4_adj_4269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_4_lut_LC_20_10_5 .C_ON=1'b0;
    defparam \c0.i33_4_lut_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i33_4_lut_LC_20_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i33_4_lut_LC_20_10_5  (
            .in0(N__55330),
            .in1(N__61859),
            .in2(N__55290),
            .in3(N__60148),
            .lcout(),
            .ltout(\c0.n89_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i45_4_lut_adj_1408_LC_20_10_6 .C_ON=1'b0;
    defparam \c0.i45_4_lut_adj_1408_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i45_4_lut_adj_1408_LC_20_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i45_4_lut_adj_1408_LC_20_10_6  (
            .in0(N__55287),
            .in1(N__60547),
            .in2(N__55281),
            .in3(N__71093),
            .lcout(\c0.n101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1619_LC_20_11_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1619_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1619_LC_20_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1619_LC_20_11_0  (
            .in0(N__71092),
            .in1(N__57186),
            .in2(N__69252),
            .in3(N__70602),
            .lcout(\c0.n22_adj_4622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_20_11_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_20_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_20_11_1  (
            .in0(N__58548),
            .in1(N__57662),
            .in2(N__59265),
            .in3(N__60818),
            .lcout(),
            .ltout(\c0.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_20_11_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_20_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_20_11_2  (
            .in0(N__58281),
            .in1(N__55478),
            .in2(N__55278),
            .in3(N__55767),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_1787_LC_20_11_3 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_1787_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_1787_LC_20_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_1787_LC_20_11_3  (
            .in0(_gnd_net_),
            .in1(N__60817),
            .in2(_gnd_net_),
            .in3(N__58280),
            .lcout(\c0.n13075 ),
            .ltout(\c0.n13075_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i37_4_lut_LC_20_11_4 .C_ON=1'b0;
    defparam \c0.i37_4_lut_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i37_4_lut_LC_20_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i37_4_lut_LC_20_11_4  (
            .in0(N__60792),
            .in1(N__68970),
            .in2(N__55257),
            .in3(N__61294),
            .lcout(),
            .ltout(\c0.n93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i47_4_lut_LC_20_11_5 .C_ON=1'b0;
    defparam \c0.i47_4_lut_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i47_4_lut_LC_20_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i47_4_lut_LC_20_11_5  (
            .in0(N__55766),
            .in1(N__60924),
            .in2(N__55254),
            .in3(N__68750),
            .lcout(\c0.n103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_3_lut_4_lut_LC_20_11_6 .C_ON=1'b0;
    defparam \c0.i13_3_lut_4_lut_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_3_lut_4_lut_LC_20_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_3_lut_4_lut_LC_20_11_6  (
            .in0(N__71091),
            .in1(N__58054),
            .in2(N__57783),
            .in3(N__60080),
            .lcout(\c0.n23156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i66_4_lut_LC_20_12_0 .C_ON=1'b0;
    defparam \c0.i66_4_lut_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i66_4_lut_LC_20_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i66_4_lut_LC_20_12_0  (
            .in0(N__62123),
            .in1(N__55434),
            .in2(N__55392),
            .in3(N__55410),
            .lcout(),
            .ltout(\c0.n147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i74_4_lut_LC_20_12_1 .C_ON=1'b0;
    defparam \c0.i74_4_lut_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i74_4_lut_LC_20_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i74_4_lut_LC_20_12_1  (
            .in0(N__61094),
            .in1(N__70229),
            .in2(N__55401),
            .in3(N__55398),
            .lcout(\c0.n155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i53_4_lut_LC_20_12_2 .C_ON=1'b0;
    defparam \c0.i53_4_lut_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i53_4_lut_LC_20_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i53_4_lut_LC_20_12_2  (
            .in0(N__57684),
            .in1(N__55632),
            .in2(N__57672),
            .in3(N__56005),
            .lcout(\c0.n134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i50_4_lut_LC_20_12_3 .C_ON=1'b0;
    defparam \c0.i50_4_lut_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i50_4_lut_LC_20_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i50_4_lut_LC_20_12_3  (
            .in0(N__70445),
            .in1(N__65576),
            .in2(N__71280),
            .in3(N__62858),
            .lcout(\c0.n131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1262_LC_20_12_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1262_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1262_LC_20_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1262_LC_20_12_4  (
            .in0(N__69837),
            .in1(N__70444),
            .in2(N__62859),
            .in3(N__55839),
            .lcout(\c0.n31_adj_4284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_3_lut_4_lut_LC_20_12_5 .C_ON=1'b0;
    defparam \c0.i15_3_lut_4_lut_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_3_lut_4_lut_LC_20_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_3_lut_4_lut_LC_20_12_5  (
            .in0(N__57667),
            .in1(N__57683),
            .in2(N__56009),
            .in3(N__60957),
            .lcout(\c0.n38_adj_4448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1411_LC_20_12_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1411_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1411_LC_20_12_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i13_4_lut_adj_1411_LC_20_12_6  (
            .in0(N__64986),
            .in1(N__70443),
            .in2(N__70787),
            .in3(N__57822),
            .lcout(\c0.n36_adj_4447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1414_LC_20_13_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1414_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1414_LC_20_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1414_LC_20_13_0  (
            .in0(N__57732),
            .in1(N__58162),
            .in2(N__58458),
            .in3(N__55368),
            .lcout(),
            .ltout(\c0.n41_adj_4452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_1416_LC_20_13_1 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_1416_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_1416_LC_20_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_adj_1416_LC_20_13_1  (
            .in0(N__55587),
            .in1(N__55593),
            .in2(N__55635),
            .in3(N__57966),
            .lcout(\c0.n24540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1415_LC_20_13_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1415_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1415_LC_20_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1415_LC_20_13_2  (
            .in0(N__60416),
            .in1(N__55631),
            .in2(N__70677),
            .in3(N__59366),
            .lcout(\c0.n39_adj_4453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1413_LC_20_13_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1413_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1413_LC_20_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1413_LC_20_13_3  (
            .in0(N__58051),
            .in1(N__70854),
            .in2(N__64059),
            .in3(N__57801),
            .lcout(\c0.n40_adj_4451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_4_lut_adj_1606_LC_20_13_4 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_4_lut_adj_1606_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_4_lut_adj_1606_LC_20_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_2_lut_3_lut_4_lut_adj_1606_LC_20_13_4  (
            .in0(N__71114),
            .in1(N__69585),
            .in2(N__60427),
            .in3(N__58053),
            .lcout(\c0.n22_adj_4244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1673_LC_20_13_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1673_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1673_LC_20_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1673_LC_20_13_5  (
            .in0(N__58049),
            .in1(N__60414),
            .in2(_gnd_net_),
            .in3(N__71113),
            .lcout(\c0.n23178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_adj_1828_LC_20_13_6 .C_ON=1'b0;
    defparam \c0.i7_2_lut_adj_1828_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_adj_1828_LC_20_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i7_2_lut_adj_1828_LC_20_13_6  (
            .in0(N__60415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58050),
            .lcout(\c0.n31_adj_4701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_LC_20_13_7 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_LC_20_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_3_lut_4_lut_LC_20_13_7  (
            .in0(N__58052),
            .in1(N__60417),
            .in2(N__65040),
            .in3(N__71115),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1847_LC_20_14_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1847_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1847_LC_20_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1847_LC_20_14_0  (
            .in0(N__61334),
            .in1(N__55760),
            .in2(N__55581),
            .in3(N__55565),
            .lcout(\c0.n13721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1599_LC_20_14_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1599_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1599_LC_20_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1599_LC_20_14_1  (
            .in0(N__55533),
            .in1(N__55524),
            .in2(N__55482),
            .in3(N__55454),
            .lcout(\c0.n23611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i85_LC_20_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i85_LC_20_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i85_LC_20_14_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i85_LC_20_14_2  (
            .in0(N__71936),
            .in1(N__69195),
            .in2(N__55779),
            .in3(N__73610),
            .lcout(\c0.data_in_frame_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1741_LC_20_14_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1741_LC_20_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1741_LC_20_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1741_LC_20_14_3  (
            .in0(_gnd_net_),
            .in1(N__55797),
            .in2(_gnd_net_),
            .in3(N__60413),
            .lcout(\c0.n8_adj_4673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i68_LC_20_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i68_LC_20_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i68_LC_20_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i68_LC_20_14_4  (
            .in0(N__72898),
            .in1(N__73608),
            .in2(N__72309),
            .in3(N__77123),
            .lcout(\c0.data_in_frame_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i84_LC_20_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i84_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i84_LC_20_14_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i84_LC_20_14_5  (
            .in0(N__69194),
            .in1(N__77122),
            .in2(N__73684),
            .in3(N__55972),
            .lcout(\c0.data_in_frame_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i69_LC_20_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i69_LC_20_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i69_LC_20_14_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i69_LC_20_14_6  (
            .in0(N__71937),
            .in1(N__73609),
            .in2(N__76047),
            .in3(N__72899),
            .lcout(\c0.data_in_frame_8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_20_14_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_20_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_LC_20_14_7  (
            .in0(N__72283),
            .in1(N__55775),
            .in2(_gnd_net_),
            .in3(N__55882),
            .lcout(\c0.n22455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_4_lut_LC_20_15_0 .C_ON=1'b0;
    defparam \c0.i29_4_lut_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i29_4_lut_LC_20_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i29_4_lut_LC_20_15_0  (
            .in0(N__55740),
            .in1(N__55686),
            .in2(N__74964),
            .in3(N__55653),
            .lcout(\c0.n65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i77_LC_20_15_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i77_LC_20_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i77_LC_20_15_2 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i77_LC_20_15_2  (
            .in0(N__71875),
            .in1(N__61245),
            .in2(N__73685),
            .in3(N__74180),
            .lcout(\c0.data_in_frame_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i46_4_lut_LC_20_15_3 .C_ON=1'b0;
    defparam \c0.i46_4_lut_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i46_4_lut_LC_20_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i46_4_lut_LC_20_15_3  (
            .in0(N__77446),
            .in1(N__55931),
            .in2(N__72006),
            .in3(N__55944),
            .lcout(\c0.n127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1805_LC_20_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1805_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1805_LC_20_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1805_LC_20_15_4  (
            .in0(_gnd_net_),
            .in1(N__58136),
            .in2(_gnd_net_),
            .in3(N__58097),
            .lcout(\c0.n5_adj_4311 ),
            .ltout(\c0.n5_adj_4311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_4_lut_adj_1357_LC_20_15_5 .C_ON=1'b0;
    defparam \c0.i29_4_lut_adj_1357_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i29_4_lut_adj_1357_LC_20_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i29_4_lut_adj_1357_LC_20_15_5  (
            .in0(N__70885),
            .in1(N__61235),
            .in2(N__55983),
            .in3(N__55965),
            .lcout(\c0.n85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1785_LC_20_15_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1785_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1785_LC_20_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1785_LC_20_15_6  (
            .in0(N__55943),
            .in1(N__65010),
            .in2(N__55932),
            .in3(N__58767),
            .lcout(\c0.n22644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i67_LC_20_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i67_LC_20_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i67_LC_20_15_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i67_LC_20_15_7  (
            .in0(N__72935),
            .in1(N__73611),
            .in2(N__55898),
            .in3(N__79110),
            .lcout(\c0.data_in_frame_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i39_2_lut_LC_20_16_0 .C_ON=1'b0;
    defparam \c0.i39_2_lut_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i39_2_lut_LC_20_16_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i39_2_lut_LC_20_16_0  (
            .in0(N__62528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62666),
            .lcout(),
            .ltout(\c0.n120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i71_4_lut_LC_20_16_1 .C_ON=1'b0;
    defparam \c0.i71_4_lut_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i71_4_lut_LC_20_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i71_4_lut_LC_20_16_1  (
            .in0(N__61890),
            .in1(N__62638),
            .in2(N__55866),
            .in3(N__55863),
            .lcout(),
            .ltout(\c0.n152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i79_4_lut_LC_20_16_2 .C_ON=1'b0;
    defparam \c0.i79_4_lut_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i79_4_lut_LC_20_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i79_4_lut_LC_20_16_2  (
            .in0(N__69760),
            .in1(N__58554),
            .in2(N__55851),
            .in3(N__55848),
            .lcout(\c0.n160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_4_lut_LC_20_16_3 .C_ON=1'b0;
    defparam \c0.i11_3_lut_4_lut_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_4_lut_LC_20_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_3_lut_4_lut_LC_20_16_3  (
            .in0(N__64340),
            .in1(N__70297),
            .in2(N__70449),
            .in3(N__55838),
            .lcout(),
            .ltout(\c0.n30_adj_4571_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1573_LC_20_16_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1573_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1573_LC_20_16_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i15_4_lut_adj_1573_LC_20_16_4  (
            .in0(N__58966),
            .in1(N__55824),
            .in2(N__55803),
            .in3(N__69804),
            .lcout(),
            .ltout(\c0.n34_adj_4600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1574_LC_20_16_5 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1574_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1574_LC_20_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1574_LC_20_16_5  (
            .in0(N__56112),
            .in1(N__69759),
            .in2(N__56103),
            .in3(N__56100),
            .lcout(\c0.n24333 ),
            .ltout(\c0.n24333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1698_LC_20_16_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1698_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1698_LC_20_16_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1698_LC_20_16_6  (
            .in0(N__62527),
            .in1(_gnd_net_),
            .in2(N__56088),
            .in3(N__62476),
            .lcout(\c0.n23661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1396_LC_20_17_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1396_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1396_LC_20_17_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1396_LC_20_17_0  (
            .in0(N__56038),
            .in1(N__72001),
            .in2(N__56073),
            .in3(N__65927),
            .lcout(\c0.n22173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i132_LC_20_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i132_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i132_LC_20_17_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i132_LC_20_17_1  (
            .in0(N__72965),
            .in1(N__80262),
            .in2(N__77098),
            .in3(N__56039),
            .lcout(\c0.data_in_frame_16_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i139_LC_20_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i139_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i139_LC_20_17_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i139_LC_20_17_2  (
            .in0(N__80259),
            .in1(N__74146),
            .in2(N__79182),
            .in3(N__58669),
            .lcout(\c0.data_in_frame_17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i131_LC_20_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i131_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i131_LC_20_17_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i131_LC_20_17_3  (
            .in0(N__72964),
            .in1(N__80261),
            .in2(N__65960),
            .in3(N__79140),
            .lcout(\c0.data_in_frame_16_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i158_LC_20_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i158_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i158_LC_20_17_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i158_LC_20_17_4  (
            .in0(N__80260),
            .in1(N__76611),
            .in2(N__71635),
            .in3(N__79784),
            .lcout(\c0.data_in_frame_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i156_LC_20_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i156_LC_20_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i156_LC_20_17_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i156_LC_20_17_5  (
            .in0(N__76610),
            .in1(N__80263),
            .in2(N__77099),
            .in3(N__59129),
            .lcout(\c0.data_in_frame_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1588_LC_20_17_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1588_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1588_LC_20_17_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1588_LC_20_17_6  (
            .in0(N__72002),
            .in1(N__62667),
            .in2(_gnd_net_),
            .in3(N__60048),
            .lcout(\c0.n22540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i80_4_lut_LC_20_17_7 .C_ON=1'b0;
    defparam \c0.i80_4_lut_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i80_4_lut_LC_20_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i80_4_lut_LC_20_17_7  (
            .in0(N__56022),
            .in1(N__58560),
            .in2(N__61212),
            .in3(N__56247),
            .lcout(\c0.n24520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1866_LC_20_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1866_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1866_LC_20_18_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1866_LC_20_18_0  (
            .in0(N__56240),
            .in1(N__61429),
            .in2(_gnd_net_),
            .in3(N__62294),
            .lcout(\c0.n22104 ),
            .ltout(\c0.n22104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i141_LC_20_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i141_LC_20_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i141_LC_20_18_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i141_LC_20_18_1  (
            .in0(N__74207),
            .in1(N__71958),
            .in2(N__56196),
            .in3(N__72238),
            .lcout(\c0.data_in_frame_17_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i140_LC_20_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i140_LC_20_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i140_LC_20_18_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i140_LC_20_18_2  (
            .in0(N__77100),
            .in1(N__74208),
            .in2(N__58829),
            .in3(N__80264),
            .lcout(\c0.data_in_frame_17_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1176_LC_20_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1176_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1176_LC_20_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1176_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(N__72237),
            .in2(_gnd_net_),
            .in3(N__58821),
            .lcout(\c0.n22822 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1708_LC_20_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1708_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1708_LC_20_18_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1708_LC_20_18_4  (
            .in0(N__77639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77579),
            .lcout(),
            .ltout(\c0.n22347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1311_LC_20_18_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1311_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1311_LC_20_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1311_LC_20_18_5  (
            .in0(N__56192),
            .in1(N__59125),
            .in2(N__56166),
            .in3(N__56159),
            .lcout(\c0.n10_adj_4315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_3_lut_adj_2043_LC_20_18_6 .C_ON=1'b0;
    defparam \c0.i13_2_lut_3_lut_adj_2043_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_3_lut_adj_2043_LC_20_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i13_2_lut_3_lut_adj_2043_LC_20_18_6  (
            .in0(N__56147),
            .in1(N__59730),
            .in2(_gnd_net_),
            .in3(N__75784),
            .lcout(\c0.n39_adj_4341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1204_LC_20_18_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1204_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1204_LC_20_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1204_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(N__63141),
            .in2(_gnd_net_),
            .in3(N__72299),
            .lcout(\c0.n10_adj_4230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_3_lut_4_lut_LC_20_19_0 .C_ON=1'b0;
    defparam \c0.i21_3_lut_4_lut_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21_3_lut_4_lut_LC_20_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_3_lut_4_lut_LC_20_19_0  (
            .in0(N__67376),
            .in1(N__67362),
            .in2(N__67415),
            .in3(N__59433),
            .lcout(\c0.n45_adj_4476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_LC_20_19_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_LC_20_19_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i6_2_lut_3_lut_LC_20_19_1  (
            .in0(N__59280),
            .in1(N__58715),
            .in2(_gnd_net_),
            .in3(N__58843),
            .lcout(\c0.n14_adj_4356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_4_lut_LC_20_19_2 .C_ON=1'b0;
    defparam \c0.i7_2_lut_4_lut_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_4_lut_LC_20_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_2_lut_4_lut_LC_20_19_2  (
            .in0(N__59333),
            .in1(N__62682),
            .in2(N__58848),
            .in3(N__60062),
            .lcout(\c0.n22_adj_4350 ),
            .ltout(\c0.n22_adj_4350_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_3_lut_LC_20_19_3 .C_ON=1'b0;
    defparam \c0.i25_3_lut_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i25_3_lut_LC_20_19_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i25_3_lut_LC_20_19_3  (
            .in0(N__59281),
            .in1(_gnd_net_),
            .in2(N__56418),
            .in3(N__56324),
            .lcout(\c0.n59_adj_4351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_adj_1991_LC_20_19_4 .C_ON=1'b0;
    defparam \c0.i8_2_lut_adj_1991_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_adj_1991_LC_20_19_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i8_2_lut_adj_1991_LC_20_19_4  (
            .in0(N__58847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59282),
            .lcout(\c0.n11_adj_4505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_LC_20_19_5 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_LC_20_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_2_lut_3_lut_LC_20_19_5  (
            .in0(N__56415),
            .in1(N__56373),
            .in2(_gnd_net_),
            .in3(N__56325),
            .lcout(\c0.n28_adj_4504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i104_LC_20_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i104_LC_20_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i104_LC_20_19_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i104_LC_20_19_6  (
            .in0(N__73598),
            .in1(N__80044),
            .in2(N__76275),
            .in3(N__63148),
            .lcout(\c0.data_in_frame_12_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_adj_1951_LC_20_19_7 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_adj_1951_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_adj_1951_LC_20_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_adj_1951_LC_20_19_7  (
            .in0(N__59348),
            .in1(N__58500),
            .in2(N__58671),
            .in3(N__81058),
            .lcout(\c0.n20_adj_4596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1473_LC_20_20_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1473_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1473_LC_20_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1473_LC_20_20_0  (
            .in0(N__75795),
            .in1(N__56610),
            .in2(N__56298),
            .in3(N__56280),
            .lcout(\c0.n23975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1994_LC_20_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1994_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1994_LC_20_20_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1994_LC_20_20_1  (
            .in0(N__74679),
            .in1(N__74529),
            .in2(N__74387),
            .in3(N__73597),
            .lcout(n22118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1746_LC_20_20_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1746_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1746_LC_20_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1746_LC_20_20_2  (
            .in0(N__56573),
            .in1(N__56595),
            .in2(N__70818),
            .in3(N__66709),
            .lcout(\c0.n9_adj_4521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1568_LC_20_20_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1568_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1568_LC_20_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1568_LC_20_20_3  (
            .in0(N__56493),
            .in1(N__56604),
            .in2(N__81114),
            .in3(N__59031),
            .lcout(\c0.n23733 ),
            .ltout(\c0.n23733_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1591_LC_20_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1591_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1591_LC_20_20_4 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_1591_LC_20_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56598),
            .in3(N__56594),
            .lcout(\c0.n20314 ),
            .ltout(\c0.n20314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1512_LC_20_20_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1512_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1512_LC_20_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1512_LC_20_20_5  (
            .in0(N__56894),
            .in1(N__56572),
            .in2(N__56529),
            .in3(N__56858),
            .lcout(\c0.n13_adj_4492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1424_LC_20_20_6 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1424_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1424_LC_20_20_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_1424_LC_20_20_6  (
            .in0(N__74817),
            .in1(N__56526),
            .in2(N__59636),
            .in3(N__56499),
            .lcout(\c0.n37_adj_4458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_4_lut_adj_1702_LC_20_21_0 .C_ON=1'b0;
    defparam \c0.i9_3_lut_4_lut_adj_1702_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_4_lut_adj_1702_LC_20_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_3_lut_4_lut_adj_1702_LC_20_21_0  (
            .in0(N__72321),
            .in1(N__77872),
            .in2(N__73401),
            .in3(N__77816),
            .lcout(\c0.n22_adj_4597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i105_LC_20_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i105_LC_20_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i105_LC_20_21_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i105_LC_20_21_1  (
            .in0(N__75493),
            .in1(N__75421),
            .in2(N__58304),
            .in3(N__80615),
            .lcout(\c0.data_in_frame_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i233_LC_20_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i233_LC_20_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i233_LC_20_21_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i233_LC_20_21_2  (
            .in0(N__75420),
            .in1(N__56483),
            .in2(N__80673),
            .in3(N__56684),
            .lcout(\c0.data_in_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i240_LC_20_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i240_LC_20_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i240_LC_20_21_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i240_LC_20_21_3  (
            .in0(N__56482),
            .in1(N__76227),
            .in2(N__75426),
            .in3(N__56904),
            .lcout(\c0.data_in_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1429_LC_20_21_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1429_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1429_LC_20_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1429_LC_20_21_4  (
            .in0(N__56903),
            .in1(N__56895),
            .in2(_gnd_net_),
            .in3(N__56862),
            .lcout(\c0.n12_adj_4466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1745_LC_20_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1745_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1745_LC_20_21_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1745_LC_20_21_5  (
            .in0(N__56817),
            .in1(N__77287),
            .in2(_gnd_net_),
            .in3(N__59561),
            .lcout(),
            .ltout(\c0.n11_adj_4474_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1433_LC_20_21_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1433_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1433_LC_20_21_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1433_LC_20_21_6  (
            .in0(N__56766),
            .in1(N__63226),
            .in2(N__56760),
            .in3(N__56757),
            .lcout(\c0.n18_adj_4475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i112_LC_20_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i112_LC_20_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i112_LC_20_21_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i112_LC_20_21_7  (
            .in0(N__75494),
            .in1(N__75422),
            .in2(N__62847),
            .in3(N__76228),
            .lcout(\c0.data_in_frame_13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1455_LC_20_22_0 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1455_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1455_LC_20_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1455_LC_20_22_0  (
            .in0(N__58719),
            .in1(N__64134),
            .in2(N__56712),
            .in3(N__56691),
            .lcout(\c0.n44_adj_4501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_324_2_lut_3_lut_LC_20_22_1 .C_ON=1'b0;
    defparam \c0.i1_rep_324_2_lut_3_lut_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_324_2_lut_3_lut_LC_20_22_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_rep_324_2_lut_3_lut_LC_20_22_1  (
            .in0(N__56652),
            .in1(_gnd_net_),
            .in2(N__67152),
            .in3(N__57014),
            .lcout(\c0.n25446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1748_LC_20_22_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1748_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1748_LC_20_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1748_LC_20_22_2  (
            .in0(N__57015),
            .in1(N__67147),
            .in2(N__56685),
            .in3(N__56650),
            .lcout(),
            .ltout(\c0.n43_adj_4463_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_4_lut_adj_1426_LC_20_22_3 .C_ON=1'b0;
    defparam \c0.i32_4_lut_adj_1426_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i32_4_lut_adj_1426_LC_20_22_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i32_4_lut_adj_1426_LC_20_22_3  (
            .in0(N__76742),
            .in1(N__56669),
            .in2(N__56655),
            .in3(N__63786),
            .lcout(\c0.n74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_adj_1744_LC_20_22_4 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_adj_1744_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_adj_1744_LC_20_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_adj_1744_LC_20_22_4  (
            .in0(N__57016),
            .in1(N__67148),
            .in2(N__67327),
            .in3(N__56651),
            .lcout(\c0.n42_adj_4540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1234_LC_20_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1234_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1234_LC_20_22_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1234_LC_20_22_5  (
            .in0(N__67149),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57017),
            .lcout(\c0.n13911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_4_lut_adj_1505_LC_20_22_6 .C_ON=1'b0;
    defparam \c0.i33_4_lut_adj_1505_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i33_4_lut_adj_1505_LC_20_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i33_4_lut_adj_1505_LC_20_22_6  (
            .in0(N__63264),
            .in1(N__56973),
            .in2(N__59796),
            .in3(N__59808),
            .lcout(),
            .ltout(\c0.n23921_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1508_LC_20_22_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1508_LC_20_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1508_LC_20_22_7 .LUT_INIT=16'b1001111101101111;
    LogicCell40 \c0.i3_4_lut_adj_1508_LC_20_22_7  (
            .in0(N__56964),
            .in1(N__56955),
            .in2(N__56949),
            .in3(N__57113),
            .lcout(\c0.n21_adj_4547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_2_lut_4_lut_adj_1732_LC_20_23_0 .C_ON=1'b0;
    defparam \c0.i10_2_lut_4_lut_adj_1732_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_2_lut_4_lut_adj_1732_LC_20_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_2_lut_4_lut_adj_1732_LC_20_23_0  (
            .in0(N__67559),
            .in1(N__68366),
            .in2(N__75938),
            .in3(N__68280),
            .lcout(\c0.n31_adj_4542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1493_LC_20_23_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1493_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1493_LC_20_23_1 .LUT_INIT=16'b1111111110110111;
    LogicCell40 \c0.i14_4_lut_adj_1493_LC_20_23_1  (
            .in0(N__66768),
            .in1(N__56934),
            .in2(N__68295),
            .in3(N__57120),
            .lcout(\c0.n32_adj_4533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i210_LC_20_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i210_LC_20_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i210_LC_20_23_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i210_LC_20_23_2  (
            .in0(N__69204),
            .in1(N__75138),
            .in2(N__63731),
            .in3(N__79457),
            .lcout(\c0.data_in_frame_26_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i40_4_lut_adj_1468_LC_20_23_3 .C_ON=1'b0;
    defparam \c0.i40_4_lut_adj_1468_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i40_4_lut_adj_1468_LC_20_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i40_4_lut_adj_1468_LC_20_23_3  (
            .in0(N__63263),
            .in1(N__56910),
            .in2(N__75636),
            .in3(N__59505),
            .lcout(\c0.n82_adj_4517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i194_LC_20_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i194_LC_20_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i194_LC_20_23_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i194_LC_20_23_4  (
            .in0(N__72989),
            .in1(N__75137),
            .in2(N__64179),
            .in3(N__79456),
            .lcout(\c0.data_in_frame_24_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1494_LC_20_23_7 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1494_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1494_LC_20_23_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i11_3_lut_adj_1494_LC_20_23_7  (
            .in0(N__67297),
            .in1(N__77341),
            .in2(_gnd_net_),
            .in3(N__66831),
            .lcout(\c0.n32_adj_4534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_3_lut_LC_20_24_0 .C_ON=1'b0;
    defparam \c0.i29_3_lut_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i29_3_lut_LC_20_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i29_3_lut_LC_20_24_0  (
            .in0(N__64085),
            .in1(N__59782),
            .in2(_gnd_net_),
            .in3(N__59896),
            .lcout(),
            .ltout(\c0.n71_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i39_4_lut_LC_20_24_1 .C_ON=1'b0;
    defparam \c0.i39_4_lut_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i39_4_lut_LC_20_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i39_4_lut_LC_20_24_1  (
            .in0(N__57174),
            .in1(N__67033),
            .in2(N__57162),
            .in3(N__59985),
            .lcout(),
            .ltout(\c0.n81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1480_LC_20_24_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1480_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1480_LC_20_24_2 .LUT_INIT=16'b1110111111111110;
    LogicCell40 \c0.i10_4_lut_adj_1480_LC_20_24_2  (
            .in0(N__57155),
            .in1(N__59955),
            .in2(N__57129),
            .in3(N__57126),
            .lcout(\c0.n28_adj_4523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1492_LC_20_24_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1492_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1492_LC_20_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1492_LC_20_24_3  (
            .in0(N__57114),
            .in1(N__57080),
            .in2(_gnd_net_),
            .in3(N__67506),
            .lcout(),
            .ltout(\c0.n23_adj_4532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1495_LC_20_24_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1495_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1495_LC_20_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1495_LC_20_24_4  (
            .in0(N__67797),
            .in1(N__77898),
            .in2(N__57048),
            .in3(N__67819),
            .lcout(),
            .ltout(\c0.n38_adj_4535_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_1502_LC_20_24_5 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_1502_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_1502_LC_20_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_1502_LC_20_24_5  (
            .in0(N__67748),
            .in1(N__57045),
            .in2(N__57039),
            .in3(N__57036),
            .lcout(\c0.n15_adj_4497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1978_LC_20_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1978_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1978_LC_20_25_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_1978_LC_20_25_7  (
            .in0(_gnd_net_),
            .in1(N__61380),
            .in2(_gnd_net_),
            .in3(N__62318),
            .lcout(\c0.n12_adj_4672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1833_LC_21_6_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1833_LC_21_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1833_LC_21_6_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1833_LC_21_6_2  (
            .in0(_gnd_net_),
            .in1(N__69354),
            .in2(_gnd_net_),
            .in3(N__64531),
            .lcout(\c0.n13998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_1767_LC_21_7_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_1767_LC_21_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_1767_LC_21_7_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i3_3_lut_adj_1767_LC_21_7_0  (
            .in0(N__60594),
            .in1(N__60204),
            .in2(_gnd_net_),
            .in3(N__68120),
            .lcout(\c0.n8_adj_4677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i79_LC_21_7_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i79_LC_21_7_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i79_LC_21_7_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i79_LC_21_7_2  (
            .in0(N__73717),
            .in1(N__74150),
            .in2(N__57417),
            .in3(N__73291),
            .lcout(\c0.data_in_frame_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_21_7_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_21_7_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_21_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i44_LC_21_7_3  (
            .in0(N__77106),
            .in1(N__69462),
            .in2(_gnd_net_),
            .in3(N__57366),
            .lcout(data_in_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i87_LC_21_7_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i87_LC_21_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i87_LC_21_7_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i87_LC_21_7_4  (
            .in0(N__73718),
            .in1(N__69185),
            .in2(N__61781),
            .in3(N__73292),
            .lcout(\c0.data_in_frame_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_21_7_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_21_7_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_21_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i43_LC_21_7_5  (
            .in0(N__57324),
            .in1(N__69461),
            .in2(_gnd_net_),
            .in3(N__79106),
            .lcout(data_in_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1582_LC_21_7_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1582_LC_21_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1582_LC_21_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1582_LC_21_7_7  (
            .in0(_gnd_net_),
            .in1(N__64049),
            .in2(_gnd_net_),
            .in3(N__69330),
            .lcout(\c0.n7_adj_4603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1609_LC_21_8_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1609_LC_21_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1609_LC_21_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1609_LC_21_8_0  (
            .in0(N__61044),
            .in1(N__57192),
            .in2(N__57309),
            .in3(N__57245),
            .lcout(\c0.n23554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_21_8_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_21_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_21_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i45_LC_21_8_1  (
            .in0(N__57461),
            .in1(N__71968),
            .in2(_gnd_net_),
            .in3(N__69459),
            .lcout(data_in_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78806),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1608_LC_21_8_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1608_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1608_LC_21_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1608_LC_21_8_2  (
            .in0(N__57951),
            .in1(N__60634),
            .in2(N__57447),
            .in3(N__60203),
            .lcout(\c0.n12_adj_4612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_4_lut_adj_1662_LC_21_8_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_4_lut_adj_1662_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_4_lut_adj_1662_LC_21_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_4_lut_adj_1662_LC_21_8_3  (
            .in0(N__68928),
            .in1(N__64490),
            .in2(N__72585),
            .in3(N__69584),
            .lcout(\c0.n15_adj_4444 ),
            .ltout(\c0.n15_adj_4444_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i46_4_lut_adj_1407_LC_21_8_4 .C_ON=1'b0;
    defparam \c0.i46_4_lut_adj_1407_LC_21_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i46_4_lut_adj_1407_LC_21_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i46_4_lut_adj_1407_LC_21_8_4  (
            .in0(N__61466),
            .in1(N__57428),
            .in2(N__57510),
            .in3(N__69492),
            .lcout(\c0.n102_adj_4445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_1672_LC_21_8_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_1672_LC_21_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_1672_LC_21_8_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_1672_LC_21_8_5  (
            .in0(N__60632),
            .in1(_gnd_net_),
            .in2(N__57462),
            .in3(N__57494),
            .lcout(\c0.n11_adj_4656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1668_LC_21_8_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1668_LC_21_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1668_LC_21_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1668_LC_21_8_6  (
            .in0(N__57495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57460),
            .lcout(\c0.n6_adj_4611 ),
            .ltout(\c0.n6_adj_4611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i35_2_lut_4_lut_LC_21_8_7 .C_ON=1'b0;
    defparam \c0.i35_2_lut_4_lut_LC_21_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i35_2_lut_4_lut_LC_21_8_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i35_2_lut_4_lut_LC_21_8_7  (
            .in0(N__60633),
            .in1(N__57950),
            .in2(N__57438),
            .in3(N__61043),
            .lcout(\c0.n91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i57_LC_21_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i57_LC_21_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i57_LC_21_9_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i57_LC_21_9_0  (
            .in0(N__80922),
            .in1(N__70166),
            .in2(N__64502),
            .in3(N__80737),
            .lcout(\c0.data_in_frame_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_21_9_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_21_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_21_9_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i7_LC_21_9_1  (
            .in0(N__70165),
            .in1(N__73294),
            .in2(N__60648),
            .in3(N__72924),
            .lcout(\c0.data_in_frame_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_21_9_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_21_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_21_9_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i23_LC_21_9_2  (
            .in0(N__73293),
            .in1(N__70167),
            .in2(N__60746),
            .in3(N__69150),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1631_LC_21_9_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1631_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1631_LC_21_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1631_LC_21_9_3  (
            .in0(N__60283),
            .in1(N__60737),
            .in2(_gnd_net_),
            .in3(N__68495),
            .lcout(\c0.n23302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_21_9_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_21_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_21_9_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i5_LC_21_9_4  (
            .in0(N__68496),
            .in1(N__71959),
            .in2(N__72966),
            .in3(N__70022),
            .lcout(\c0.data_in_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i165_LC_21_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i165_LC_21_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i165_LC_21_9_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i165_LC_21_9_5  (
            .in0(N__79986),
            .in1(N__59702),
            .in2(N__71969),
            .in3(N__80426),
            .lcout(\c0.data_in_frame_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_21_9_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_21_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_21_9_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i6_LC_21_9_6  (
            .in0(N__60301),
            .in1(N__79646),
            .in2(N__72967),
            .in3(N__70023),
            .lcout(\c0.data_in_frame_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_21_9_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_21_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_21_9_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i4_LC_21_9_7  (
            .in0(N__70164),
            .in1(N__77111),
            .in2(N__68121),
            .in3(N__72923),
            .lcout(\c0.data_in_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1898_LC_21_10_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1898_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1898_LC_21_10_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_adj_1898_LC_21_10_0  (
            .in0(N__67915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68096),
            .lcout(\c0.n10_adj_4722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1873_LC_21_10_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1873_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1873_LC_21_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1873_LC_21_10_2  (
            .in0(_gnd_net_),
            .in1(N__65678),
            .in2(_gnd_net_),
            .in3(N__57957),
            .lcout(\c0.n15_adj_4450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_21_10_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_21_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_21_10_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i22_LC_21_10_3  (
            .in0(N__69156),
            .in1(N__70141),
            .in2(N__67943),
            .in3(N__79589),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1595_LC_21_10_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1595_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1595_LC_21_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1595_LC_21_10_4  (
            .in0(N__67914),
            .in1(N__68497),
            .in2(_gnd_net_),
            .in3(N__68095),
            .lcout(\c0.n13453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_21_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_21_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_21_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_21_10_5  (
            .in0(N__75186),
            .in1(N__68437),
            .in2(_gnd_net_),
            .in3(N__58128),
            .lcout(data_in_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i164_LC_21_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i164_LC_21_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i164_LC_21_10_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i164_LC_21_10_6  (
            .in0(N__79953),
            .in1(N__80425),
            .in2(N__75765),
            .in3(N__77130),
            .lcout(\c0.data_in_frame_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_2_lut_4_lut_LC_21_10_7 .C_ON=1'b0;
    defparam \c0.i25_2_lut_4_lut_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i25_2_lut_4_lut_LC_21_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_2_lut_4_lut_LC_21_10_7  (
            .in0(N__57536),
            .in1(N__64827),
            .in2(N__64902),
            .in3(N__64779),
            .lcout(\c0.n61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_1233_LC_21_11_0 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_1233_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_1233_LC_21_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_1233_LC_21_11_0  (
            .in0(_gnd_net_),
            .in1(N__60884),
            .in2(_gnd_net_),
            .in3(N__62070),
            .lcout(\c0.n17_adj_4224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i54_4_lut_LC_21_11_1 .C_ON=1'b0;
    defparam \c0.i54_4_lut_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i54_4_lut_LC_21_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i54_4_lut_LC_21_11_1  (
            .in0(N__57864),
            .in1(N__57855),
            .in2(N__61503),
            .in3(N__57849),
            .lcout(),
            .ltout(\c0.n110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i55_4_lut_LC_21_11_2 .C_ON=1'b0;
    defparam \c0.i55_4_lut_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i55_4_lut_LC_21_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i55_4_lut_LC_21_11_2  (
            .in0(N__57843),
            .in1(N__57837),
            .in2(N__57825),
            .in3(N__57738),
            .lcout(\c0.n24465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1621_LC_21_11_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1621_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1621_LC_21_11_3 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1621_LC_21_11_3  (
            .in0(N__62071),
            .in1(N__57730),
            .in2(N__60895),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_frame_0__7__N_2579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_2_lut_3_lut_4_lut_LC_21_11_4 .C_ON=1'b0;
    defparam \c0.i31_2_lut_3_lut_4_lut_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i31_2_lut_3_lut_4_lut_LC_21_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i31_2_lut_3_lut_4_lut_LC_21_11_4  (
            .in0(N__57728),
            .in1(N__58155),
            .in2(N__57800),
            .in3(N__60942),
            .lcout(\c0.n87 ),
            .ltout(\c0.n87_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i50_4_lut_adj_1410_LC_21_11_5 .C_ON=1'b0;
    defparam \c0.i50_4_lut_adj_1410_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i50_4_lut_adj_1410_LC_21_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i50_4_lut_adj_1410_LC_21_11_5  (
            .in0(N__57765),
            .in1(N__57753),
            .in2(N__57741),
            .in3(N__64389),
            .lcout(\c0.n106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1780_LC_21_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1780_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1780_LC_21_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1780_LC_21_11_6  (
            .in0(N__57729),
            .in1(N__60883),
            .in2(N__61596),
            .in3(N__62069),
            .lcout(\c0.n7_adj_4304 ),
            .ltout(\c0.n7_adj_4304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1283_LC_21_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1283_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1283_LC_21_11_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1283_LC_21_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57675),
            .in3(N__57661),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1902_LC_21_12_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1902_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1902_LC_21_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1902_LC_21_12_0  (
            .in0(N__58048),
            .in1(N__57606),
            .in2(N__61083),
            .in3(N__71080),
            .lcout(\c0.n27_adj_4725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i49_3_lut_4_lut_LC_21_12_1 .C_ON=1'b0;
    defparam \c0.i49_3_lut_4_lut_LC_21_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i49_3_lut_4_lut_LC_21_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i49_3_lut_4_lut_LC_21_12_1  (
            .in0(N__72397),
            .in1(N__58253),
            .in2(N__72483),
            .in3(N__60029),
            .lcout(\c0.n130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1863_LC_21_12_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1863_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1863_LC_21_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1863_LC_21_12_2  (
            .in0(N__58230),
            .in1(N__58212),
            .in2(N__58200),
            .in3(N__65096),
            .lcout(\c0.n22_adj_4259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_LC_21_12_3 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_LC_21_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_LC_21_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_2_lut_3_lut_LC_21_12_3  (
            .in0(N__65706),
            .in1(_gnd_net_),
            .in2(N__60953),
            .in3(N__57960),
            .lcout(\c0.n18_adj_4314 ),
            .ltout(\c0.n18_adj_4314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_4_lut_adj_1678_LC_21_12_4 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_4_lut_adj_1678_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_4_lut_adj_1678_LC_21_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_2_lut_3_lut_4_lut_adj_1678_LC_21_12_4  (
            .in0(N__71095),
            .in1(N__58132),
            .in2(N__58101),
            .in3(N__58098),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_1895_LC_21_12_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_1895_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_1895_LC_21_12_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i3_2_lut_adj_1895_LC_21_12_5  (
            .in0(N__71079),
            .in1(N__58047),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n22230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1412_LC_21_12_6 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1412_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1412_LC_21_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1412_LC_21_12_6  (
            .in0(N__70225),
            .in1(N__64345),
            .in2(N__65295),
            .in3(N__57972),
            .lcout(\c0.n42_adj_4449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_4_lut_4_lut_LC_21_12_7 .C_ON=1'b0;
    defparam \c0.i9_3_lut_4_lut_4_lut_LC_21_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_4_lut_4_lut_LC_21_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_3_lut_4_lut_4_lut_LC_21_12_7  (
            .in0(N__65705),
            .in1(N__71094),
            .in2(N__60952),
            .in3(N__57959),
            .lcout(\c0.n24_adj_4689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1377_LC_21_13_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1377_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1377_LC_21_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1377_LC_21_13_0  (
            .in0(N__78852),
            .in1(N__66863),
            .in2(N__73038),
            .in3(N__57888),
            .lcout(\c0.n41_adj_4360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2040_LC_21_13_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2040_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2040_LC_21_13_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_2040_LC_21_13_2  (
            .in0(N__58447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70439),
            .lcout(\c0.n31 ),
            .ltout(\c0.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_adj_1228_LC_21_13_3 .C_ON=1'b0;
    defparam \c0.i23_4_lut_adj_1228_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_adj_1228_LC_21_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_adj_1228_LC_21_13_3  (
            .in0(N__61293),
            .in1(N__58331),
            .in2(N__58410),
            .in3(N__58407),
            .lcout(\c0.n53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_21_13_4 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_21_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_LC_21_13_4  (
            .in0(N__58377),
            .in1(N__60558),
            .in2(N__58350),
            .in3(N__58341),
            .lcout(\c0.n23267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i115_LC_21_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i115_LC_21_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i115_LC_21_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i115_LC_21_13_5  (
            .in0(N__79168),
            .in1(N__59205),
            .in2(_gnd_net_),
            .in3(N__58332),
            .lcout(data_in_frame_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1747_LC_21_13_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1747_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1747_LC_21_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1747_LC_21_13_6  (
            .in0(N__58313),
            .in1(N__60557),
            .in2(N__58323),
            .in3(N__61292),
            .lcout(\c0.n23491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_21_13_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_21_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_21_13_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0__i51_LC_21_13_7  (
            .in0(N__68433),
            .in1(_gnd_net_),
            .in2(N__79193),
            .in3(N__58314),
            .lcout(data_in_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_21_14_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_21_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_21_14_0  (
            .in0(N__76037),
            .in1(N__77845),
            .in2(N__76070),
            .in3(N__81032),
            .lcout(\c0.n22205 ),
            .ltout(\c0.n22205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1696_LC_21_14_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1696_LC_21_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1696_LC_21_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1696_LC_21_14_1  (
            .in0(N__58305),
            .in1(N__60819),
            .in2(N__58284),
            .in3(N__58279),
            .lcout(\c0.n22589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_4_lut_LC_21_14_2 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_4_lut_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_4_lut_LC_21_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_2_lut_3_lut_4_lut_LC_21_14_2  (
            .in0(N__66053),
            .in1(N__77846),
            .in2(N__76048),
            .in3(N__77776),
            .lcout(\c0.n22_adj_4243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1652_LC_21_14_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1652_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1652_LC_21_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1652_LC_21_14_3  (
            .in0(N__72577),
            .in1(N__66052),
            .in2(_gnd_net_),
            .in3(N__69580),
            .lcout(\c0.n23598 ),
            .ltout(\c0.n23598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1723_LC_21_14_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1723_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1723_LC_21_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1723_LC_21_14_4  (
            .in0(_gnd_net_),
            .in1(N__77844),
            .in2(N__58503),
            .in3(N__81031),
            .lcout(\c0.n13128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_21_14_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_21_14_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_LC_21_14_5  (
            .in0(_gnd_net_),
            .in1(N__63032),
            .in2(_gnd_net_),
            .in3(N__72284),
            .lcout(\c0.n9_adj_4208 ),
            .ltout(\c0.n9_adj_4208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1890_LC_21_14_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1890_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1890_LC_21_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1890_LC_21_14_6  (
            .in0(N__73400),
            .in1(N__58496),
            .in2(N__58485),
            .in3(N__77777),
            .lcout(\c0.n22304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_LC_21_14_7 .C_ON=1'b0;
    defparam \c0.i26_4_lut_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_LC_21_14_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i26_4_lut_LC_21_14_7  (
            .in0(N__61122),
            .in1(N__68190),
            .in2(N__68879),
            .in3(N__62875),
            .lcout(\c0.n107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1883_LC_21_15_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1883_LC_21_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1883_LC_21_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1883_LC_21_15_0  (
            .in0(N__59260),
            .in1(N__59053),
            .in2(N__62615),
            .in3(N__58472),
            .lcout(\c0.n13892 ),
            .ltout(\c0.n13892_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1789_LC_21_15_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1789_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1789_LC_21_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1789_LC_21_15_1  (
            .in0(N__74714),
            .in1(N__66097),
            .in2(N__58461),
            .in3(N__58872),
            .lcout(\c0.n6215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1604_LC_21_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1604_LC_21_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1604_LC_21_15_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1604_LC_21_15_2  (
            .in0(N__61648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62808),
            .lcout(\c0.n22662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i95_LC_21_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i95_LC_21_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i95_LC_21_15_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i95_LC_21_15_3  (
            .in0(N__76654),
            .in1(N__73705),
            .in2(N__58451),
            .in3(N__73299),
            .lcout(\c0.data_in_frame_11_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1948_LC_21_15_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1948_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1948_LC_21_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1948_LC_21_15_4  (
            .in0(N__59352),
            .in1(N__59081),
            .in2(N__58670),
            .in3(N__58425),
            .lcout(\c0.n13797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1538_LC_21_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1538_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1538_LC_21_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1538_LC_21_15_5  (
            .in0(N__74713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58662),
            .lcout(\c0.n14088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1223_LC_21_15_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1223_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1223_LC_21_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1223_LC_21_15_6  (
            .in0(N__72631),
            .in1(N__72581),
            .in2(N__65748),
            .in3(N__65798),
            .lcout(\c0.n22547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1623_LC_21_16_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1623_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1623_LC_21_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1623_LC_21_16_2  (
            .in0(N__65112),
            .in1(N__70926),
            .in2(N__58638),
            .in3(N__65154),
            .lcout(\c0.n22825 ),
            .ltout(\c0.n22825_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1730_LC_21_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1730_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1730_LC_21_16_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1730_LC_21_16_3  (
            .in0(N__72165),
            .in1(_gnd_net_),
            .in2(N__58623),
            .in3(N__72210),
            .lcout(\c0.n22751 ),
            .ltout(\c0.n22751_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i68_4_lut_LC_21_16_4 .C_ON=1'b0;
    defparam \c0.i68_4_lut_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i68_4_lut_LC_21_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i68_4_lut_LC_21_16_4  (
            .in0(N__58620),
            .in1(N__58587),
            .in2(N__58572),
            .in3(N__58569),
            .lcout(\c0.n149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1632_LC_21_16_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1632_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1632_LC_21_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1632_LC_21_16_5  (
            .in0(N__65370),
            .in1(N__74962),
            .in2(_gnd_net_),
            .in3(N__61815),
            .lcout(\c0.n22586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i59_4_lut_LC_21_16_6 .C_ON=1'b0;
    defparam \c0.i59_4_lut_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i59_4_lut_LC_21_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i59_4_lut_LC_21_16_6  (
            .in0(N__65717),
            .in1(N__71116),
            .in2(N__65779),
            .in3(N__77792),
            .lcout(\c0.n140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1575_LC_21_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1575_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1575_LC_21_16_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1575_LC_21_16_7  (
            .in0(N__66096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66565),
            .lcout(\c0.n22843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1224_LC_21_17_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1224_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1224_LC_21_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1224_LC_21_17_0  (
            .in0(N__61796),
            .in1(N__63152),
            .in2(N__74718),
            .in3(N__61698),
            .lcout(\c0.n22_adj_4245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1279_LC_21_17_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1279_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1279_LC_21_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1279_LC_21_17_1  (
            .in0(N__66006),
            .in1(N__58700),
            .in2(_gnd_net_),
            .in3(N__72078),
            .lcout(\c0.n22514 ),
            .ltout(\c0.n22514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1871_LC_21_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1871_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1871_LC_21_17_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1871_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__58704),
            .in3(N__72103),
            .lcout(\c0.n22803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i129_LC_21_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i129_LC_21_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i129_LC_21_17_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i129_LC_21_17_3  (
            .in0(N__80746),
            .in1(N__72982),
            .in2(N__72110),
            .in3(N__80265),
            .lcout(\c0.data_in_frame_16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i130_LC_21_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i130_LC_21_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i130_LC_21_17_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i130_LC_21_17_4  (
            .in0(N__75253),
            .in1(N__58701),
            .in2(N__72992),
            .in3(N__80266),
            .lcout(\c0.data_in_frame_16_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i110_LC_21_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i110_LC_21_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i110_LC_21_17_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i110_LC_21_17_5  (
            .in0(N__79727),
            .in1(N__75499),
            .in2(N__66016),
            .in3(N__75373),
            .lcout(\c0.data_in_frame_13_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i111_LC_21_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i111_LC_21_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i111_LC_21_17_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i111_LC_21_17_6  (
            .in0(N__75498),
            .in1(N__73335),
            .in2(N__72088),
            .in3(N__75374),
            .lcout(\c0.data_in_frame_13_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1534_LC_21_17_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1534_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1534_LC_21_17_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i5_3_lut_adj_1534_LC_21_17_7  (
            .in0(N__73944),
            .in1(N__59724),
            .in2(_gnd_net_),
            .in3(N__66336),
            .lcout(\c0.n14_adj_4566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1729_LC_21_18_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1729_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1729_LC_21_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1729_LC_21_18_0  (
            .in0(N__58980),
            .in1(N__72681),
            .in2(N__58782),
            .in3(N__70549),
            .lcout(\c0.n14165 ),
            .ltout(\c0.n14165_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1521_LC_21_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1521_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1521_LC_21_18_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_1521_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__58674),
            .in3(N__62360),
            .lcout(\c0.n4_adj_4345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1681_LC_21_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1681_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1681_LC_21_18_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1681_LC_21_18_2  (
            .in0(N__58777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59025),
            .lcout(),
            .ltout(\c0.n4_adj_4658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1786_LC_21_18_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1786_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1786_LC_21_18_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1786_LC_21_18_3  (
            .in0(N__62407),
            .in1(N__62483),
            .in2(N__58983),
            .in3(N__58979),
            .lcout(),
            .ltout(\c0.n12_adj_4682_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1788_LC_21_18_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1788_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1788_LC_21_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1788_LC_21_18_4  (
            .in0(N__58938),
            .in1(N__58725),
            .in2(N__58902),
            .in3(N__58899),
            .lcout(\c0.n22249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1903_LC_21_18_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1903_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1903_LC_21_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1903_LC_21_18_5  (
            .in0(N__63430),
            .in1(N__63347),
            .in2(N__71631),
            .in3(N__58854),
            .lcout(\c0.n24534 ),
            .ltout(\c0.n24534_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1366_LC_21_18_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1366_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1366_LC_21_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1366_LC_21_18_6  (
            .in0(N__58828),
            .in1(N__58803),
            .in2(N__58797),
            .in3(N__62009),
            .lcout(\c0.n12_adj_4346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1618_LC_21_18_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1618_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1618_LC_21_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1618_LC_21_18_7  (
            .in0(N__70548),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58778),
            .lcout(\c0.n4_adj_4621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1561_LC_21_19_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1561_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1561_LC_21_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1561_LC_21_19_0  (
            .in0(N__77674),
            .in1(N__72123),
            .in2(N__77705),
            .in3(N__77812),
            .lcout(\c0.n44_adj_4588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_4_lut_LC_21_19_2 .C_ON=1'b0;
    defparam \c0.i9_2_lut_4_lut_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_4_lut_LC_21_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_2_lut_4_lut_LC_21_19_2  (
            .in0(N__60061),
            .in1(N__72347),
            .in2(N__59334),
            .in3(N__62687),
            .lcout(\c0.n12_adj_4500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_1892_LC_21_19_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1892_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1892_LC_21_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1892_LC_21_19_3  (
            .in0(N__65787),
            .in1(N__61746),
            .in2(N__59058),
            .in3(N__61797),
            .lcout(\c0.n6_adj_4587 ),
            .ltout(\c0.n6_adj_4587_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1889_LC_21_19_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1889_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1889_LC_21_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1889_LC_21_19_4  (
            .in0(N__77673),
            .in1(N__59370),
            .in2(N__59355),
            .in3(N__77811),
            .lcout(\c0.n13461 ),
            .ltout(\c0.n13461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1697_LC_21_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1697_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1697_LC_21_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1697_LC_21_19_5  (
            .in0(N__66496),
            .in1(N__59329),
            .in2(N__59310),
            .in3(N__72242),
            .lcout(\c0.n6227 ),
            .ltout(\c0.n6227_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1398_LC_21_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1398_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1398_LC_21_19_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i2_3_lut_adj_1398_LC_21_19_6  (
            .in0(_gnd_net_),
            .in1(N__62686),
            .in2(N__59307),
            .in3(N__59304),
            .lcout(\c0.n21301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1265_LC_21_19_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1265_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1265_LC_21_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1265_LC_21_19_7  (
            .in0(N__62424),
            .in1(N__62411),
            .in2(N__66501),
            .in3(N__60060),
            .lcout(\c0.n19_adj_4291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1879_LC_21_20_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1879_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1879_LC_21_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1879_LC_21_20_0  (
            .in0(N__59261),
            .in1(N__62720),
            .in2(N__62603),
            .in3(N__59088),
            .lcout(\c0.n21414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i120_LC_21_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i120_LC_21_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i120_LC_21_20_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i120_LC_21_20_1  (
            .in0(N__76385),
            .in1(N__59148),
            .in2(_gnd_net_),
            .in3(N__62591),
            .lcout(data_in_frame_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78752),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1548_LC_21_20_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1548_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1548_LC_21_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1548_LC_21_20_3  (
            .in0(N__59130),
            .in1(N__59109),
            .in2(N__62331),
            .in3(N__62010),
            .lcout(\c0.n23300 ),
            .ltout(\c0.n23300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1567_LC_21_20_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1567_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1567_LC_21_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1567_LC_21_20_4  (
            .in0(N__59082),
            .in1(N__59057),
            .in2(N__59034),
            .in3(N__62721),
            .lcout(\c0.n21_adj_4594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1388_LC_21_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1388_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1388_LC_21_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1388_LC_21_20_5  (
            .in0(_gnd_net_),
            .in1(N__59456),
            .in2(_gnd_net_),
            .in3(N__67180),
            .lcout(\c0.n4_adj_4347 ),
            .ltout(\c0.n4_adj_4347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1376_LC_21_20_6 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1376_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1376_LC_21_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1376_LC_21_20_6  (
            .in0(N__59484),
            .in1(N__80136),
            .in2(N__59463),
            .in3(N__77229),
            .lcout(\c0.n40_adj_4359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i186_LC_21_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i186_LC_21_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i186_LC_21_20_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i186_LC_21_20_7  (
            .in0(N__80328),
            .in1(N__80966),
            .in2(N__59460),
            .in3(N__75224),
            .lcout(\c0.data_in_frame_23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78752),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1700_LC_21_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1700_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1700_LC_21_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1700_LC_21_21_0  (
            .in0(N__73034),
            .in1(N__65904),
            .in2(_gnd_net_),
            .in3(N__63299),
            .lcout(\c0.n22698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_adj_1576_LC_21_21_1 .C_ON=1'b0;
    defparam \c0.i7_2_lut_adj_1576_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_adj_1576_LC_21_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i7_2_lut_adj_1576_LC_21_21_1  (
            .in0(N__66661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66597),
            .lcout(\c0.n30_adj_4357 ),
            .ltout(\c0.n30_adj_4357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1375_LC_21_21_2 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1375_LC_21_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1375_LC_21_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1375_LC_21_21_2  (
            .in0(N__59720),
            .in1(N__66950),
            .in2(N__59445),
            .in3(N__59434),
            .lcout(),
            .ltout(\c0.n42_adj_4358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_21_21_3 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_21_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_LC_21_21_3  (
            .in0(N__59403),
            .in1(N__61926),
            .in2(N__59397),
            .in3(N__59394),
            .lcout(\c0.n34_adj_4361 ),
            .ltout(\c0.n34_adj_4361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1464_LC_21_21_4 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1464_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1464_LC_21_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1464_LC_21_21_4  (
            .in0(N__59385),
            .in1(N__59376),
            .in2(N__59379),
            .in3(N__63170),
            .lcout(\c0.n42_adj_4510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1553_LC_21_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1553_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1553_LC_21_21_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1553_LC_21_21_5  (
            .in0(_gnd_net_),
            .in1(N__75847),
            .in2(_gnd_net_),
            .in3(N__66751),
            .lcout(\c0.n14148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1421_LC_21_21_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1421_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1421_LC_21_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1421_LC_21_21_6  (
            .in0(N__61927),
            .in1(N__66525),
            .in2(N__59731),
            .in3(N__59676),
            .lcout(\c0.n22426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1527_LC_21_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1527_LC_21_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1527_LC_21_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1527_LC_21_21_7  (
            .in0(_gnd_net_),
            .in1(N__67313),
            .in2(_gnd_net_),
            .in3(N__67260),
            .lcout(\c0.n5_adj_4486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_334_2_lut_4_lut_LC_21_22_0 .C_ON=1'b0;
    defparam \c0.i1_rep_334_2_lut_4_lut_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_334_2_lut_4_lut_LC_21_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_rep_334_2_lut_4_lut_LC_21_22_0  (
            .in0(N__67251),
            .in1(N__59589),
            .in2(N__64168),
            .in3(N__67550),
            .lcout(\c0.n25456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1509_LC_21_22_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1509_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1509_LC_21_22_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i11_4_lut_adj_1509_LC_21_22_1  (
            .in0(N__67499),
            .in1(N__59663),
            .in2(N__59640),
            .in3(N__73943),
            .lcout(\c0.n26_adj_4548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1718_LC_21_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1718_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1718_LC_21_22_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1718_LC_21_22_2  (
            .in0(N__64158),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59588),
            .lcout(\c0.n13468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1518_LC_21_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1518_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1518_LC_21_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1518_LC_21_22_3  (
            .in0(_gnd_net_),
            .in1(N__67549),
            .in2(_gnd_net_),
            .in3(N__67250),
            .lcout(\c0.n13490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_3_lut_4_lut_LC_21_22_4 .C_ON=1'b0;
    defparam \c0.i24_3_lut_4_lut_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i24_3_lut_4_lut_LC_21_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_3_lut_4_lut_LC_21_22_4  (
            .in0(N__78026),
            .in1(N__59562),
            .in2(N__59532),
            .in3(N__67500),
            .lcout(),
            .ltout(\c0.n66_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_4_lut_adj_1427_LC_21_22_5 .C_ON=1'b0;
    defparam \c0.i33_4_lut_adj_1427_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i33_4_lut_adj_1427_LC_21_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i33_4_lut_adj_1427_LC_21_22_5  (
            .in0(N__67314),
            .in1(N__59499),
            .in2(N__59508),
            .in3(N__63599),
            .lcout(\c0.n75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_LC_21_22_6 .C_ON=1'b0;
    defparam \c0.i4_3_lut_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_LC_21_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_3_lut_LC_21_22_6  (
            .in0(N__77376),
            .in1(N__74893),
            .in2(_gnd_net_),
            .in3(N__67593),
            .lcout(\c0.n46_adj_4461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_1927_LC_21_22_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_1927_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_1927_LC_21_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_1927_LC_21_22_7  (
            .in0(N__63230),
            .in1(N__68312),
            .in2(_gnd_net_),
            .in3(N__63636),
            .lcout(\c0.n25_adj_4469 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1499_LC_21_23_0 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1499_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1499_LC_21_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1499_LC_21_23_0  (
            .in0(N__67089),
            .in1(N__59919),
            .in2(N__59787),
            .in3(N__59897),
            .lcout(\c0.n53_adj_4538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1510_LC_21_23_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1510_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1510_LC_21_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1510_LC_21_23_1  (
            .in0(N__74778),
            .in1(N__67592),
            .in2(N__59880),
            .in3(N__63598),
            .lcout(),
            .ltout(\c0.n24_adj_4550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1511_LC_21_23_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1511_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1511_LC_21_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1511_LC_21_23_2  (
            .in0(N__59838),
            .in1(N__59826),
            .in2(N__59820),
            .in3(N__73773),
            .lcout(\c0.n21010 ),
            .ltout(\c0.n21010_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_LC_21_23_3 .C_ON=1'b0;
    defparam \c0.i27_4_lut_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_LC_21_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_LC_21_23_3  (
            .in0(N__64089),
            .in1(N__63686),
            .in2(N__59817),
            .in3(N__59814),
            .lcout(\c0.n61_adj_4543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_adj_1501_LC_21_23_4 .C_ON=1'b0;
    defparam \c0.i28_4_lut_adj_1501_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_adj_1501_LC_21_23_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i28_4_lut_adj_1501_LC_21_23_4  (
            .in0(N__59802),
            .in1(N__63567),
            .in2(N__63739),
            .in3(N__63849),
            .lcout(\c0.n62_adj_4541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_adj_1450_LC_21_23_5 .C_ON=1'b0;
    defparam \c0.i4_3_lut_adj_1450_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_adj_1450_LC_21_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i4_3_lut_adj_1450_LC_21_23_5  (
            .in0(_gnd_net_),
            .in1(N__64138),
            .in2(N__67873),
            .in3(N__59786),
            .lcout(\c0.n18_adj_4493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1454_LC_21_24_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1454_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1454_LC_21_24_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i12_4_lut_adj_1454_LC_21_24_1  (
            .in0(N__59763),
            .in1(N__63791),
            .in2(N__75702),
            .in3(N__63642),
            .lcout(),
            .ltout(\c0.n26_adj_4499_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1458_LC_21_24_2 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1458_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1458_LC_21_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1458_LC_21_24_2  (
            .in0(N__62553),
            .in1(N__59754),
            .in2(N__59745),
            .in3(N__63848),
            .lcout(),
            .ltout(\c0.n24441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1506_LC_21_24_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1506_LC_21_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1506_LC_21_24_3 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i12_4_lut_adj_1506_LC_21_24_3  (
            .in0(N__63453),
            .in1(N__63855),
            .in2(N__60003),
            .in3(N__67398),
            .lcout(\c0.n30_adj_4545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_adj_1467_LC_21_24_4 .C_ON=1'b0;
    defparam \c0.i30_4_lut_adj_1467_LC_21_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_adj_1467_LC_21_24_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i30_4_lut_adj_1467_LC_21_24_4  (
            .in0(N__63680),
            .in1(N__63847),
            .in2(N__63741),
            .in3(N__63653),
            .lcout(\c0.n72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i177_LC_21_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i177_LC_21_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i177_LC_21_24_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i177_LC_21_24_5  (
            .in0(N__63499),
            .in1(N__80672),
            .in2(_gnd_net_),
            .in3(N__78915),
            .lcout(data_in_frame_22_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1469_LC_21_24_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1469_LC_21_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1469_LC_21_24_7 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \c0.i2_4_lut_adj_1469_LC_21_24_7  (
            .in0(N__59979),
            .in1(N__67005),
            .in2(N__59967),
            .in3(N__63810),
            .lcout(\c0.n20_adj_4518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i227_LC_21_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i227_LC_21_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i227_LC_21_25_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i227_LC_21_25_0  (
            .in0(N__80079),
            .in1(N__79167),
            .in2(N__63828),
            .in3(N__79482),
            .lcout(\c0.data_in_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78797),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20984_4_lut_LC_22_7_4 .C_ON=1'b0;
    defparam \c0.i20984_4_lut_LC_22_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20984_4_lut_LC_22_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20984_4_lut_LC_22_7_4  (
            .in0(N__67941),
            .in1(N__60644),
            .in2(N__60798),
            .in3(N__60304),
            .lcout(\c0.n24751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1839_LC_22_8_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1839_LC_22_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1839_LC_22_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1839_LC_22_8_0  (
            .in0(_gnd_net_),
            .in1(N__64033),
            .in2(_gnd_net_),
            .in3(N__61767),
            .lcout(\c0.n6_adj_4632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1766_LC_22_8_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1766_LC_22_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1766_LC_22_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i6_4_lut_adj_1766_LC_22_8_2  (
            .in0(N__60303),
            .in1(N__60208),
            .in2(N__68543),
            .in3(N__60637),
            .lcout(),
            .ltout(\c0.n14_adj_4676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1768_LC_22_8_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1768_LC_22_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1768_LC_22_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i7_4_lut_adj_1768_LC_22_8_3  (
            .in0(N__69582),
            .in1(N__64068),
            .in2(N__59934),
            .in3(N__68094),
            .lcout(\c0.data_out_frame_0__7__N_2777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1762_LC_22_8_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1762_LC_22_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1762_LC_22_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1762_LC_22_8_4  (
            .in0(N__68849),
            .in1(N__60636),
            .in2(N__68542),
            .in3(N__69581),
            .lcout(\c0.n24016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20982_4_lut_LC_22_8_5 .C_ON=1'b0;
    defparam \c0.i20982_4_lut_LC_22_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20982_4_lut_LC_22_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20982_4_lut_LC_22_8_5  (
            .in0(N__69583),
            .in1(N__64778),
            .in2(N__60228),
            .in3(N__68795),
            .lcout(\c0.n24749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1935_LC_22_8_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1935_LC_22_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1935_LC_22_8_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.i13_4_lut_adj_1935_LC_22_8_6  (
            .in0(N__68848),
            .in1(N__60566),
            .in2(N__72586),
            .in3(N__60431),
            .lcout(\c0.n37_adj_4738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1881_LC_22_8_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1881_LC_22_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1881_LC_22_8_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1881_LC_22_8_7  (
            .in0(N__72570),
            .in1(N__60302),
            .in2(N__60227),
            .in3(N__68093),
            .lcout(\c0.n24_adj_4717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_2049_LC_22_9_0 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_2049_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_2049_LC_22_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i4_2_lut_adj_2049_LC_22_9_0  (
            .in0(N__60155),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61262),
            .lcout(),
            .ltout(\c0.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_LC_22_9_1 .C_ON=1'b0;
    defparam \c0.i24_4_lut_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_LC_22_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_LC_22_9_1  (
            .in0(N__60012),
            .in1(N__60135),
            .in2(N__60120),
            .in3(N__60117),
            .lcout(),
            .ltout(\c0.n54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_4_lut_adj_1230_LC_22_9_2 .C_ON=1'b0;
    defparam \c0.i29_4_lut_adj_1230_LC_22_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i29_4_lut_adj_1230_LC_22_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i29_4_lut_adj_1230_LC_22_9_2  (
            .in0(N__60099),
            .in1(N__60654),
            .in2(N__60087),
            .in3(N__60084),
            .lcout(\c0.n13821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_22_9_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_22_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_22_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_LC_22_9_3  (
            .in0(N__69894),
            .in1(N__64008),
            .in2(N__64229),
            .in3(N__68141),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_adj_1865_LC_22_9_4 .C_ON=1'b0;
    defparam \c0.i7_2_lut_adj_1865_LC_22_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_adj_1865_LC_22_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i7_2_lut_adj_1865_LC_22_9_4  (
            .in0(_gnd_net_),
            .in1(N__68840),
            .in2(_gnd_net_),
            .in3(N__68081),
            .lcout(\c0.n37 ),
            .ltout(\c0.n37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1869_LC_22_9_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1869_LC_22_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1869_LC_22_9_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1869_LC_22_9_5  (
            .in0(N__64012),
            .in1(N__68028),
            .in2(N__60753),
            .in3(N__68140),
            .lcout(\c0.n22647 ),
            .ltout(\c0.n22647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1877_LC_22_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1877_LC_22_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1877_LC_22_9_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1877_LC_22_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60750),
            .in3(N__68958),
            .lcout(\c0.n16_adj_4716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20980_4_lut_LC_22_9_7 .C_ON=1'b0;
    defparam \c0.i20980_4_lut_LC_22_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i20980_4_lut_LC_22_9_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20980_4_lut_LC_22_9_7  (
            .in0(N__68082),
            .in1(N__68752),
            .in2(N__60747),
            .in3(N__68029),
            .lcout(\c0.n24747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_1614_LC_22_10_0 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_1614_LC_22_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_1614_LC_22_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_1614_LC_22_10_0  (
            .in0(N__68733),
            .in1(N__68512),
            .in2(N__65696),
            .in3(N__68846),
            .lcout(),
            .ltout(\c0.n14_adj_4616_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1899_LC_22_10_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1899_LC_22_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1899_LC_22_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1899_LC_22_10_1  (
            .in0(N__68781),
            .in1(N__60699),
            .in2(N__60693),
            .in3(N__64006),
            .lcout(\c0.data_out_frame_0__7__N_2743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i38_LC_22_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i38_LC_22_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i38_LC_22_10_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i38_LC_22_10_2  (
            .in0(N__79588),
            .in1(N__79988),
            .in2(N__65697),
            .in3(N__70146),
            .lcout(\c0.data_in_frame_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78799),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_LC_22_10_3 .C_ON=1'b0;
    defparam \c0.i25_4_lut_LC_22_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_LC_22_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_LC_22_10_3  (
            .in0(N__64293),
            .in1(N__60690),
            .in2(N__60666),
            .in3(N__68034),
            .lcout(\c0.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i33_LC_22_10_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i33_LC_22_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i33_LC_22_10_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i33_LC_22_10_4  (
            .in0(N__80742),
            .in1(N__79987),
            .in2(N__60899),
            .in3(N__70145),
            .lcout(\c0.data_in_frame_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78799),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1864_LC_22_10_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1864_LC_22_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1864_LC_22_10_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1864_LC_22_10_5  (
            .in0(N__68780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68671),
            .lcout(\c0.n5_adj_4711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_LC_22_10_6 .C_ON=1'b0;
    defparam \c0.i9_3_lut_LC_22_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_LC_22_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i9_3_lut_LC_22_10_6  (
            .in0(N__60891),
            .in1(N__61101),
            .in2(_gnd_net_),
            .in3(N__60854),
            .lcout(\c0.n24_adj_4724 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i39_LC_22_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i39_LC_22_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i39_LC_22_10_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i39_LC_22_10_7  (
            .in0(N__70144),
            .in1(N__73289),
            .in2(N__80032),
            .in3(N__64007),
            .lcout(\c0.data_in_frame_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78799),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1882_LC_22_11_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1882_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1882_LC_22_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1882_LC_22_11_0  (
            .in0(N__61057),
            .in1(N__60987),
            .in2(N__60796),
            .in3(N__60912),
            .lcout(),
            .ltout(\c0.n28_adj_4718_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1891_LC_22_11_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1891_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1891_LC_22_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1891_LC_22_11_1  (
            .in0(N__60981),
            .in1(N__68531),
            .in2(N__60969),
            .in3(N__60966),
            .lcout(\c0.n23_adj_4599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1872_LC_22_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1872_LC_22_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1872_LC_22_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1872_LC_22_11_2  (
            .in0(_gnd_net_),
            .in1(N__64259),
            .in2(_gnd_net_),
            .in3(N__69546),
            .lcout(\c0.n4_adj_4446 ),
            .ltout(\c0.n4_adj_4446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1876_LC_22_11_3 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1876_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1876_LC_22_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_3_lut_adj_1876_LC_22_11_3  (
            .in0(_gnd_net_),
            .in1(N__68727),
            .in2(N__60915),
            .in3(N__61288),
            .lcout(\c0.n26_adj_4714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_22_11_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_22_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_22_11_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i17_LC_22_11_4  (
            .in0(N__80741),
            .in1(N__70018),
            .in2(N__60797),
            .in3(N__69091),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78791),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1757_LC_22_11_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1757_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1757_LC_22_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1757_LC_22_11_5  (
            .in0(N__60774),
            .in1(N__60882),
            .in2(_gnd_net_),
            .in3(N__60855),
            .lcout(\c0.n23597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1705_LC_22_11_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1705_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1705_LC_22_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1705_LC_22_11_6  (
            .in0(N__68959),
            .in1(N__60773),
            .in2(N__61298),
            .in3(N__64260),
            .lcout(\c0.n10_adj_4664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_LC_22_11_7 .C_ON=1'b0;
    defparam \c0.i12_3_lut_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_LC_22_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i12_3_lut_LC_22_11_7  (
            .in0(N__61255),
            .in1(N__70694),
            .in2(_gnd_net_),
            .in3(N__67985),
            .lcout(\c0.n48_adj_4227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i69_4_lut_LC_22_12_0 .C_ON=1'b0;
    defparam \c0.i69_4_lut_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i69_4_lut_LC_22_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i69_4_lut_LC_22_12_0  (
            .in0(N__61113),
            .in1(N__70715),
            .in2(N__65369),
            .in3(N__69700),
            .lcout(\c0.n150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_1179_LC_22_12_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_1179_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_1179_LC_22_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_1179_LC_22_12_1  (
            .in0(_gnd_net_),
            .in1(N__65201),
            .in2(_gnd_net_),
            .in3(N__65220),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_1665_LC_22_12_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_1665_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_1665_LC_22_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_1665_LC_22_12_2  (
            .in0(N__65221),
            .in1(N__65202),
            .in2(_gnd_net_),
            .in3(N__65108),
            .lcout(\c0.n13651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1200_LC_22_12_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1200_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1200_LC_22_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1200_LC_22_12_3  (
            .in0(N__64562),
            .in1(N__61111),
            .in2(N__64686),
            .in3(N__71119),
            .lcout(),
            .ltout(\c0.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_LC_22_12_4 .C_ON=1'b0;
    defparam \c0.i14_3_lut_LC_22_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_LC_22_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i14_3_lut_LC_22_12_4  (
            .in0(_gnd_net_),
            .in1(N__61175),
            .in2(N__61152),
            .in3(N__61149),
            .lcout(\c0.n23528 ),
            .ltout(\c0.n23528_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_22_12_5 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_22_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_22_12_5  (
            .in0(N__65988),
            .in1(N__64967),
            .in2(N__61128),
            .in3(N__61341),
            .lcout(),
            .ltout(\c0.n34_adj_4278_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1259_LC_22_12_6 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1259_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1259_LC_22_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1259_LC_22_12_6  (
            .in0(N__66227),
            .in1(N__68604),
            .in2(N__61125),
            .in3(N__68532),
            .lcout(\c0.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_2_lut_LC_22_12_7 .C_ON=1'b0;
    defparam \c0.i24_2_lut_LC_22_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i24_2_lut_LC_22_12_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i24_2_lut_LC_22_12_7  (
            .in0(N__64563),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61112),
            .lcout(\c0.n60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1848_LC_22_13_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1848_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1848_LC_22_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1848_LC_22_13_0  (
            .in0(N__62119),
            .in1(N__71209),
            .in2(N__64966),
            .in3(N__71118),
            .lcout(),
            .ltout(\c0.n30_adj_4705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1850_LC_22_13_1 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1850_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1850_LC_22_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1850_LC_22_13_1  (
            .in0(N__69758),
            .in1(N__69693),
            .in2(N__61347),
            .in3(N__62033),
            .lcout(\c0.n23523 ),
            .ltout(\c0.n23523_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_LC_22_13_2 .C_ON=1'b0;
    defparam \c0.i11_3_lut_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_LC_22_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_3_lut_LC_22_13_2  (
            .in0(_gnd_net_),
            .in1(N__65591),
            .in2(N__61344),
            .in3(N__65549),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1728_LC_22_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1728_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1728_LC_22_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1728_LC_22_13_3  (
            .in0(N__66246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65525),
            .lcout(\c0.n4_adj_4261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i99_LC_22_13_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i99_LC_22_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i99_LC_22_13_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i99_LC_22_13_4  (
            .in0(N__80060),
            .in1(N__73665),
            .in2(N__65039),
            .in3(N__79209),
            .lcout(\c0.data_in_frame_12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_2013_LC_22_13_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_2013_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_2013_LC_22_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_2013_LC_22_13_5  (
            .in0(N__64191),
            .in1(N__70672),
            .in2(_gnd_net_),
            .in3(N__65638),
            .lcout(\c0.n6_adj_4209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i72_LC_22_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i72_LC_22_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i72_LC_22_13_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i72_LC_22_13_6  (
            .in0(N__76378),
            .in1(N__65639),
            .in2(N__72978),
            .in3(N__73666),
            .lcout(\c0.data_in_frame_8_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1838_LC_22_14_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1838_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1838_LC_22_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1838_LC_22_14_0  (
            .in0(N__65631),
            .in1(N__61333),
            .in2(N__61479),
            .in3(N__61488),
            .lcout(\c0.n7_adj_4634 ),
            .ltout(\c0.n7_adj_4634_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1775_LC_22_14_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1775_LC_22_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1775_LC_22_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1775_LC_22_14_1  (
            .in0(N__71177),
            .in1(N__70958),
            .in2(N__61305),
            .in3(N__65297),
            .lcout(\c0.n5807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1776_LC_22_14_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1776_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1776_LC_22_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1776_LC_22_14_2  (
            .in0(N__65296),
            .in1(N__64506),
            .in2(N__71176),
            .in3(N__61738),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i40_4_lut_LC_22_14_3 .C_ON=1'b0;
    defparam \c0.i40_4_lut_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i40_4_lut_LC_22_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i40_4_lut_LC_22_14_3  (
            .in0(N__61589),
            .in1(N__61782),
            .in2(N__61745),
            .in3(N__65630),
            .lcout(),
            .ltout(\c0.n96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i48_4_lut_adj_1406_LC_22_14_4 .C_ON=1'b0;
    defparam \c0.i48_4_lut_adj_1406_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i48_4_lut_adj_1406_LC_22_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i48_4_lut_adj_1406_LC_22_14_4  (
            .in0(N__61475),
            .in1(N__61487),
            .in2(N__61560),
            .in3(N__61557),
            .lcout(\c0.n104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1242_LC_22_14_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1242_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1242_LC_22_14_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1242_LC_22_14_5  (
            .in0(_gnd_net_),
            .in1(N__69301),
            .in2(_gnd_net_),
            .in3(N__70618),
            .lcout(\c0.n7_adj_4253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_22_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_22_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_22_14_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0__i52_LC_22_14_6  (
            .in0(N__68432),
            .in1(_gnd_net_),
            .in2(N__77121),
            .in3(N__77856),
            .lcout(data_in_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1241_LC_22_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1241_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1241_LC_22_14_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1241_LC_22_14_7  (
            .in0(N__76036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65327),
            .lcout(\c0.n5_adj_4252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1676_LC_22_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1676_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1676_LC_22_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1676_LC_22_15_0  (
            .in0(N__61852),
            .in1(N__61467),
            .in2(N__65337),
            .in3(N__65226),
            .lcout(\c0.n13734 ),
            .ltout(\c0.n13734_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_1675_LC_22_15_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_1675_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_1675_LC_22_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_1675_LC_22_15_1  (
            .in0(N__61741),
            .in1(_gnd_net_),
            .in2(N__61440),
            .in3(N__65772),
            .lcout(\c0.n18_adj_4580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1719_LC_22_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1719_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1719_LC_22_15_2 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1719_LC_22_15_2  (
            .in0(N__61437),
            .in1(N__61392),
            .in2(_gnd_net_),
            .in3(N__62271),
            .lcout(\c0.n22120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1656_LC_22_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1656_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1656_LC_22_15_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1656_LC_22_15_3  (
            .in0(_gnd_net_),
            .in1(N__65331),
            .in2(_gnd_net_),
            .in3(N__61851),
            .lcout(\c0.n22176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1583_LC_22_15_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1583_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1583_LC_22_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1583_LC_22_15_5  (
            .in0(N__64373),
            .in1(N__65150),
            .in2(N__61833),
            .in3(N__65111),
            .lcout(\c0.n13738 ),
            .ltout(\c0.n13738_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1893_LC_22_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1893_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1893_LC_22_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1893_LC_22_15_6  (
            .in0(N__61811),
            .in1(N__61739),
            .in2(N__61800),
            .in3(N__61792),
            .lcout(\c0.n22782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1667_LC_22_15_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1667_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1667_LC_22_15_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1667_LC_22_15_7  (
            .in0(N__61740),
            .in1(N__61691),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n5_adj_4310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_1855_LC_22_16_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_1855_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_1855_LC_22_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_1855_LC_22_16_0  (
            .in0(_gnd_net_),
            .in1(N__62141),
            .in2(_gnd_net_),
            .in3(N__62132),
            .lcout(),
            .ltout(\c0.n39_adj_4708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_adj_1857_LC_22_16_1 .C_ON=1'b0;
    defparam \c0.i28_4_lut_adj_1857_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_adj_1857_LC_22_16_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i28_4_lut_adj_1857_LC_22_16_1  (
            .in0(N__66161),
            .in1(N__62799),
            .in2(N__61680),
            .in3(N__61629),
            .lcout(),
            .ltout(\c0.n64_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i34_4_lut_LC_22_16_2 .C_ON=1'b0;
    defparam \c0.i34_4_lut_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i34_4_lut_LC_22_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i34_4_lut_LC_22_16_2  (
            .in0(N__61677),
            .in1(N__69765),
            .in2(N__61662),
            .in3(N__69701),
            .lcout(\c0.n70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1856_LC_22_16_3 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1856_LC_22_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1856_LC_22_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1856_LC_22_16_3  (
            .in0(N__72468),
            .in1(N__66010),
            .in2(N__61659),
            .in3(N__65435),
            .lcout(\c0.n55_adj_4709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1227_LC_22_16_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1227_LC_22_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1227_LC_22_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1227_LC_22_16_4  (
            .in0(N__68982),
            .in1(N__65009),
            .in2(N__61623),
            .in3(N__64655),
            .lcout(\c0.n10_adj_4247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i43_4_lut_LC_22_16_5 .C_ON=1'b0;
    defparam \c0.i43_4_lut_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i43_4_lut_LC_22_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i43_4_lut_LC_22_16_5  (
            .in0(N__73392),
            .in1(N__62742),
            .in2(N__62806),
            .in3(N__66464),
            .lcout(\c0.n124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1417_LC_22_16_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1417_LC_22_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1417_LC_22_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1417_LC_22_16_6  (
            .in0(N__65436),
            .in1(N__62142),
            .in2(N__62807),
            .in3(N__62133),
            .lcout(\c0.n12_adj_4455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_22_17_0 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_22_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_LC_22_17_0  (
            .in0(N__62124),
            .in1(N__62886),
            .in2(N__64989),
            .in3(N__62091),
            .lcout(),
            .ltout(\c0.n59_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i35_4_lut_LC_22_17_1 .C_ON=1'b0;
    defparam \c0.i35_4_lut_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i35_4_lut_LC_22_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i35_4_lut_LC_22_17_1  (
            .in0(N__62052),
            .in1(N__62037),
            .in2(N__62022),
            .in3(N__62019),
            .lcout(\c0.n24444 ),
            .ltout(\c0.n24444_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_22_17_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_22_17_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_LC_22_17_2  (
            .in0(N__62919),
            .in1(N__62887),
            .in2(N__62013),
            .in3(N__62756),
            .lcout(\c0.n13604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1523_LC_22_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1523_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1523_LC_22_17_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_1523_LC_22_17_3  (
            .in0(N__62757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62356),
            .lcout(\c0.n21282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1264_LC_22_17_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1264_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1264_LC_22_17_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i2_3_lut_adj_1264_LC_22_17_4  (
            .in0(_gnd_net_),
            .in1(N__61995),
            .in2(N__62361),
            .in3(N__62758),
            .lcout(\c0.n23224 ),
            .ltout(\c0.n23224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_2028_LC_22_17_5 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_2028_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_2028_LC_22_17_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_2028_LC_22_17_5  (
            .in0(N__61949),
            .in1(N__66608),
            .in2(N__61938),
            .in3(N__66364),
            .lcout(\c0.n21409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1577_LC_22_17_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1577_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1577_LC_22_17_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1577_LC_22_17_6  (
            .in0(N__61902),
            .in1(N__62710),
            .in2(N__66117),
            .in3(N__62688),
            .lcout(\c0.n10_adj_4602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_2027_LC_22_17_7 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_2027_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_2027_LC_22_17_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_2027_LC_22_17_7  (
            .in0(N__72021),
            .in1(N__66335),
            .in2(N__69645),
            .in3(N__66365),
            .lcout(\c0.n21404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1630_LC_22_18_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1630_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1630_LC_22_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1630_LC_22_18_0  (
            .in0(N__62355),
            .in1(N__62613),
            .in2(N__62643),
            .in3(N__66133),
            .lcout(\c0.n10_adj_4630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_2034_LC_22_18_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_2034_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_2034_LC_22_18_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_2034_LC_22_18_1  (
            .in0(N__62639),
            .in1(N__62994),
            .in2(N__62616),
            .in3(N__62354),
            .lcout(\c0.n12_adj_4246 ),
            .ltout(\c0.n12_adj_4246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1419_LC_22_18_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1419_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1419_LC_22_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1419_LC_22_18_2  (
            .in0(N__71646),
            .in1(N__62766),
            .in2(N__62559),
            .in3(N__66134),
            .lcout(\c0.n23691 ),
            .ltout(\c0.n23691_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1371_LC_22_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1371_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1371_LC_22_18_3 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_1371_LC_22_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62556),
            .in3(N__66871),
            .lcout(\c0.n20543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1581_LC_22_18_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1581_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1581_LC_22_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1581_LC_22_18_4  (
            .in0(N__62532),
            .in1(N__62493),
            .in2(_gnd_net_),
            .in3(N__62487),
            .lcout(\c0.n14189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_1706_LC_22_18_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1706_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1706_LC_22_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1706_LC_22_18_5  (
            .in0(N__62463),
            .in1(N__62423),
            .in2(N__62412),
            .in3(N__62353),
            .lcout(\c0.n7_adj_4581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_3_i3_2_lut_LC_22_18_7 .C_ON=1'b0;
    defparam \c0.select_367_Select_3_i3_2_lut_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_3_i3_2_lut_LC_22_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_3_i3_2_lut_LC_22_18_7  (
            .in0(_gnd_net_),
            .in1(N__62295),
            .in2(_gnd_net_),
            .in3(N__71537),
            .lcout(\c0.n3_adj_4430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_1852_LC_22_19_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_1852_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_1852_LC_22_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_1852_LC_22_19_0  (
            .in0(_gnd_net_),
            .in1(N__62920),
            .in2(_gnd_net_),
            .in3(N__62894),
            .lcout(\c0.n20467 ),
            .ltout(\c0.n20467_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_1754_LC_22_19_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_1754_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_1754_LC_22_19_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_1754_LC_22_19_1  (
            .in0(N__62768),
            .in1(N__62939),
            .in2(N__62985),
            .in3(N__75939),
            .lcout(\c0.n17_adj_4354 ),
            .ltout(\c0.n17_adj_4354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_1373_LC_22_19_2 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_1373_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_1373_LC_22_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_adj_1373_LC_22_19_2  (
            .in0(N__63522),
            .in1(N__62981),
            .in2(N__62943),
            .in3(N__67351),
            .lcout(\c0.n58_adj_4355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1689_LC_22_19_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1689_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1689_LC_22_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1689_LC_22_19_3  (
            .in0(N__62769),
            .in1(N__62940),
            .in2(N__62927),
            .in3(N__62895),
            .lcout(\c0.n21295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3286_2_lut_LC_22_19_4 .C_ON=1'b0;
    defparam \c0.i3286_2_lut_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3286_2_lut_LC_22_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3286_2_lut_LC_22_19_4  (
            .in0(N__72089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62848),
            .lcout(\c0.n5965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i103_LC_22_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i103_LC_22_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i103_LC_22_19_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i103_LC_22_19_5  (
            .in0(N__80016),
            .in1(N__73708),
            .in2(N__73347),
            .in3(N__62795),
            .lcout(\c0.data_in_frame_12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78753),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i183_LC_22_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i183_LC_22_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i183_LC_22_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i183_LC_22_19_6  (
            .in0(N__63523),
            .in1(N__73331),
            .in2(_gnd_net_),
            .in3(N__78904),
            .lcout(data_in_frame_22_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78753),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1225_LC_22_19_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1225_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1225_LC_22_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1225_LC_22_19_7  (
            .in0(N__62767),
            .in1(N__66135),
            .in2(N__77209),
            .in3(N__62727),
            .lcout(\c0.n21299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1547_LC_22_20_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1547_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1547_LC_22_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1547_LC_22_20_0  (
            .in0(N__63108),
            .in1(N__63120),
            .in2(N__72594),
            .in3(N__66033),
            .lcout(\c0.n23453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_2_lut_4_lut_LC_22_20_1 .C_ON=1'b0;
    defparam \c0.i10_2_lut_4_lut_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_2_lut_4_lut_LC_22_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_2_lut_4_lut_LC_22_20_1  (
            .in0(N__72319),
            .in1(N__77879),
            .in2(N__63156),
            .in3(N__77810),
            .lcout(\c0.n25_adj_4579 ),
            .ltout(\c0.n25_adj_4579_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1707_LC_22_20_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1707_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1707_LC_22_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1707_LC_22_20_2  (
            .in0(N__63096),
            .in1(N__66032),
            .in2(N__63114),
            .in3(N__65385),
            .lcout(\c0.n23433 ),
            .ltout(\c0.n23433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_4_lut_LC_22_20_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_4_lut_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_4_lut_LC_22_20_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i17_4_lut_4_lut_LC_22_20_3  (
            .in0(N__72320),
            .in1(_gnd_net_),
            .in2(N__63111),
            .in3(N__77578),
            .lcout(\c0.n43_adj_4661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_LC_22_20_4 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_LC_22_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i9_2_lut_3_lut_LC_22_20_4  (
            .in0(N__63107),
            .in1(_gnd_net_),
            .in2(N__74963),
            .in3(N__65427),
            .lcout(\c0.n24_adj_4655 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_1910_LC_22_20_5 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_1910_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_1910_LC_22_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_adj_1910_LC_22_20_5  (
            .in0(N__63090),
            .in1(N__63069),
            .in2(N__63063),
            .in3(N__65814),
            .lcout(),
            .ltout(\c0.n50_adj_4340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_1361_LC_22_20_6 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_1361_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_1361_LC_22_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_adj_1361_LC_22_20_6  (
            .in0(N__63051),
            .in1(N__63039),
            .in2(N__63021),
            .in3(N__66375),
            .lcout(\c0.n28_adj_4343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1571_LC_22_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1571_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1571_LC_22_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1571_LC_22_21_0  (
            .in0(_gnd_net_),
            .in1(N__65903),
            .in2(_gnd_net_),
            .in3(N__63295),
            .lcout(\c0.n22375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1448_LC_22_21_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1448_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1448_LC_22_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_1448_LC_22_21_1  (
            .in0(N__63011),
            .in1(N__67082),
            .in2(N__75700),
            .in3(N__63790),
            .lcout(\c0.n39_adj_4487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1965_LC_22_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1965_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1965_LC_22_21_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1965_LC_22_21_2  (
            .in0(N__63345),
            .in1(N__63379),
            .in2(_gnd_net_),
            .in3(N__66919),
            .lcout(\c0.n12559 ),
            .ltout(\c0.n12559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_1731_LC_22_21_3 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1731_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1731_LC_22_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1731_LC_22_21_3  (
            .in0(N__73033),
            .in1(N__66750),
            .in2(N__63474),
            .in3(N__63464),
            .lcout(\c0.n21316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1457_LC_22_21_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1457_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1457_LC_22_21_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i5_3_lut_adj_1457_LC_22_21_4  (
            .in0(N__68365),
            .in1(N__77307),
            .in2(_gnd_net_),
            .in3(N__66827),
            .lcout(\c0.n24451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1966_LC_22_21_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1966_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1966_LC_22_21_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1966_LC_22_21_5  (
            .in0(N__66985),
            .in1(N__63346),
            .in2(_gnd_net_),
            .in3(N__63380),
            .lcout(\c0.n6_adj_4459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_22_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_22_21_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_22_21_6  (
            .in0(N__63440),
            .in1(N__63378),
            .in2(N__63348),
            .in3(N__65862),
            .lcout(\c0.n21275 ),
            .ltout(\c0.n21275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1400_LC_22_21_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1400_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1400_LC_22_21_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_1400_LC_22_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__63279),
            .in3(N__80135),
            .lcout(\c0.n14_adj_4440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_2_lut_4_lut_LC_22_22_0 .C_ON=1'b0;
    defparam \c0.i29_2_lut_4_lut_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i29_2_lut_4_lut_LC_22_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i29_2_lut_4_lut_LC_22_22_0  (
            .in0(N__63635),
            .in1(N__67056),
            .in2(N__63174),
            .in3(N__77955),
            .lcout(\c0.n63_adj_4516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_LC_22_22_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_LC_22_22_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i6_2_lut_LC_22_22_1  (
            .in0(N__78018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67491),
            .lcout(\c0.n48_adj_4365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_3_lut_adj_1921_LC_22_22_2 .C_ON=1'b0;
    defparam \c0.i12_2_lut_3_lut_adj_1921_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_3_lut_adj_1921_LC_22_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i12_2_lut_3_lut_adj_1921_LC_22_22_2  (
            .in0(N__63211),
            .in1(N__67163),
            .in2(_gnd_net_),
            .in3(N__68311),
            .lcout(\c0.n46 ),
            .ltout(\c0.n46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_LC_22_22_3 .C_ON=1'b0;
    defparam \c0.i23_3_lut_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_LC_22_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i23_3_lut_LC_22_22_3  (
            .in0(_gnd_net_),
            .in1(N__77938),
            .in2(N__63159),
            .in3(N__63634),
            .lcout(),
            .ltout(\c0.n57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1381_LC_22_22_4 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1381_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1381_LC_22_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1381_LC_22_22_4  (
            .in0(N__72366),
            .in1(N__66998),
            .in2(N__63621),
            .in3(N__63618),
            .lcout(\c0.n21426 ),
            .ltout(\c0.n21426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1753_LC_22_22_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1753_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1753_LC_22_22_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1753_LC_22_22_5  (
            .in0(_gnd_net_),
            .in1(N__74815),
            .in2(N__63612),
            .in3(N__63782),
            .lcout(\c0.n23032 ),
            .ltout(\c0.n23032_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1532_LC_22_22_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1532_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1532_LC_22_22_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1532_LC_22_22_6  (
            .in0(N__73809),
            .in1(N__73797),
            .in2(N__63582),
            .in3(N__67591),
            .lcout(\c0.n23209 ),
            .ltout(\c0.n23209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_1441_LC_22_22_7 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_1441_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_1441_LC_22_22_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_adj_1441_LC_22_22_7  (
            .in0(N__78019),
            .in1(N__63579),
            .in2(N__63570),
            .in3(N__67492),
            .lcout(\c0.n56_adj_4479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1928_LC_22_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1928_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1928_LC_22_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1928_LC_22_23_0  (
            .in0(N__77190),
            .in1(N__77730),
            .in2(N__73908),
            .in3(N__63561),
            .lcout(\c0.n20802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_1555_LC_22_23_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_1555_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_1555_LC_22_23_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_1555_LC_22_23_1  (
            .in0(_gnd_net_),
            .in1(N__63543),
            .in2(_gnd_net_),
            .in3(N__67164),
            .lcout(\c0.n26_adj_4470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i175_LC_22_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i175_LC_22_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i175_LC_22_23_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i175_LC_22_23_2  (
            .in0(N__67214),
            .in1(N__73326),
            .in2(_gnd_net_),
            .in3(N__67664),
            .lcout(data_in_frame_21_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1558_LC_22_23_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1558_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1558_LC_22_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1558_LC_22_23_3  (
            .in0(N__63506),
            .in1(N__77151),
            .in2(N__67218),
            .in3(N__66899),
            .lcout(\c0.n22340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1380_LC_22_23_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1380_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1380_LC_22_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1380_LC_22_23_5  (
            .in0(_gnd_net_),
            .in1(N__74811),
            .in2(_gnd_net_),
            .in3(N__63787),
            .lcout(),
            .ltout(\c0.n7_adj_4364_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1422_LC_22_23_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1422_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1422_LC_22_23_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1422_LC_22_23_6  (
            .in0(N__67213),
            .in1(N__63972),
            .in2(N__63945),
            .in3(N__63932),
            .lcout(\c0.n23031 ),
            .ltout(\c0.n23031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1430_LC_22_23_7 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1430_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1430_LC_22_23_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i15_4_lut_adj_1430_LC_22_23_7  (
            .in0(N__77958),
            .in1(N__63727),
            .in2(N__63921),
            .in3(N__63918),
            .lcout(\c0.n39_adj_4467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1461_LC_22_24_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1461_LC_22_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1461_LC_22_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1461_LC_22_24_1  (
            .in0(N__63685),
            .in1(N__74904),
            .in2(N__63888),
            .in3(N__68247),
            .lcout(\c0.n24482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1425_LC_22_24_2 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1425_LC_22_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1425_LC_22_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1425_LC_22_24_2  (
            .in0(N__63803),
            .in1(N__63788),
            .in2(N__63740),
            .in3(N__63846),
            .lcout(),
            .ltout(\c0.n36_adj_4460_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1465_LC_22_24_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1465_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1465_LC_22_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1465_LC_22_24_3  (
            .in0(N__63824),
            .in1(N__77957),
            .in2(N__63813),
            .in3(N__72372),
            .lcout(\c0.n41_adj_4511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1431_LC_22_24_4 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1431_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1431_LC_22_24_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_1431_LC_22_24_4  (
            .in0(N__63804),
            .in1(N__74816),
            .in2(N__63687),
            .in3(N__63789),
            .lcout(\c0.n38_adj_4468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1554_LC_22_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1554_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1554_LC_22_24_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1554_LC_22_24_5  (
            .in0(N__64177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66811),
            .lcout(\c0.n5_adj_4472 ),
            .ltout(\c0.n5_adj_4472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1452_LC_22_24_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1452_LC_22_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1452_LC_22_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1452_LC_22_24_6  (
            .in0(N__63735),
            .in1(N__63684),
            .in2(N__63657),
            .in3(N__63654),
            .lcout(\c0.n24_adj_4496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1738_LC_22_24_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1738_LC_22_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1738_LC_22_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1738_LC_22_24_7  (
            .in0(N__64178),
            .in1(N__66812),
            .in2(N__67863),
            .in3(N__64143),
            .lcout(\c0.n39_adj_4515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_23_7_3 .C_ON=1'b0;
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_23_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_23_7_3 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.equal_87_i9_2_lut_3_lut_LC_23_7_3  (
            .in0(N__74348),
            .in1(N__74642),
            .in2(_gnd_net_),
            .in3(N__74507),
            .lcout(\c0.n9_adj_4552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1764_LC_23_8_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1764_LC_23_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1764_LC_23_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i2_2_lut_adj_1764_LC_23_8_5  (
            .in0(_gnd_net_),
            .in1(N__68751),
            .in2(_gnd_net_),
            .in3(N__68850),
            .lcout(\c0.n10_adj_4675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i89_LC_23_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i89_LC_23_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i89_LC_23_8_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i89_LC_23_8_7  (
            .in0(N__76629),
            .in1(N__73716),
            .in2(N__64048),
            .in3(N__80740),
            .lcout(\c0.data_in_frame_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78818),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_2022_LC_23_9_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_2022_LC_23_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_2022_LC_23_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_2022_LC_23_9_0  (
            .in0(N__68108),
            .in1(N__68030),
            .in2(N__64013),
            .in3(N__68841),
            .lcout(\c0.n23282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1605_LC_23_9_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1605_LC_23_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1605_LC_23_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1605_LC_23_9_1  (
            .in0(N__68842),
            .in1(_gnd_net_),
            .in2(N__68039),
            .in3(N__68110),
            .lcout(\c0.n23283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1969_LC_23_9_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1969_LC_23_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1969_LC_23_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1969_LC_23_9_2  (
            .in0(N__67968),
            .in1(N__64491),
            .in2(N__64544),
            .in3(N__68215),
            .lcout(\c0.n8_adj_4216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i37_LC_23_9_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i37_LC_23_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i37_LC_23_9_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i37_LC_23_9_3  (
            .in0(N__70081),
            .in1(N__68677),
            .in2(N__79954),
            .in3(N__71945),
            .lcout(\c0.data_in_frame_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78815),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_23_9_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_23_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_23_9_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i20_LC_23_9_4  (
            .in0(N__77110),
            .in1(N__70082),
            .in2(N__68796),
            .in3(N__69211),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78815),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_23_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_23_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_23_9_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i21_LC_23_9_5  (
            .in0(N__69210),
            .in1(N__68038),
            .in2(N__70150),
            .in3(N__71944),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78815),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_23_9_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_23_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_23_9_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i3_LC_23_9_6  (
            .in0(N__72925),
            .in1(N__70083),
            .in2(N__79204),
            .in3(N__68843),
            .lcout(\c0.data_in_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78815),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1330_LC_23_9_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1330_LC_23_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1330_LC_23_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1330_LC_23_9_7  (
            .in0(N__67942),
            .in1(N__68527),
            .in2(N__64901),
            .in3(N__68109),
            .lcout(\c0.n21_adj_4327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1602_LC_23_10_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1602_LC_23_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1602_LC_23_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1602_LC_23_10_0  (
            .in0(N__68161),
            .in1(N__64819),
            .in2(N__70277),
            .in3(N__64212),
            .lcout(\c0.n7_adj_4226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1546_LC_23_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1546_LC_23_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1546_LC_23_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1546_LC_23_10_1  (
            .in0(N__64818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68162),
            .lcout(\c0.n4_adj_4211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i40_LC_23_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i40_LC_23_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i40_LC_23_10_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i40_LC_23_10_2  (
            .in0(N__70142),
            .in1(N__80030),
            .in2(N__76294),
            .in3(N__64820),
            .lcout(\c0.data_in_frame_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78807),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i36_LC_23_10_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i36_LC_23_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i36_LC_23_10_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i36_LC_23_10_3  (
            .in0(N__80029),
            .in1(N__70143),
            .in2(N__68969),
            .in3(N__77131),
            .lcout(\c0.data_in_frame_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78807),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1713_LC_23_10_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1713_LC_23_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1713_LC_23_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1713_LC_23_10_4  (
            .in0(N__68160),
            .in1(N__64817),
            .in2(_gnd_net_),
            .in3(N__64211),
            .lcout(\c0.n13904 ),
            .ltout(\c0.n13904_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1328_LC_23_10_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1328_LC_23_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1328_LC_23_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1328_LC_23_10_5  (
            .in0(N__67967),
            .in1(N__69480),
            .in2(N__64203),
            .in3(N__68645),
            .lcout(),
            .ltout(\c0.n19_adj_4324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1343_LC_23_10_6 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1343_LC_23_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1343_LC_23_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_3_lut_adj_1343_LC_23_10_6  (
            .in0(_gnd_net_),
            .in1(N__64200),
            .in2(N__64194),
            .in3(N__68889),
            .lcout(\c0.n22417 ),
            .ltout(\c0.n22417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_LC_23_10_7 .C_ON=1'b0;
    defparam \c0.i30_4_lut_LC_23_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_LC_23_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i30_4_lut_LC_23_10_7  (
            .in0(N__64457),
            .in1(N__64360),
            .in2(N__64416),
            .in3(N__64413),
            .lcout(\c0.n86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_4_lut_LC_23_11_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_4_lut_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_4_lut_LC_23_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_4_lut_LC_23_11_0  (
            .in0(N__69549),
            .in1(N__69481),
            .in2(N__68927),
            .in3(N__72563),
            .lcout(\c0.n13085 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_4_lut_LC_23_11_1 .C_ON=1'b0;
    defparam \c0.i20_3_lut_4_lut_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_4_lut_LC_23_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_3_lut_4_lut_LC_23_11_1  (
            .in0(N__69788),
            .in1(N__70215),
            .in2(N__69832),
            .in3(N__64341),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1997_LC_23_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1997_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1997_LC_23_11_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1997_LC_23_11_2  (
            .in0(N__74525),
            .in1(N__74632),
            .in2(N__74381),
            .in3(N__70014),
            .lcout(n22121),
            .ltout(n22121_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_23_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_23_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_23_11_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0__i55_LC_23_11_3  (
            .in0(N__64283),
            .in1(_gnd_net_),
            .in2(N__64287),
            .in3(N__73290),
            .lcout(data_in_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78800),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_23_11_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_23_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_23_11_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i2_LC_23_11_4  (
            .in0(N__72936),
            .in1(N__70016),
            .in2(N__68756),
            .in3(N__75250),
            .lcout(\c0.data_in_frame_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78800),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_23_11_5 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_23_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_23_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_23_11_5  (
            .in0(N__68726),
            .in1(N__69548),
            .in2(N__64284),
            .in3(N__64261),
            .lcout(\c0.n22322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_23_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_23_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_23_11_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i19_LC_23_11_6  (
            .in0(N__64262),
            .in1(N__79205),
            .in2(N__69170),
            .in3(N__70017),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78800),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_23_11_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_23_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_23_11_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i1_LC_23_11_7  (
            .in0(N__70015),
            .in1(N__72937),
            .in2(N__80735),
            .in3(N__69550),
            .lcout(\c0.data_in_frame_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78800),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_3_lut_LC_23_12_0 .C_ON=1'b0;
    defparam \c0.i13_2_lut_3_lut_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_3_lut_LC_23_12_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i13_2_lut_3_lut_LC_23_12_0  (
            .in0(N__64897),
            .in1(_gnd_net_),
            .in2(N__64838),
            .in3(N__64777),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_2001_LC_23_12_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_2001_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_2001_LC_23_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_2001_LC_23_12_1  (
            .in0(N__70659),
            .in1(N__65637),
            .in2(_gnd_net_),
            .in3(N__67986),
            .lcout(\c0.n20_adj_4260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_23_12_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_23_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_LC_23_12_2  (
            .in0(_gnd_net_),
            .in1(N__64965),
            .in2(_gnd_net_),
            .in3(N__64673),
            .lcout(\c0.n7_adj_4229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_23_12_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_23_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_23_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_23_12_4  (
            .in0(N__65336),
            .in1(N__70915),
            .in2(N__69384),
            .in3(N__77857),
            .lcout(\c0.n17_adj_4219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_1194_LC_23_12_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_1194_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_1194_LC_23_12_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3_2_lut_adj_1194_LC_23_12_5  (
            .in0(N__64634),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70887),
            .lcout(\c0.n9_adj_4220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_2_lut_3_lut_4_lut_LC_23_12_6 .C_ON=1'b0;
    defparam \c0.i11_2_lut_3_lut_4_lut_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_2_lut_3_lut_4_lut_LC_23_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_2_lut_3_lut_4_lut_LC_23_12_6  (
            .in0(N__70886),
            .in1(N__64633),
            .in2(N__69884),
            .in3(N__64605),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1711_LC_23_12_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1711_LC_23_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1711_LC_23_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1711_LC_23_12_7  (
            .in0(_gnd_net_),
            .in1(N__68732),
            .in2(N__64554),
            .in3(N__69557),
            .lcout(\c0.n23406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i125_LC_23_13_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i125_LC_23_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i125_LC_23_13_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i125_LC_23_13_0  (
            .in0(N__80923),
            .in1(N__73667),
            .in2(N__66273),
            .in3(N__71781),
            .lcout(\c0.data_in_frame_15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78783),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1190_LC_23_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1190_LC_23_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1190_LC_23_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1190_LC_23_13_1  (
            .in0(_gnd_net_),
            .in1(N__64545),
            .in2(_gnd_net_),
            .in3(N__64501),
            .lcout(\c0.n22650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1598_LC_23_13_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1598_LC_23_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1598_LC_23_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1598_LC_23_13_2  (
            .in0(N__65222),
            .in1(N__65200),
            .in2(N__70598),
            .in3(N__65110),
            .lcout(),
            .ltout(\c0.n14_adj_4609_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1615_LC_23_13_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1615_LC_23_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1615_LC_23_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1615_LC_23_13_3  (
            .in0(N__70498),
            .in1(N__65160),
            .in2(N__65163),
            .in3(N__69321),
            .lcout(\c0.n22748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1974_LC_23_13_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1974_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1974_LC_23_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1974_LC_23_13_4  (
            .in0(N__65633),
            .in1(N__70645),
            .in2(_gnd_net_),
            .in3(N__65127),
            .lcout(\c0.n10_adj_4617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_2014_LC_23_13_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_2014_LC_23_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_2014_LC_23_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_2014_LC_23_13_5  (
            .in0(N__70591),
            .in1(N__65632),
            .in2(N__70658),
            .in3(N__65143),
            .lcout(),
            .ltout(\c0.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1192_LC_23_13_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1192_LC_23_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1192_LC_23_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1192_LC_23_13_6  (
            .in0(N__69320),
            .in1(N__65126),
            .in2(N__65115),
            .in3(N__65109),
            .lcout(\c0.n5813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1201_LC_23_13_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1201_LC_23_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1201_LC_23_13_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1201_LC_23_13_7  (
            .in0(N__70527),
            .in1(_gnd_net_),
            .in2(N__65035),
            .in3(_gnd_net_),
            .lcout(\c0.n13809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i94_LC_23_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i94_LC_23_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i94_LC_23_14_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i94_LC_23_14_0  (
            .in0(N__76674),
            .in1(N__73696),
            .in2(N__64987),
            .in3(N__79698),
            .lcout(\c0.data_in_frame_11_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i127_LC_23_14_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i127_LC_23_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i127_LC_23_14_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i127_LC_23_14_1  (
            .in0(N__73692),
            .in1(N__80941),
            .in2(N__70506),
            .in3(N__73336),
            .lcout(\c0.data_in_frame_15_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1515_LC_23_14_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1515_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1515_LC_23_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1515_LC_23_14_2  (
            .in0(N__64914),
            .in1(N__69609),
            .in2(N__70458),
            .in3(N__70469),
            .lcout(\c0.n22508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i73_LC_23_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i73_LC_23_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i73_LC_23_14_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i73_LC_23_14_3  (
            .in0(N__73694),
            .in1(N__74178),
            .in2(N__80747),
            .in3(N__70620),
            .lcout(\c0.data_in_frame_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_adj_1861_LC_23_14_5 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_adj_1861_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_adj_1861_LC_23_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_adj_1861_LC_23_14_5  (
            .in0(N__72559),
            .in1(N__71268),
            .in2(N__72482),
            .in3(N__72396),
            .lcout(\c0.n23_adj_4665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i123_LC_23_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i123_LC_23_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i123_LC_23_14_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i123_LC_23_14_6  (
            .in0(N__80940),
            .in1(N__73695),
            .in2(N__65368),
            .in3(N__79185),
            .lcout(\c0.data_in_frame_15_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i71_LC_23_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i71_LC_23_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i71_LC_23_14_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i71_LC_23_14_7  (
            .in0(N__73693),
            .in1(N__72940),
            .in2(N__69325),
            .in3(N__73337),
            .lcout(\c0.data_in_frame_8_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i70_LC_23_15_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i70_LC_23_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i70_LC_23_15_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i70_LC_23_15_0  (
            .in0(N__73688),
            .in1(N__72941),
            .in2(N__79728),
            .in3(N__65335),
            .lcout(\c0.data_in_frame_8_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1637_LC_23_15_1 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1637_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1637_LC_23_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1637_LC_23_15_1  (
            .in0(N__68634),
            .in1(N__70899),
            .in2(N__65304),
            .in3(N__65654),
            .lcout(),
            .ltout(\c0.n28_adj_4637_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1638_LC_23_15_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1638_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1638_LC_23_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1638_LC_23_15_2  (
            .in0(N__65253),
            .in1(N__65244),
            .in2(N__65247),
            .in3(N__65232),
            .lcout(\c0.n22319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1636_LC_23_15_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1636_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1636_LC_23_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1636_LC_23_15_3  (
            .in0(N__65493),
            .in1(N__69380),
            .in2(N__65511),
            .in3(N__70848),
            .lcout(\c0.n24_adj_4636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1635_LC_23_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1635_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1635_LC_23_15_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1635_LC_23_15_4  (
            .in0(N__66271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65238),
            .lcout(\c0.n16_adj_4635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1807_LC_23_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1807_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1807_LC_23_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1807_LC_23_15_5  (
            .in0(N__68679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65704),
            .lcout(\c0.n5_adj_4631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1596_LC_23_15_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1596_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1596_LC_23_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1596_LC_23_15_6  (
            .in0(N__65703),
            .in1(N__68633),
            .in2(N__65655),
            .in3(N__68678),
            .lcout(\c0.n13474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1191_LC_23_15_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1191_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1191_LC_23_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1191_LC_23_15_7  (
            .in0(_gnd_net_),
            .in1(N__69313),
            .in2(_gnd_net_),
            .in3(N__65640),
            .lcout(\c0.n22602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1984_LC_23_16_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1984_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1984_LC_23_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1984_LC_23_16_1  (
            .in0(N__68189),
            .in1(N__65595),
            .in2(N__65580),
            .in3(N__65553),
            .lcout(\c0.n31_adj_4743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1193_LC_23_16_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1193_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1193_LC_23_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1193_LC_23_16_2  (
            .in0(N__70847),
            .in1(N__65526),
            .in2(N__65510),
            .in3(N__65492),
            .lcout(),
            .ltout(\c0.n16_adj_4218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_4_lut_adj_1769_LC_23_16_3 .C_ON=1'b0;
    defparam \c0.i9_3_lut_4_lut_adj_1769_LC_23_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_4_lut_adj_1769_LC_23_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_3_lut_4_lut_adj_1769_LC_23_16_3  (
            .in0(N__76082),
            .in1(N__65475),
            .in2(N__65466),
            .in3(N__81057),
            .lcout(\c0.n13767 ),
            .ltout(\c0.n13767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1716_LC_23_16_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1716_LC_23_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1716_LC_23_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1716_LC_23_16_4  (
            .in0(N__71675),
            .in1(N__72196),
            .in2(N__65463),
            .in3(N__65453),
            .lcout(\c0.n6_adj_4454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1679_LC_23_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1679_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1679_LC_23_16_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1679_LC_23_16_5  (
            .in0(_gnd_net_),
            .in1(N__74961),
            .in2(_gnd_net_),
            .in3(N__65419),
            .lcout(\c0.n14_adj_4619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1418_LC_23_17_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1418_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1418_LC_23_17_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1418_LC_23_17_0  (
            .in0(N__66018),
            .in1(N__66189),
            .in2(N__66183),
            .in3(N__66162),
            .lcout(\c0.n23507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i169_LC_23_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i169_LC_23_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i169_LC_23_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i169_LC_23_17_1  (
            .in0(N__80733),
            .in1(N__66116),
            .in2(_gnd_net_),
            .in3(N__67657),
            .lcout(data_in_frame_21_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i137_LC_23_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i137_LC_23_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i137_LC_23_17_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i137_LC_23_17_2  (
            .in0(N__74187),
            .in1(N__80395),
            .in2(N__66098),
            .in3(N__80734),
            .lcout(\c0.data_in_frame_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_2_lut_3_lut_adj_2024_LC_23_17_4 .C_ON=1'b0;
    defparam \c0.i11_2_lut_3_lut_adj_2024_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_2_lut_3_lut_adj_2024_LC_23_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i11_2_lut_3_lut_adj_2024_LC_23_17_4  (
            .in0(N__72638),
            .in1(N__76052),
            .in2(_gnd_net_),
            .in3(N__66060),
            .lcout(\c0.n26_adj_4578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1239_LC_23_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1239_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1239_LC_23_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1239_LC_23_17_5  (
            .in0(_gnd_net_),
            .in1(N__65980),
            .in2(_gnd_net_),
            .in3(N__66017),
            .lcout(\c0.n22518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i144_LC_23_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i144_LC_23_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i144_LC_23_17_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i144_LC_23_17_6  (
            .in0(N__74188),
            .in1(N__76393),
            .in2(N__65987),
            .in3(N__80396),
            .lcout(\c0.data_in_frame_17_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1350_LC_23_17_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1350_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1350_LC_23_17_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_1350_LC_23_17_7  (
            .in0(N__65959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65931),
            .lcout(\c0.n5_adj_4335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1562_LC_23_18_0 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1562_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1562_LC_23_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i16_4_lut_adj_1562_LC_23_18_0  (
            .in0(N__71645),
            .in1(N__72036),
            .in2(N__65902),
            .in3(N__65861),
            .lcout(\c0.n42_adj_4589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_4_lut_adj_1693_LC_23_18_1 .C_ON=1'b0;
    defparam \c0.i11_3_lut_4_lut_adj_1693_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_4_lut_adj_1693_LC_23_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_3_lut_4_lut_adj_1693_LC_23_18_1  (
            .in0(N__65805),
            .in1(N__65786),
            .in2(N__65747),
            .in3(N__65721),
            .lcout(\c0.n24_adj_4618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i180_LC_23_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i180_LC_23_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i180_LC_23_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i180_LC_23_18_2  (
            .in0(N__77044),
            .in1(N__73750),
            .in2(_gnd_net_),
            .in3(N__78895),
            .lcout(data_in_frame_22_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1240_LC_23_18_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1240_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1240_LC_23_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1240_LC_23_18_4  (
            .in0(_gnd_net_),
            .in1(N__72017),
            .in2(_gnd_net_),
            .in3(N__66355),
            .lcout(\c0.n7_adj_4251 ),
            .ltout(\c0.n7_adj_4251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1537_LC_23_18_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1537_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1537_LC_23_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1537_LC_23_18_5  (
            .in0(N__75778),
            .in1(N__69630),
            .in2(N__66339),
            .in3(N__66333),
            .lcout(\c0.n4_adj_4568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1516_LC_23_18_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1516_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1516_LC_23_18_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1516_LC_23_18_6  (
            .in0(N__66334),
            .in1(N__66393),
            .in2(N__69640),
            .in3(N__66315),
            .lcout(\c0.n21412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i184_LC_23_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i184_LC_23_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i184_LC_23_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i184_LC_23_18_7  (
            .in0(N__78896),
            .in1(N__76289),
            .in2(_gnd_net_),
            .in3(N__66302),
            .lcout(data_in_frame_22_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i142_LC_23_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i142_LC_23_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i142_LC_23_19_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i142_LC_23_19_0  (
            .in0(N__74205),
            .in1(N__79759),
            .in2(N__66500),
            .in3(N__80415),
            .lcout(\c0.data_in_frame_17_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78766),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1626_LC_23_19_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1626_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1626_LC_23_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1626_LC_23_19_1  (
            .in0(N__66288),
            .in1(N__66272),
            .in2(N__67071),
            .in3(N__69608),
            .lcout(\c0.n15_adj_4624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i147_LC_23_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i147_LC_23_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i147_LC_23_19_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i147_LC_23_19_2  (
            .in0(N__69180),
            .in1(N__80416),
            .in2(N__79051),
            .in3(N__66242),
            .lcout(\c0.data_in_frame_18_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78766),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i149_LC_23_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i149_LC_23_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i149_LC_23_19_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i149_LC_23_19_3  (
            .in0(N__80412),
            .in1(N__69181),
            .in2(N__66220),
            .in3(N__71953),
            .lcout(\c0.data_in_frame_18_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78766),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1535_LC_23_19_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1535_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1535_LC_23_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1535_LC_23_19_4  (
            .in0(N__66666),
            .in1(N__66612),
            .in2(N__66521),
            .in3(N__66593),
            .lcout(\c0.n15_adj_4569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i152_LC_23_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i152_LC_23_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i152_LC_23_19_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i152_LC_23_19_5  (
            .in0(N__80413),
            .in1(N__69182),
            .in2(N__76325),
            .in3(N__66552),
            .lcout(\c0.data_in_frame_18_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78766),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i182_LC_23_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i182_LC_23_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i182_LC_23_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i182_LC_23_19_6  (
            .in0(N__66517),
            .in1(N__79758),
            .in2(_gnd_net_),
            .in3(N__78891),
            .lcout(data_in_frame_22_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78766),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i187_LC_23_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i187_LC_23_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i187_LC_23_19_7 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_in_frame_0__i187_LC_23_19_7  (
            .in0(N__80414),
            .in1(N__78994),
            .in2(N__80986),
            .in3(N__77266),
            .lcout(\c0.data_in_frame_23_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78766),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i181_LC_23_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i181_LC_23_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i181_LC_23_20_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i181_LC_23_20_1  (
            .in0(N__71943),
            .in1(N__75558),
            .in2(_gnd_net_),
            .in3(N__78897),
            .lcout(data_in_frame_22_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1625_LC_23_20_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1625_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1625_LC_23_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1625_LC_23_20_2  (
            .in0(N__66495),
            .in1(N__71247),
            .in2(_gnd_net_),
            .in3(N__66465),
            .lcout(),
            .ltout(\c0.n14_adj_4623_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1627_LC_23_20_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1627_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1627_LC_23_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1627_LC_23_20_3  (
            .in0(N__77573),
            .in1(N__72489),
            .in2(N__66444),
            .in3(N__66441),
            .lcout(\c0.n13963 ),
            .ltout(\c0.n13963_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1563_LC_23_20_4 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1563_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1563_LC_23_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1563_LC_23_20_4  (
            .in0(N__66435),
            .in1(N__66756),
            .in2(N__66396),
            .in3(N__66392),
            .lcout(\c0.n40_adj_4342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1526_LC_23_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1526_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1526_LC_23_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1526_LC_23_20_6  (
            .in0(N__68262),
            .in1(N__67151),
            .in2(_gnd_net_),
            .in3(N__75962),
            .lcout(\c0.n22495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i162_LC_23_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i162_LC_23_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i162_LC_23_20_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i162_LC_23_20_7  (
            .in0(N__79983),
            .in1(N__80397),
            .in2(N__75229),
            .in3(N__67070),
            .lcout(\c0.data_in_frame_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_adj_1379_LC_23_21_0 .C_ON=1'b0;
    defparam \c0.i13_2_lut_adj_1379_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_adj_1379_LC_23_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i13_2_lut_adj_1379_LC_23_21_0  (
            .in0(_gnd_net_),
            .in1(N__67055),
            .in2(_gnd_net_),
            .in3(N__67037),
            .lcout(\c0.n28_adj_4363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1483_LC_23_21_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1483_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1483_LC_23_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1483_LC_23_21_1  (
            .in0(N__77150),
            .in1(N__66984),
            .in2(N__66957),
            .in3(N__66930),
            .lcout(),
            .ltout(\c0.n10_adj_4524_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1485_LC_23_21_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1485_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1485_LC_23_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1485_LC_23_21_2  (
            .in0(_gnd_net_),
            .in1(N__75946),
            .in2(N__66903),
            .in3(N__66898),
            .lcout(\c0.n24576 ),
            .ltout(\c0.n24576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1471_LC_23_21_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1471_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1471_LC_23_21_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1471_LC_23_21_3  (
            .in0(N__66813),
            .in1(N__78025),
            .in2(N__66771),
            .in3(N__66687),
            .lcout(\c0.n14_adj_4519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1703_LC_23_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1703_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1703_LC_23_21_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1703_LC_23_21_4  (
            .in0(N__66752),
            .in1(_gnd_net_),
            .in2(N__75857),
            .in3(N__66714),
            .lcout(\c0.n22686 ),
            .ltout(\c0.n22686_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1432_LC_23_21_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1432_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1432_LC_23_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1432_LC_23_21_5  (
            .in0(N__70575),
            .in1(N__66681),
            .in2(N__66669),
            .in3(N__78024),
            .lcout(\c0.n37_adj_4473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i198_LC_23_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i198_LC_23_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i198_LC_23_21_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i198_LC_23_21_6  (
            .in0(N__72991),
            .in1(N__79703),
            .in2(N__74870),
            .in3(N__79489),
            .lcout(\c0.data_in_frame_24_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78784),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1737_LC_23_22_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1737_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1737_LC_23_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1737_LC_23_22_0  (
            .in0(N__67552),
            .in1(N__67255),
            .in2(N__77394),
            .in3(N__67501),
            .lcout(),
            .ltout(\c0.n30_adj_4489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_23_22_1 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_23_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_LC_23_22_1  (
            .in0(N__67328),
            .in1(N__67461),
            .in2(N__67455),
            .in3(N__67452),
            .lcout(),
            .ltout(\c0.n45_adj_4490_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_adj_1456_LC_23_22_2 .C_ON=1'b0;
    defparam \c0.i23_4_lut_adj_1456_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_adj_1456_LC_23_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_adj_1456_LC_23_22_2  (
            .in0(N__67335),
            .in1(N__67793),
            .in2(N__67446),
            .in3(N__67386),
            .lcout(),
            .ltout(\c0.n48_adj_4503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_1459_LC_23_22_3 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_1459_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_1459_LC_23_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_adj_1459_LC_23_22_3  (
            .in0(N__67443),
            .in1(N__67434),
            .in2(N__67422),
            .in3(N__67419),
            .lcout(\c0.n24573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_3_lut_LC_23_22_4 .C_ON=1'b0;
    defparam \c0.i16_3_lut_LC_23_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i16_3_lut_LC_23_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i16_3_lut_LC_23_22_4  (
            .in0(N__78020),
            .in1(N__77956),
            .in2(_gnd_net_),
            .in3(N__67820),
            .lcout(\c0.n41_adj_4488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_1552_LC_23_22_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_1552_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_1552_LC_23_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_1552_LC_23_22_5  (
            .in0(_gnd_net_),
            .in1(N__67380),
            .in2(_gnd_net_),
            .in3(N__67361),
            .lcout(\c0.n27_adj_4502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1740_LC_23_22_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1740_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1740_LC_23_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1740_LC_23_22_6  (
            .in0(N__67551),
            .in1(N__77391),
            .in2(N__67329),
            .in3(N__67256),
            .lcout(\c0.n21_adj_4481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1930_LC_23_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1930_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1930_LC_23_23_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1930_LC_23_23_0  (
            .in0(N__73899),
            .in1(N__67212),
            .in2(N__77189),
            .in3(N__67193),
            .lcout(\c0.n23_adj_4582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i219_LC_23_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i219_LC_23_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i219_LC_23_23_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i219_LC_23_23_1  (
            .in0(N__76693),
            .in1(N__67862),
            .in2(N__79191),
            .in3(N__79476),
            .lcout(\c0.data_in_frame_27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78801),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_LC_23_23_2 .C_ON=1'b0;
    defparam \c0.i20_3_lut_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_LC_23_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i20_3_lut_LC_23_23_2  (
            .in0(N__67824),
            .in1(N__67792),
            .in2(_gnd_net_),
            .in3(N__67773),
            .lcout(),
            .ltout(\c0.n44_adj_4471_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_adj_1434_LC_23_23_3 .C_ON=1'b0;
    defparam \c0.i23_4_lut_adj_1434_LC_23_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_adj_1434_LC_23_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_adj_1434_LC_23_23_3  (
            .in0(N__67767),
            .in1(N__67761),
            .in2(N__67752),
            .in3(N__67749),
            .lcout(),
            .ltout(\c0.n24362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1490_LC_23_23_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1490_LC_23_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1490_LC_23_23_4 .LUT_INIT=16'b1111011011111001;
    LogicCell40 \c0.i8_4_lut_adj_1490_LC_23_23_4  (
            .in0(N__67725),
            .in1(N__67716),
            .in2(N__67695),
            .in3(N__67692),
            .lcout(\c0.n26_adj_4530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i176_LC_23_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i176_LC_23_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i176_LC_23_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i176_LC_23_24_0  (
            .in0(N__77187),
            .in1(N__76274),
            .in2(_gnd_net_),
            .in3(N__67665),
            .lcout(data_in_frame_21_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78808),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1517_LC_23_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1517_LC_23_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1517_LC_23_24_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1517_LC_23_24_1  (
            .in0(_gnd_net_),
            .in1(N__73751),
            .in2(_gnd_net_),
            .in3(N__75732),
            .lcout(\c0.n22632 ),
            .ltout(\c0.n22632_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1525_LC_23_24_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1525_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1525_LC_23_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1525_LC_23_24_2  (
            .in0(_gnd_net_),
            .in1(N__73900),
            .in2(N__67566),
            .in3(N__81006),
            .lcout(\c0.n20358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1479_LC_23_24_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1479_LC_23_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1479_LC_23_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1479_LC_23_24_3  (
            .in0(N__68278),
            .in1(N__67563),
            .in2(_gnd_net_),
            .in3(N__75951),
            .lcout(),
            .ltout(\c0.n22362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1488_LC_23_24_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1488_LC_23_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1488_LC_23_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1488_LC_23_24_4  (
            .in0(N__68228),
            .in1(N__68370),
            .in2(N__68319),
            .in3(N__68316),
            .lcout(\c0.n13_adj_4527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1449_LC_23_24_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1449_LC_23_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1449_LC_23_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1449_LC_23_24_5  (
            .in0(N__68279),
            .in1(N__77351),
            .in2(N__68241),
            .in3(N__68261),
            .lcout(\c0.n12_adj_4491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i231_LC_23_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i231_LC_23_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i231_LC_23_24_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i231_LC_23_24_6  (
            .in0(N__79471),
            .in1(N__68240),
            .in2(N__80080),
            .in3(N__73330),
            .lcout(\c0.data_in_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78808),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i229_LC_23_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i229_LC_23_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i229_LC_23_24_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i229_LC_23_24_7  (
            .in0(N__80031),
            .in1(N__68229),
            .in2(N__71970),
            .in3(N__79472),
            .lcout(\c0.data_in_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78808),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1870_LC_24_9_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1870_LC_24_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1870_LC_24_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1870_LC_24_9_0  (
            .in0(N__69491),
            .in1(N__68923),
            .in2(N__68216),
            .in3(N__68646),
            .lcout(\c0.n28_adj_4286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_24_9_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_24_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_24_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i41_LC_24_9_2  (
            .in0(N__80748),
            .in1(N__69460),
            .in2(_gnd_net_),
            .in3(N__68163),
            .lcout(data_in_frame_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78819),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_3_lut_4_lut_LC_24_9_4 .C_ON=1'b0;
    defparam \c0.i18_3_lut_4_lut_LC_24_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i18_3_lut_4_lut_LC_24_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_3_lut_4_lut_LC_24_9_4  (
            .in0(N__68145),
            .in1(N__68122),
            .in2(N__68040),
            .in3(N__68847),
            .lcout(\c0.n42_adj_4746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i58_LC_24_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i58_LC_24_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i58_LC_24_9_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i58_LC_24_9_5  (
            .in0(N__75261),
            .in1(N__80843),
            .in2(N__67984),
            .in3(N__70187),
            .lcout(\c0.data_in_frame_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78819),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_LC_24_10_0 .C_ON=1'b0;
    defparam \c0.i7_2_lut_LC_24_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_LC_24_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i7_2_lut_LC_24_10_0  (
            .in0(_gnd_net_),
            .in1(N__68901),
            .in2(_gnd_net_),
            .in3(N__67934),
            .lcout(\c0.n24_adj_4213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1802_LC_24_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1802_LC_24_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1802_LC_24_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1802_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(N__68957),
            .in2(_gnd_net_),
            .in3(N__68669),
            .lcout(),
            .ltout(\c0.n6_adj_4687_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1803_LC_24_10_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1803_LC_24_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1803_LC_24_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1803_LC_24_10_2  (
            .in0(N__68793),
            .in1(N__68728),
            .in2(N__68931),
            .in3(N__68844),
            .lcout(\c0.n23274 ),
            .ltout(\c0.n23274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1319_LC_24_10_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1319_LC_24_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1319_LC_24_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1319_LC_24_10_3  (
            .in0(N__68900),
            .in1(N__69500),
            .in2(N__68892),
            .in3(N__68622),
            .lcout(\c0.n20_adj_4316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_adj_1721_LC_24_10_4 .C_ON=1'b0;
    defparam \c0.i12_3_lut_adj_1721_LC_24_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_adj_1721_LC_24_10_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i12_3_lut_adj_1721_LC_24_10_4  (
            .in0(N__68624),
            .in1(_gnd_net_),
            .in2(N__69504),
            .in3(N__68571),
            .lcout(\c0.n29_adj_4287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_4_lut_adj_1695_LC_24_10_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_4_lut_adj_1695_LC_24_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_4_lut_adj_1695_LC_24_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_3_lut_4_lut_adj_1695_LC_24_10_5  (
            .in0(N__68845),
            .in1(N__68794),
            .in2(N__68749),
            .in3(N__68670),
            .lcout(\c0.n23276 ),
            .ltout(\c0.n23276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1183_LC_24_10_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1183_LC_24_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1183_LC_24_10_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1183_LC_24_10_6  (
            .in0(N__68623),
            .in1(_gnd_net_),
            .in2(N__68607),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_24_10_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_24_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_24_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_24_10_7  (
            .in0(N__68600),
            .in1(N__68570),
            .in2(N__68559),
            .in3(N__68544),
            .lcout(\c0.n23343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_24_11_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_24_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_24_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i54_LC_24_11_0  (
            .in0(N__79622),
            .in1(N__68395),
            .in2(_gnd_net_),
            .in3(N__69264),
            .lcout(data_in_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1302_LC_24_11_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1302_LC_24_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1302_LC_24_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1302_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(N__72528),
            .in2(_gnd_net_),
            .in3(N__69547),
            .lcout(\c0.n22701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1804_LC_24_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1804_LC_24_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1804_LC_24_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1804_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(N__69262),
            .in2(_gnd_net_),
            .in3(N__71117),
            .lcout(\c0.n5_adj_4323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_24_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_24_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_24_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i42_LC_24_11_3  (
            .in0(N__69450),
            .in1(N__75251),
            .in2(_gnd_net_),
            .in3(N__70284),
            .lcout(data_in_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_89_i9_2_lut_3_lut_LC_24_11_4 .C_ON=1'b0;
    defparam \c0.equal_89_i9_2_lut_3_lut_LC_24_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.equal_89_i9_2_lut_3_lut_LC_24_11_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.equal_89_i9_2_lut_3_lut_LC_24_11_4  (
            .in0(N__74358),
            .in1(N__74631),
            .in2(_gnd_net_),
            .in3(N__74500),
            .lcout(\c0.n9 ),
            .ltout(\c0.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i145_LC_24_11_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i145_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i145_LC_24_11_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i145_LC_24_11_5  (
            .in0(N__80696),
            .in1(N__80427),
            .in2(N__69387),
            .in3(N__69275),
            .lcout(\c0.data_in_frame_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1617_LC_24_11_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1617_LC_24_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1617_LC_24_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1617_LC_24_11_6  (
            .in0(N__69376),
            .in1(N__69329),
            .in2(N__69276),
            .in3(N__69263),
            .lcout(\c0.n19_adj_4620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_24_11_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_24_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_24_11_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i18_LC_24_11_7  (
            .in0(N__69068),
            .in1(N__75252),
            .in2(N__70087),
            .in3(N__72529),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i61_LC_24_12_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i61_LC_24_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i61_LC_24_12_0 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i61_LC_24_12_0  (
            .in0(N__70193),
            .in1(N__80944),
            .in2(N__70347),
            .in3(N__71902),
            .lcout(\c0.data_in_frame_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1203_LC_24_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1203_LC_24_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1203_LC_24_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1203_LC_24_12_1  (
            .in0(_gnd_net_),
            .in1(N__69825),
            .in2(_gnd_net_),
            .in3(N__69792),
            .lcout(\c0.n22392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i78_LC_24_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i78_LC_24_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i78_LC_24_12_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i78_LC_24_12_2  (
            .in0(N__70425),
            .in1(N__73703),
            .in2(N__79649),
            .in3(N__74117),
            .lcout(\c0.data_in_frame_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_13_i3_2_lut_LC_24_12_3 .C_ON=1'b0;
    defparam \c0.select_367_Select_13_i3_2_lut_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_13_i3_2_lut_LC_24_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_13_i3_2_lut_LC_24_12_3  (
            .in0(_gnd_net_),
            .in1(N__70401),
            .in2(_gnd_net_),
            .in3(N__71529),
            .lcout(\c0.n3_adj_4410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_2_lut_3_lut_LC_24_12_4 .C_ON=1'b0;
    defparam \c0.i10_2_lut_3_lut_LC_24_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_2_lut_3_lut_LC_24_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i10_2_lut_3_lut_LC_24_12_4  (
            .in0(N__69860),
            .in1(N__70328),
            .in2(_gnd_net_),
            .in3(N__70264),
            .lcout(\c0.n40_adj_4288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i60_LC_24_12_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i60_LC_24_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i60_LC_24_12_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.data_in_frame_0__i60_LC_24_12_5  (
            .in0(N__80943),
            .in1(N__70194),
            .in2(N__77132),
            .in3(N__69861),
            .lcout(\c0.data_in_frame_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i97_LC_24_12_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i97_LC_24_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i97_LC_24_12_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i97_LC_24_12_6  (
            .in0(N__80718),
            .in1(N__79948),
            .in2(N__69833),
            .in3(N__73704),
            .lcout(\c0.data_in_frame_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i98_LC_24_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i98_LC_24_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i98_LC_24_12_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i98_LC_24_12_7  (
            .in0(N__73702),
            .in1(N__75257),
            .in2(N__80009),
            .in3(N__69793),
            .lcout(\c0.data_in_frame_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78802),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_2020_LC_24_13_0 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_2020_LC_24_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_2020_LC_24_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_2020_LC_24_13_0  (
            .in0(N__70683),
            .in1(N__69761),
            .in2(N__70971),
            .in3(N__69702),
            .lcout(\c0.n13253 ),
            .ltout(\c0.n13253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1624_LC_24_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1624_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1624_LC_24_13_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1624_LC_24_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69648),
            .in3(N__69644),
            .lcout(\c0.n22828 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_2018_LC_24_13_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_2018_LC_24_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_2018_LC_24_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_2018_LC_24_13_2  (
            .in0(N__70788),
            .in1(N__70749),
            .in2(N__70716),
            .in3(N__70701),
            .lcout(\c0.n27_adj_4748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i92_LC_24_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i92_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i92_LC_24_14_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i92_LC_24_14_0  (
            .in0(N__73690),
            .in1(N__76530),
            .in2(N__70673),
            .in3(N__77091),
            .lcout(\c0.data_in_frame_11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1178_LC_24_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1178_LC_24_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1178_LC_24_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1178_LC_24_14_2  (
            .in0(_gnd_net_),
            .in1(N__70850),
            .in2(_gnd_net_),
            .in3(N__70619),
            .lcout(\c0.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i159_LC_24_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i159_LC_24_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i159_LC_24_14_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i159_LC_24_14_3  (
            .in0(N__80399),
            .in1(N__76529),
            .in2(N__77649),
            .in3(N__73276),
            .lcout(\c0.data_in_frame_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i228_LC_24_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i228_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i228_LC_24_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i228_LC_24_14_4  (
            .in0(N__79491),
            .in1(N__79952),
            .in2(N__70571),
            .in3(N__77090),
            .lcout(\c0.data_in_frame_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i126_LC_24_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i126_LC_24_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i126_LC_24_14_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i126_LC_24_14_6  (
            .in0(N__73689),
            .in1(N__80942),
            .in2(N__71246),
            .in3(N__79702),
            .lcout(\c0.data_in_frame_15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i100_LC_24_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i100_LC_24_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i100_LC_24_14_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i100_LC_24_14_7  (
            .in0(N__77092),
            .in1(N__73691),
            .in2(N__70550),
            .in3(N__79947),
            .lcout(\c0.data_in_frame_12_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1727_LC_24_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1727_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1727_LC_24_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1727_LC_24_15_0  (
            .in0(_gnd_net_),
            .in1(N__70505),
            .in2(_gnd_net_),
            .in3(N__71674),
            .lcout(\c0.n22379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1514_LC_24_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1514_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1514_LC_24_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1514_LC_24_15_1  (
            .in0(_gnd_net_),
            .in1(N__73055),
            .in2(_gnd_net_),
            .in3(N__71269),
            .lcout(\c0.n6_adj_4559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i143_LC_24_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i143_LC_24_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i143_LC_24_15_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i143_LC_24_15_3  (
            .in0(N__74116),
            .in1(N__80385),
            .in2(N__73307),
            .in3(N__71270),
            .lcout(\c0.data_in_frame_17_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1715_LC_24_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1715_LC_24_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1715_LC_24_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1715_LC_24_15_4  (
            .in0(N__71242),
            .in1(N__72195),
            .in2(_gnd_net_),
            .in3(N__71673),
            .lcout(\c0.n22605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_2016_LC_24_15_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_2016_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_2016_LC_24_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_2016_LC_24_15_5  (
            .in0(N__71219),
            .in1(N__71175),
            .in2(N__71148),
            .in3(N__71126),
            .lcout(\c0.n30_adj_4747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1634_LC_24_15_7 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1634_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1634_LC_24_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1634_LC_24_15_7  (
            .in0(N__70959),
            .in1(N__70932),
            .in2(N__72464),
            .in3(N__70922),
            .lcout(\c0.n25_adj_4633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i76_LC_24_16_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i76_LC_24_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i76_LC_24_16_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i76_LC_24_16_0  (
            .in0(N__74157),
            .in1(N__73687),
            .in2(N__77133),
            .in3(N__70876),
            .lcout(\c0.data_in_frame_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i91_LC_24_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i91_LC_24_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i91_LC_24_16_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i91_LC_24_16_1  (
            .in0(N__73686),
            .in1(N__76525),
            .in2(N__79184),
            .in3(N__70849),
            .lcout(\c0.data_in_frame_11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i226_LC_24_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i226_LC_24_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i226_LC_24_16_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i226_LC_24_16_2  (
            .in0(N__79490),
            .in1(N__75178),
            .in2(N__70808),
            .in3(N__80008),
            .lcout(\c0.data_in_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i108_LC_24_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i108_LC_24_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i108_LC_24_16_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i108_LC_24_16_3  (
            .in0(N__75399),
            .in1(N__77124),
            .in2(N__72215),
            .in3(N__75507),
            .lcout(\c0.data_in_frame_13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1236_LC_24_16_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1236_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1236_LC_24_16_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1236_LC_24_16_4  (
            .in0(_gnd_net_),
            .in1(N__77440),
            .in2(_gnd_net_),
            .in3(N__77405),
            .lcout(\c0.n14081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i107_LC_24_16_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i107_LC_24_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i107_LC_24_16_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i107_LC_24_16_5  (
            .in0(N__75398),
            .in1(N__75506),
            .in2(N__79183),
            .in3(N__72463),
            .lcout(\c0.data_in_frame_13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78767),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_4_lut_adj_2033_LC_24_16_6 .C_ON=1'b0;
    defparam \c0.i3_2_lut_4_lut_adj_2033_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_4_lut_adj_2033_LC_24_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_4_lut_adj_2033_LC_24_16_6  (
            .in0(N__72152),
            .in1(N__72252),
            .in2(N__72214),
            .in3(N__72318),
            .lcout(\c0.n16_adj_4627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1685_LC_24_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1685_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1685_LC_24_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1685_LC_24_16_7  (
            .in0(N__72251),
            .in1(N__72206),
            .in2(_gnd_net_),
            .in3(N__72153),
            .lcout(\c0.n4_adj_4586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1238_LC_24_17_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1238_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1238_LC_24_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1238_LC_24_17_1  (
            .in0(N__72111),
            .in1(N__72090),
            .in2(N__72060),
            .in3(N__72032),
            .lcout(\c0.n10_adj_4250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i133_LC_24_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i133_LC_24_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i133_LC_24_17_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i133_LC_24_17_3  (
            .in0(N__72938),
            .in1(N__80431),
            .in2(N__71946),
            .in3(N__71988),
            .lcout(\c0.data_in_frame_16_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i109_LC_24_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i109_LC_24_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i109_LC_24_17_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i109_LC_24_17_4  (
            .in0(N__75500),
            .in1(N__75415),
            .in2(N__71679),
            .in3(N__71906),
            .lcout(\c0.data_in_frame_13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1709_LC_24_17_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1709_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1709_LC_24_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1709_LC_24_17_6  (
            .in0(_gnd_net_),
            .in1(N__73081),
            .in2(_gnd_net_),
            .in3(N__71627),
            .lcout(\c0.n16_adj_4666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_367_Select_18_i3_2_lut_LC_24_17_7 .C_ON=1'b0;
    defparam \c0.select_367_Select_18_i3_2_lut_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_367_Select_18_i3_2_lut_LC_24_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_367_Select_18_i3_2_lut_LC_24_17_7  (
            .in0(_gnd_net_),
            .in1(N__71589),
            .in2(_gnd_net_),
            .in3(N__71544),
            .lcout(\c0.n3_adj_4400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i178_LC_24_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i178_LC_24_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i178_LC_24_18_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.data_in_frame_0__i178_LC_24_18_0  (
            .in0(_gnd_net_),
            .in1(N__75177),
            .in2(N__73083),
            .in3(N__78890),
            .lcout(data_in_frame_22_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i121_LC_24_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i121_LC_24_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i121_LC_24_18_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i121_LC_24_18_2  (
            .in0(N__80973),
            .in1(N__73706),
            .in2(N__73396),
            .in3(N__80719),
            .lcout(\c0.data_in_frame_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i191_LC_24_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i191_LC_24_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i191_LC_24_18_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i191_LC_24_18_3  (
            .in0(N__73300),
            .in1(N__80323),
            .in2(N__75830),
            .in3(N__80974),
            .lcout(\c0.data_in_frame_23_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1378_LC_24_18_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1378_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1378_LC_24_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1378_LC_24_18_4  (
            .in0(N__75566),
            .in1(N__73734),
            .in2(N__73082),
            .in3(N__75823),
            .lcout(\c0.n29_adj_4362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i163_LC_24_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i163_LC_24_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i163_LC_24_18_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i163_LC_24_18_5  (
            .in0(N__80007),
            .in1(N__80322),
            .in2(N__73059),
            .in3(N__79148),
            .lcout(\c0.data_in_frame_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i190_LC_24_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i190_LC_24_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i190_LC_24_18_6 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_in_frame_0__i190_LC_24_18_6  (
            .in0(N__80320),
            .in1(N__80975),
            .in2(N__79756),
            .in3(N__73020),
            .lcout(\c0.data_in_frame_23_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i136_LC_24_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i136_LC_24_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i136_LC_24_18_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i136_LC_24_18_7  (
            .in0(N__72939),
            .in1(N__80321),
            .in2(N__72682),
            .in3(N__76293),
            .lcout(\c0.data_in_frame_16_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1616_LC_24_19_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1616_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1616_LC_24_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1616_LC_24_19_0  (
            .in0(N__72642),
            .in1(N__72612),
            .in2(N__72606),
            .in3(N__72587),
            .lcout(\c0.n22288 ),
            .ltout(\c0.n22288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1862_LC_24_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1862_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1862_LC_24_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1862_LC_24_19_1  (
            .in0(_gnd_net_),
            .in1(N__72472),
            .in2(N__72417),
            .in3(N__72413),
            .lcout(\c0.n14160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i138_LC_24_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i138_LC_24_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i138_LC_24_19_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i138_LC_24_19_2  (
            .in0(N__80401),
            .in1(N__74156),
            .in2(N__74712),
            .in3(N__75047),
            .lcout(\c0.data_in_frame_17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1998_LC_24_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1998_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1998_LC_24_19_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1998_LC_24_19_3  (
            .in0(N__74678),
            .in1(N__74524),
            .in2(N__74388),
            .in3(N__80400),
            .lcout(n22110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i202_LC_24_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i202_LC_24_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i202_LC_24_19_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i202_LC_24_19_4  (
            .in0(N__74206),
            .in1(N__75046),
            .in2(N__73939),
            .in3(N__79481),
            .lcout(\c0.data_in_frame_25_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i161_LC_24_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i161_LC_24_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i161_LC_24_19_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i161_LC_24_19_5  (
            .in0(N__80095),
            .in1(N__80617),
            .in2(N__73901),
            .in3(N__80403),
            .lcout(\c0.data_in_frame_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i153_LC_24_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i153_LC_24_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i153_LC_24_19_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i153_LC_24_19_7  (
            .in0(N__76683),
            .in1(N__80402),
            .in2(N__73863),
            .in3(N__80618),
            .lcout(\c0.data_in_frame_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1528_LC_24_20_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1528_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1528_LC_24_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1528_LC_24_20_0  (
            .in0(N__75614),
            .in1(N__74772),
            .in2(N__75562),
            .in3(N__75708),
            .lcout(\c0.n12_adj_4564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1726_LC_24_20_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1726_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1726_LC_24_20_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1726_LC_24_20_1  (
            .in0(N__75785),
            .in1(N__73796),
            .in2(_gnd_net_),
            .in3(N__75729),
            .lcout(\c0.n6_adj_4462 ),
            .ltout(\c0.n6_adj_4462_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_3_lut_LC_24_20_2 .C_ON=1'b0;
    defparam \c0.i12_2_lut_3_lut_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_3_lut_LC_24_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i12_2_lut_3_lut_LC_24_20_2  (
            .in0(_gnd_net_),
            .in1(N__75548),
            .in2(N__73776),
            .in3(N__75612),
            .lcout(\c0.n22562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_rep_362_2_lut_3_lut_LC_24_20_3 .C_ON=1'b0;
    defparam \c0.i6_rep_362_2_lut_3_lut_LC_24_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_rep_362_2_lut_3_lut_LC_24_20_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i6_rep_362_2_lut_3_lut_LC_24_20_3  (
            .in0(N__74773),
            .in1(_gnd_net_),
            .in2(N__73752),
            .in3(N__75731),
            .lcout(\c0.n25484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_24_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_24_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_24_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_24_20_4  (
            .in0(N__75549),
            .in1(N__75613),
            .in2(N__75996),
            .in3(N__76726),
            .lcout(\c0.n22769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1428_LC_24_20_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1428_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1428_LC_24_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1428_LC_24_20_6  (
            .in0(N__75947),
            .in1(N__75873),
            .in2(N__75858),
            .in3(N__75810),
            .lcout(\c0.n14_adj_4465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1389_LC_24_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1389_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1389_LC_24_20_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1389_LC_24_20_7  (
            .in0(N__75786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75730),
            .lcout(\c0.n4_adj_4369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_3_lut_4_lut_LC_24_21_0 .C_ON=1'b0;
    defparam \c0.i31_3_lut_4_lut_LC_24_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i31_3_lut_4_lut_LC_24_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i31_3_lut_4_lut_LC_24_21_0  (
            .in0(N__74768),
            .in1(N__75553),
            .in2(N__75701),
            .in3(N__75620),
            .lcout(\c0.n73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_2_lut_LC_24_21_1 .C_ON=1'b0;
    defparam \c0.i20_2_lut_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20_2_lut_LC_24_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i20_2_lut_LC_24_21_1  (
            .in0(N__75621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75554),
            .lcout(\c0.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i106_LC_24_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i106_LC_24_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i106_LC_24_21_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i106_LC_24_21_3  (
            .in0(N__75492),
            .in1(N__75416),
            .in2(N__75228),
            .in3(N__74933),
            .lcout(\c0.data_in_frame_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1592_LC_24_21_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1592_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1592_LC_24_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1592_LC_24_21_5  (
            .in0(N__77392),
            .in1(N__74903),
            .in2(N__74866),
            .in3(N__74841),
            .lcout(\c0.n6718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1714_LC_24_21_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1714_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1714_LC_24_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1714_LC_24_21_6  (
            .in0(N__81002),
            .in1(N__77298),
            .in2(N__74774),
            .in3(N__74745),
            .lcout(\c0.n20239 ),
            .ltout(\c0.n20239_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1423_LC_24_21_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1423_LC_24_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1423_LC_24_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1423_LC_24_21_7  (
            .in0(N__77393),
            .in1(N__79226),
            .in2(N__77355),
            .in3(N__77352),
            .lcout(\c0.n10_adj_4457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1773_LC_24_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1773_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1773_LC_24_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1773_LC_24_22_3  (
            .in0(N__77188),
            .in1(N__77726),
            .in2(_gnd_net_),
            .in3(N__77217),
            .lcout(\c0.n6_adj_4668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1560_LC_24_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1560_LC_24_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1560_LC_24_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1560_LC_24_22_5  (
            .in0(_gnd_net_),
            .in1(N__77280),
            .in2(_gnd_net_),
            .in3(N__76797),
            .lcout(\c0.n13314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1774_LC_24_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1774_LC_24_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1774_LC_24_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1774_LC_24_23_0  (
            .in0(N__77216),
            .in1(N__77180),
            .in2(_gnd_net_),
            .in3(N__77638),
            .lcout(\c0.n20350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i188_LC_24_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i188_LC_24_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i188_LC_24_23_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_in_frame_0__i188_LC_24_23_2  (
            .in0(N__80987),
            .in1(N__77058),
            .in2(N__76815),
            .in3(N__80433),
            .lcout(\c0.data_in_frame_23_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1444_LC_24_23_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1444_LC_24_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1444_LC_24_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1444_LC_24_23_3  (
            .in0(N__76776),
            .in1(N__76767),
            .in2(N__76758),
            .in3(N__76741),
            .lcout(\c0.n30_adj_4482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i160_LC_24_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i160_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i160_LC_24_23_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i160_LC_24_23_6  (
            .in0(N__76582),
            .in1(N__80432),
            .in2(N__77569),
            .in3(N__76394),
            .lcout(\c0.data_in_frame_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_1647_LC_26_16_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_1647_LC_26_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_1647_LC_26_16_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_1647_LC_26_16_5  (
            .in0(_gnd_net_),
            .in1(N__76086),
            .in2(_gnd_net_),
            .in3(N__76053),
            .lcout(\c0.n19_adj_4595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_26_19_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_26_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_26_19_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i5_2_lut_LC_26_19_1  (
            .in0(N__77883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77817),
            .lcout(\c0.n18 ),
            .ltout(\c0.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1710_LC_26_19_2 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1710_LC_26_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1710_LC_26_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1710_LC_26_19_2  (
            .in0(N__81103),
            .in1(N__77501),
            .in2(N__77754),
            .in3(N__77489),
            .lcout(\c0.n28_adj_4667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_4_lut_LC_26_19_4 .C_ON=1'b0;
    defparam \c0.i9_3_lut_4_lut_LC_26_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_4_lut_LC_26_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_3_lut_4_lut_LC_26_19_4  (
            .in0(N__77453),
            .in1(N__77508),
            .in2(N__77655),
            .in3(N__77417),
            .lcout(),
            .ltout(\c0.n24_adj_4653_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1712_LC_26_19_5 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1712_LC_26_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1712_LC_26_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1712_LC_26_19_5  (
            .in0(N__77751),
            .in1(N__77739),
            .in2(N__77733),
            .in3(N__81071),
            .lcout(\c0.n22369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_1650_LC_26_19_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_1650_LC_26_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_1650_LC_26_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_1650_LC_26_19_7  (
            .in0(_gnd_net_),
            .in1(N__77709),
            .in2(_gnd_net_),
            .in3(N__77687),
            .lcout(\c0.n17_adj_4626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1669_LC_26_20_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1669_LC_26_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1669_LC_26_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1669_LC_26_20_4  (
            .in0(N__77650),
            .in1(N__77574),
            .in2(_gnd_net_),
            .in3(N__77517),
            .lcout(\c0.n15_adj_4625 ),
            .ltout(\c0.n15_adj_4625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1628_LC_26_20_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1628_LC_26_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1628_LC_26_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1628_LC_26_20_5  (
            .in0(N__77502),
            .in1(N__77490),
            .in2(N__77466),
            .in3(N__77463),
            .lcout(\c0.n24_adj_4628 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1692_LC_26_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1692_LC_26_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1692_LC_26_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1692_LC_26_21_1  (
            .in0(N__78841),
            .in1(N__77457),
            .in2(_gnd_net_),
            .in3(N__77421),
            .lcout(),
            .ltout(\c0.n14_adj_4629_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1629_LC_26_21_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1629_LC_26_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1629_LC_26_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1629_LC_26_21_2  (
            .in0(N__81104),
            .in1(N__81081),
            .in2(N__81075),
            .in3(N__81072),
            .lcout(\c0.n22234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i185_LC_26_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i185_LC_26_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i185_LC_26_21_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_in_frame_0__i185_LC_26_21_3  (
            .in0(N__80918),
            .in1(N__80729),
            .in2(N__80131),
            .in3(N__80430),
            .lcout(\c0.data_in_frame_23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78811),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i230_LC_26_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i230_LC_26_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i230_LC_26_21_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i230_LC_26_21_4  (
            .in0(N__80051),
            .in1(N__79757),
            .in2(N__79227),
            .in3(N__79488),
            .lcout(\c0.data_in_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78811),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i179_LC_26_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i179_LC_26_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i179_LC_26_21_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i179_LC_26_21_6  (
            .in0(N__79192),
            .in1(N__78842),
            .in2(_gnd_net_),
            .in3(N__78911),
            .lcout(data_in_frame_22_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__78811),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_1491_LC_26_23_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_1491_LC_26_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_1491_LC_26_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_1491_LC_26_23_5  (
            .in0(_gnd_net_),
            .in1(N__78027),
            .in2(_gnd_net_),
            .in3(N__77954),
            .lcout(\c0.n24_adj_4531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
